//# 38 inputs
//# 304 outputs
//# 1426 D-type flipflops
//# 7805 inverters
//# 11448 gates (5516 ANDs + 2126 NANDs + 2621 ORs + 1185 NORs)



module s38584 (clock, g35, g36, g6744, g6745, g6746, g6747,
     g6748, g6749, g6750, g6751, g6752, g6753, g7243, g7245, g7257,
     g7260, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277,
     g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g8403,
     g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788,
     g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920,
     g9019, g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680,
     g9682, g9741, g9743, g9817, g10122, g10306, g10500, g10527,
     g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238,
     g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923,
     g13039, g13049, g13068, g13085, g13099, g13259, g13272, g13865,
     g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147,
     g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597,
     g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779,
     g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693,
     g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955,
     g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577,
     g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678,
     g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760,
     g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092,
     g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101,
     g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763,
     g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727,
     g23002, g23190, g23612, g23652, g23683, g23759, g24151, g25114,
     g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586,
     g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877,
     g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212,
     g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220,
     g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656,
     g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429,
     g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874,
     g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950,
     g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236,
     g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436,
     g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919,
     g34921, g34923, g34925, g34927, g34956, g34972);
  input clock, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749,
       g6750, g6751, g6752, g6753;
  output g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178,
       g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353,
       g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785,
       g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917,
       g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
       g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306,
       g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770,
       g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832,
       g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259,
       g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096,
       g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451,
       g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738,
       g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659,
       g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874,
       g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423,
       g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649,
       g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739,
       g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845,
       g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099,
       g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652,
       g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292,
       g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759,
       g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584,
       g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875,
       g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210,
       g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218,
       g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332,
       g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863,
       g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636,
       g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948,
       g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234,
       g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425,
       g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915,
       g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972;
  wire clock, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749,
       g6750, g6751, g6752, g6753;
  wire g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178,
       g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353,
       g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785,
       g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917,
       g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
       g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306,
       g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770,
       g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832,
       g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259,
       g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096,
       g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451,
       g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738,
       g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659,
       g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874,
       g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423,
       g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649,
       g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739,
       g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845,
       g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099,
       g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652,
       g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292,
       g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759,
       g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584,
       g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875,
       g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210,
       g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218,
       g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332,
       g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863,
       g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636,
       g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948,
       g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234,
       g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425,
       g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915,
       g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972;
  wire g37, g55, g142, g146, g150, g153, g157, g160;
  wire g164, g168, g174, g182, g191, g203, g209, g218;
  wire g222, g225, g232, g239, g246, g255, g262, g269;
  wire g278, g283, g287, g291, g294, g298, g301, g305;
  wire g311, g316, g319, g324, g329, g333, g336, g341;
  wire g347, g351, g355, g358, g370, g376, g385, g392;
  wire g401, g405, g411, g417, g424, g429, g433, g437;
  wire g441, g446, g452, g460, g475, g479, g482, g490;
  wire g496, g499, g504, g513, g518, g534, g538, g542;
  wire g546, g550, g554, g645, g650, g655, g661, g667;
  wire g671, g676, g681, g686, g691, g699, g703, g718;
  wire g723, g728, g732, g736, g739, g744, g749, g753;
  wire g758, g763, g767, g772, g776, g781, g785, g790;
  wire g794, g807, g812, g817, g822, g827, g832, g837;
  wire g843, g847, g854, g862, g872, g890, g896, g956;
  wire g962, g969, g976, g979, g990, g996, g1002, g1008;
  wire g1018, g1024, g1030, g1036, g1041, g1046, g1052, g1061;
  wire g1070, g1087, g1094, g1099, g1105, g1111, g1124, g1129;
  wire g1135, g1141, g1146, g1152, g1171, g1178, g1183, g1189;
  wire g1193, g1199, g1205, g1211, g1216, g1221, g1236, g1300;
  wire g1306, g1312, g1319, g1322, g1333, g1339, g1345, g1351;
  wire g1361, g1367, g1373, g1379, g1384, g1389, g1395, g1404;
  wire g1413, g1430, g1437, g1442, g1448, g1454, g1467, g1472;
  wire g1478, g1484, g1489, g1495, g1514, g1521, g1526, g1532;
  wire g1536, g1542, g1548, g1554, g1559, g1564, g1579, g1585;
  wire g1592, g1600, g1604, g1608, g1612, g1616, g1620, g1624;
  wire g1632, g1636, g1644, g1648, g1657, g1664, g1668, g1677;
  wire g1682, g1687, g1691, g1696, g1700, g1706, g1710, g1714;
  wire g1720, g1724, g1728, g1736, g1740, g1744, g1748, g1752;
  wire g1756, g1760, g1768, g1772, g1779, g1783, g1792, g1798;
  wire g1802, g1811, g1816, g1821, g1825, g1830, g1834, g1840;
  wire g1844, g1848, g1854, g1858, g1862, g1870, g1874, g1878;
  wire g1882, g1886, g1890, g1894, g1902, g1906, g1913, g1917;
  wire g1926, g1932, g1936, g1945, g1950, g1955, g1959, g1964;
  wire g1968, g1974, g1978, g1982, g1988, g1992, g1996, g2004;
  wire g2008, g2012, g2016, g2020, g2024, g2028, g2036, g2040;
  wire g2047, g2051, g2060, g2066, g2070, g2079, g2084, g2089;
  wire g2093, g2098, g2102, g2108, g2112, g2116, g2122, g2126;
  wire g2153, g2161, g2165, g2169, g2173, g2177, g2181, g2185;
  wire g2193, g2197, g2204, g2208, g2217, g2223, g2227, g2236;
  wire g2241, g2246, g2250, g2255, g2259, g2265, g2269, g2273;
  wire g2279, g2283, g2287, g2295, g2299, g2303, g2307, g2311;
  wire g2315, g2319, g2327, g2331, g2338, g2342, g2351, g2357;
  wire g2361, g2370, g2375, g2380, g2384, g2389, g2393, g2399;
  wire g2403, g2407, g2413, g2417, g2421, g2429, g2433, g2437;
  wire g2441, g2445, g2449, g2453, g2461, g2465, g2472, g2476;
  wire g2485, g2491, g2495, g2504, g2509, g2514, g2518, g2523;
  wire g2527, g2533, g2537, g2541, g2547, g2551, g2555, g2563;
  wire g2567, g2571, g2575, g2579, g2583, g2587, g2595, g2599;
  wire g2606, g2610, g2619, g2625, g2629, g2638, g2643, g2648;
  wire g2652, g2657, g2661, g2667, g2671, g2675, g2681, g2685;
  wire g2724, g2729, g2735, g2759, g2763, g2767, g2771, g2775;
  wire g2779, g2783, g2787, g2791, g2795, g2799, g2803, g2807;
  wire g2811, g2815, g2819, g2823, g2827, g2831, g2834, g2844;
  wire g2848, g2852, g2856, g2860, g2864, g2868, g2873, g2878;
  wire g2882, g2886, g2890, g2894, g2898, g2902, g2907, g2912;
  wire g2917, g2922, g2927, g2932, g2936, g2941, g2946, g2950;
  wire g2955, g2960, g2965, g2970, g2975, g2980, g2984, g2988;
  wire g2994, g2999, g3003, g3050, g3100, g3106, g3111, g3115;
  wire g3119, g3125, g3129, g3133, g3139, g3143, g3147, g3155;
  wire g3161, g3171, g3179, g3187, g3191, g3195, g3199, g3203;
  wire g3207, g3211, g3215, g3219, g3223, g3227, g3231, g3235;
  wire g3239, g3243, g3247, g3251, g3255, g3259, g3263, g3329;
  wire g3333, g3338, g3343, g3347, g3401, g3451, g3457, g3462;
  wire g3466, g3470, g3476, g3480, g3484, g3490, g3494, g3498;
  wire g3506, g3512, g3522, g3530, g3538, g3542, g3546, g3550;
  wire g3554, g3558, g3562, g3566, g3570, g3574, g3578, g3582;
  wire g3586, g3590, g3594, g3598, g3602, g3606, g3610, g3614;
  wire g3680, g3684, g3689, g3694, g3698, g3752, g3802, g3808;
  wire g3813, g3817, g3821, g3827, g3831, g3835, g3841, g3845;
  wire g3849, g3857, g3863, g3873, g3881, g3889, g3893, g3897;
  wire g3901, g3905, g3909, g3913, g3917, g3921, g3925, g3929;
  wire g3933, g3937, g3941, g3945, g3949, g3953, g3957, g3961;
  wire g3965, g4031, g4035, g4040, g4045, g4049, g4057, g4064;
  wire g4072, g4076, g4082, g4087, g4093, g4098, g4104, g4108;
  wire g4112, g4116, g4119, g4122, g4141, g4146, g4153, g4157;
  wire g4172, g4176, g4180, g4235, g4239, g4242, g4245, g4249;
  wire g4253, g4258, g4264, g4269, g4273, g4281, g4291, g4297;
  wire g4300, g4308, g4311, g4322, g4340, g4349, g4358, g4366;
  wire g4369, g4375, g4382, g4388, g4392, g4401, g4405, g4411;
  wire g4417, g4420, g4423, g4427, g4430, g4434, g4438, g4443;
  wire g4452, g4455, g4456, g4459, g4462, g4467, g4477, g4480;
  wire g4483, g4486, g4489, g4492, g4495, g4498, g4501, g4504;
  wire g4512, g4515, g4519, g4521, g4527, g4531, g4534, g4540;
  wire g4543, g4546, g4549, g4552, g4555, g4558, g4561, g4564;
  wire g4567, g4570, g4572, g4575, g4578, g4584, g4593, g4601;
  wire g4608, g4621, g4628, g4633, g4643, g4646, g4653, g4659;
  wire g4664, g4669, g4674, g4681, g4688, g4698, g4704, g4709;
  wire g4743, g4749, g4754, g4760, g4765, g4771, g4776, g4785;
  wire g4793, g4801, g4821, g4826, g4831, g4836, g4843, g4849;
  wire g4854, g4859, g4864, g4871, g4878, g4888, g4894, g4899;
  wire g4933, g4939, g4944, g4950, g4955, g4961, g4966, g4975;
  wire g4983, g4991, g5011, g5016, g5022, g5029, g5033, g5037;
  wire g5041, g5046, g5052, g5057, g5062, g5069, g5073, g5077;
  wire g5080, g5084, g5092, g5097, g5109, g5112, g5115, g5120;
  wire g5124, g5128, g5134, g5138, g5142, g5148, g5152, g5156;
  wire g5164, g5170, g5180, g5188, g5196, g5200, g5204, g5208;
  wire g5212, g5216, g5220, g5224, g5228, g5232, g5236, g5240;
  wire g5244, g5248, g5252, g5256, g5260, g5264, g5268, g5272;
  wire g5297, g5339, g5348, g5352, g5406, g5456, g5462, g5467;
  wire g5471, g5475, g5481, g5485, g5489, g5495, g5499, g5503;
  wire g5511, g5517, g5527, g5535, g5543, g5547, g5551, g5555;
  wire g5559, g5563, g5567, g5571, g5575, g5579, g5583, g5587;
  wire g5591, g5595, g5599, g5603, g5607, g5611, g5615, g5619;
  wire g5685, g5689, g5694, g5698, g5752, g5802, g5808, g5813;
  wire g5817, g5821, g5827, g5831, g5835, g5841, g5845, g5849;
  wire g5857, g5863, g5873, g5881, g5889, g5893, g5897, g5901;
  wire g5905, g5909, g5913, g5917, g5921, g5925, g5929, g5933;
  wire g5937, g5941, g5945, g5949, g5953, g5957, g5961, g5965;
  wire g6031, g6035, g6040, g6044, g6098, g6148, g6154, g6159;
  wire g6163, g6167, g6173, g6177, g6181, g6187, g6191, g6195;
  wire g6203, g6209, g6219, g6227, g6235, g6239, g6243, g6247;
  wire g6251, g6255, g6259, g6263, g6267, g6271, g6275, g6279;
  wire g6283, g6287, g6291, g6295, g6299, g6303, g6307, g6311;
  wire g6377, g6381, g6386, g6390, g6444, g6494, g6500, g6505;
  wire g6509, g6513, g6519, g6523, g6527, g6533, g6537, g6541;
  wire g6549, g6555, g6565, g6573, g6581, g6585, g6589, g6593;
  wire g6597, g6601, g6605, g6609, g6613, g6617, g6621, g6625;
  wire g6629, g6633, g6637, g6641, g6645, g6649, g6653, g6657;
  wire g6723, g6727, g6732, g6736, g_5902, g_5903, n_0, n_1;
  wire n_2, n_3, n_4, n_5, n_6, n_7, n_9, n_10;
  wire n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18;
  wire n_20, n_21, n_22, n_23, n_24, n_26, n_27, n_29;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_41, n_42, n_43, n_44, n_46, n_47;
  wire n_49, n_50, n_52, n_53, n_54, n_56, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_66, n_67, n_68, n_70;
  wire n_71, n_72, n_74, n_77, n_80, n_81, n_83, n_85;
  wire n_86, n_87, n_88, n_90, n_91, n_96, n_99, n_102;
  wire n_103, n_104, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_113, n_117, n_120, n_122, n_123, n_126, n_127, n_128;
  wire n_129, n_130, n_132, n_134, n_135, n_136, n_137, n_139;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_150, n_151, n_152, n_155, n_156, n_159, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_169, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179;
  wire n_181, n_182, n_183, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_203, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_218, n_219;
  wire n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_237;
  wire n_238, n_239, n_241, n_242, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431;
  wire n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439;
  wire n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_531, n_532, n_533, n_534, n_535;
  wire n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543;
  wire n_544, n_545, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560;
  wire n_561, n_564, n_565, n_566, n_567, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_577, n_578, n_579;
  wire n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587;
  wire n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595;
  wire n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603;
  wire n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611;
  wire n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619;
  wire n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627;
  wire n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635;
  wire n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643;
  wire n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651;
  wire n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659;
  wire n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667;
  wire n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683;
  wire n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691;
  wire n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755;
  wire n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763;
  wire n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779;
  wire n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787;
  wire n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811;
  wire n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819;
  wire n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827;
  wire n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835;
  wire n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843;
  wire n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851;
  wire n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859;
  wire n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867;
  wire n_868, n_869, n_870, n_871, n_872, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884;
  wire n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892;
  wire n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900;
  wire n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956;
  wire n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964;
  wire n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972;
  wire n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980;
  wire n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988;
  wire n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996;
  wire n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004;
  wire n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012;
  wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028;
  wire n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036;
  wire n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044;
  wire n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052;
  wire n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060;
  wire n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068;
  wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086;
  wire n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1097, n_1099;
  wire n_1100, n_1101, n_1103, n_1105, n_1106, n_1109, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135;
  wire n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143;
  wire n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151;
  wire n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159;
  wire n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167;
  wire n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175;
  wire n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183;
  wire n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191;
  wire n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1218;
  wire n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226;
  wire n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234;
  wire n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242;
  wire n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250;
  wire n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258;
  wire n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266;
  wire n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274;
  wire n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282;
  wire n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290;
  wire n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298;
  wire n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306;
  wire n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314;
  wire n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322;
  wire n_1323, n_1324, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331;
  wire n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339;
  wire n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347;
  wire n_1348, n_1349, n_1350, n_1351, n_1352, n_1354, n_1355, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413;
  wire n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421;
  wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
  wire n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437;
  wire n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445;
  wire n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1460, n_1461, n_1462;
  wire n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470;
  wire n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478;
  wire n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486;
  wire n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494;
  wire n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502;
  wire n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510;
  wire n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518;
  wire n_1519, n_1520, n_1521, n_1522, n_1523, n_1525, n_1526, n_1527;
  wire n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535;
  wire n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543;
  wire n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551;
  wire n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567;
  wire n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575;
  wire n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583;
  wire n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591;
  wire n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599;
  wire n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607;
  wire n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623;
  wire n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632;
  wire n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640;
  wire n_1641, n_1642, n_1643, n_1644, n_1646, n_1647, n_1648, n_1649;
  wire n_1650, n_1651, n_1652, n_1653, n_1654, n_1656, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675;
  wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683;
  wire n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691;
  wire n_1692, n_1693, n_1694, n_1696, n_1697, n_1698, n_1699, n_1700;
  wire n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708;
  wire n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716;
  wire n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724;
  wire n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732;
  wire n_1733, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759;
  wire n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767;
  wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775;
  wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815;
  wire n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  wire n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839;
  wire n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847;
  wire n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855;
  wire n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863;
  wire n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871;
  wire n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879;
  wire n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887;
  wire n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895;
  wire n_1897, n_1898, n_1899, n_1901, n_1902, n_1903, n_1904, n_1905;
  wire n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913;
  wire n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921;
  wire n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929;
  wire n_1930, n_1931, n_1932, n_1933, n_1934, n_1936, n_1937, n_1938;
  wire n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946;
  wire n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954;
  wire n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962;
  wire n_1963, n_1964, n_1965, n_1966, n_1967, n_1971, n_1972, n_1973;
  wire n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981;
  wire n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989;
  wire n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997;
  wire n_1998, n_2000, n_2001, n_2002, n_2004, n_2005, n_2006, n_2007;
  wire n_2008, n_2009, n_2010, n_2011, n_2013, n_2014, n_2015, n_2016;
  wire n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024;
  wire n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032;
  wire n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040;
  wire n_2041, n_2042, n_2043, n_2044, n_2046, n_2047, n_2049, n_2050;
  wire n_2051, n_2052, n_2053, n_2054, n_2055, n_2057, n_2058, n_2059;
  wire n_2060, n_2061, n_2062, n_2063, n_2064, n_2066, n_2067, n_2068;
  wire n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076;
  wire n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084;
  wire n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092;
  wire n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100;
  wire n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108;
  wire n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116;
  wire n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124;
  wire n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132;
  wire n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140;
  wire n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148;
  wire n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157;
  wire n_2158, n_2159, n_2160, n_2162, n_2163, n_2164, n_2165, n_2166;
  wire n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174;
  wire n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182;
  wire n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2191;
  wire n_2193, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201;
  wire n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209;
  wire n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217;
  wire n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225;
  wire n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233;
  wire n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241;
  wire n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249;
  wire n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257;
  wire n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265;
  wire n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273;
  wire n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281;
  wire n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289;
  wire n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297;
  wire n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305;
  wire n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313;
  wire n_2314, n_2315, n_2316, n_2317, n_2319, n_2320, n_2321, n_2322;
  wire n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331;
  wire n_2333, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341;
  wire n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349;
  wire n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357;
  wire n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365;
  wire n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373;
  wire n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381;
  wire n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389;
  wire n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397;
  wire n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405;
  wire n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413;
  wire n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421;
  wire n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429;
  wire n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437;
  wire n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445;
  wire n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453;
  wire n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461;
  wire n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469;
  wire n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477;
  wire n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485;
  wire n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493;
  wire n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501;
  wire n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509;
  wire n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517;
  wire n_2518, n_2519, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526;
  wire n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534;
  wire n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542;
  wire n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550;
  wire n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558;
  wire n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566;
  wire n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574;
  wire n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582;
  wire n_2583, n_2584, n_2588, n_2589, n_2591, n_2592, n_2593, n_2594;
  wire n_2595, n_2597, n_2598, n_2599, n_2601, n_2602, n_2603, n_2604;
  wire n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612;
  wire n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620;
  wire n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628;
  wire n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636;
  wire n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644;
  wire n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652;
  wire n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660;
  wire n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668;
  wire n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676;
  wire n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684;
  wire n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692;
  wire n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700;
  wire n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708;
  wire n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716;
  wire n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724;
  wire n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, n_2732;
  wire n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740;
  wire n_2741, n_2742, n_2743, n_2745, n_2746, n_2747, n_2748, n_2749;
  wire n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757;
  wire n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765;
  wire n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773;
  wire n_2774, n_2775, n_2776, n_2778, n_2779, n_2780, n_2781, n_2782;
  wire n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790;
  wire n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798;
  wire n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806;
  wire n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814;
  wire n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822;
  wire n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2832;
  wire n_2833, n_2834, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841;
  wire n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849;
  wire n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857;
  wire n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865;
  wire n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873;
  wire n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881;
  wire n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889;
  wire n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897;
  wire n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905;
  wire n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913;
  wire n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921;
  wire n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929;
  wire n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937;
  wire n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945;
  wire n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953;
  wire n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961;
  wire n_2962, n_2963, n_2964, n_2966, n_2967, n_2968, n_2969, n_2970;
  wire n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978;
  wire n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986;
  wire n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994;
  wire n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, n_3002;
  wire n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010;
  wire n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018;
  wire n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3026, n_3027;
  wire n_3031, n_3032, n_3033, n_3034, n_3035, n_3037, n_3038, n_3040;
  wire n_3041, n_3043, n_3044, n_3045, n_3046, n_3048, n_3049, n_3050;
  wire n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058;
  wire n_3060, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068;
  wire n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3076, n_3077;
  wire n_3079, n_3081, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088;
  wire n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096;
  wire n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104;
  wire n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112;
  wire n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120;
  wire n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128;
  wire n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136;
  wire n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144;
  wire n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152;
  wire n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160;
  wire n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168;
  wire n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176;
  wire n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184;
  wire n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192;
  wire n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200;
  wire n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208;
  wire n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216;
  wire n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224;
  wire n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232;
  wire n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240;
  wire n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248;
  wire n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256;
  wire n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264;
  wire n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272;
  wire n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280;
  wire n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288;
  wire n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296;
  wire n_3297, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305;
  wire n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313;
  wire n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321;
  wire n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3330;
  wire n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338;
  wire n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346;
  wire n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354;
  wire n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3362, n_3363;
  wire n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, n_3371;
  wire n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379;
  wire n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387;
  wire n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396;
  wire n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404;
  wire n_3405, n_3406, n_3407, n_3408, n_3410, n_3415, n_3418, n_3419;
  wire n_3421, n_3422, n_3423, n_3424, n_3425, n_3427, n_3428, n_3429;
  wire n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437;
  wire n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445;
  wire n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453;
  wire n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461;
  wire n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469;
  wire n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477;
  wire n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485;
  wire n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493;
  wire n_3494, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502;
  wire n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3510;
  wire n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3519;
  wire n_3521, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529;
  wire n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537;
  wire n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545;
  wire n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553;
  wire n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561;
  wire n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569;
  wire n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577;
  wire n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585;
  wire n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593;
  wire n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3601, n_3602;
  wire n_3603, n_3604, n_3605, n_3606, n_3608, n_3609, n_3610, n_3611;
  wire n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619;
  wire n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627;
  wire n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635;
  wire n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643;
  wire n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651;
  wire n_3652, n_3653, n_3654, n_3655, n_3656, n_3658, n_3659, n_3660;
  wire n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668;
  wire n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3677;
  wire n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685;
  wire n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693;
  wire n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701;
  wire n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708, n_3709;
  wire n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, n_3717;
  wire n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725;
  wire n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733;
  wire n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741;
  wire n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, n_3749;
  wire n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757;
  wire n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765;
  wire n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773;
  wire n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781;
  wire n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788, n_3789;
  wire n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797;
  wire n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805;
  wire n_3806, n_3807, n_3808, n_3809, n_3811, n_3812, n_3813, n_3814;
  wire n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822;
  wire n_3823, n_3824, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831;
  wire n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839;
  wire n_3840, n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847;
  wire n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855;
  wire n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863;
  wire n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, n_3871;
  wire n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879;
  wire n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, n_3887, n_3888;
  wire n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896;
  wire n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904;
  wire n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912;
  wire n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920;
  wire n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928;
  wire n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936;
  wire n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944;
  wire n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952;
  wire n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960;
  wire n_3961, n_3962, n_3963, n_3964, n_3966, n_3967, n_3968, n_3969;
  wire n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977;
  wire n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985;
  wire n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993;
  wire n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001;
  wire n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009;
  wire n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, n_4017, n_4018;
  wire n_4019, n_4020, n_4022, n_4024, n_4028, n_4030, n_4031, n_4032;
  wire n_4033, n_4034, n_4035, n_4036, n_4037, n_4039, n_4040, n_4041;
  wire n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049;
  wire n_4050, n_4051, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058;
  wire n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066;
  wire n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074;
  wire n_4075, n_4076, n_4077, n_4078, n_4079, n_4081, n_4082, n_4083;
  wire n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091;
  wire n_4092, n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099;
  wire n_4100, n_4101, n_4102, n_4103, n_4104, n_4105, n_4106, n_4108;
  wire n_4109, n_4110, n_4111, n_4112, n_4113, n_4114, n_4115, n_4116;
  wire n_4117, n_4118, n_4119, n_4120, n_4121, n_4122, n_4123, n_4124;
  wire n_4125, n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132;
  wire n_4133, n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140;
  wire n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148;
  wire n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157;
  wire n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165;
  wire n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173;
  wire n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181;
  wire n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190;
  wire n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198;
  wire n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206;
  wire n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214;
  wire n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222;
  wire n_4223, n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230;
  wire n_4231, n_4232, n_4233, n_4235, n_4236, n_4237, n_4238, n_4239;
  wire n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247;
  wire n_4248, n_4249, n_4250, n_4252, n_4253, n_4254, n_4255, n_4256;
  wire n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264;
  wire n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272;
  wire n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280;
  wire n_4281, n_4282, n_4283, n_4285, n_4286, n_4287, n_4288, n_4289;
  wire n_4290, n_4291, n_4292, n_4293, n_4294, n_4295, n_4296, n_4297;
  wire n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, n_4304, n_4305;
  wire n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313;
  wire n_4314, n_4315, n_4316, n_4317, n_4319, n_4320, n_4321, n_4322;
  wire n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330;
  wire n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338;
  wire n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, n_4346;
  wire n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355;
  wire n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4363, n_4364;
  wire n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372;
  wire n_4373, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381;
  wire n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388, n_4389;
  wire n_4390, n_4391, n_4392, n_4393, n_4394, n_4395, n_4396, n_4397;
  wire n_4398, n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405;
  wire n_4406, n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413;
  wire n_4414, n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, n_4421;
  wire n_4422, n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429;
  wire n_4430, n_4431, n_4432, n_4433, n_4434, n_4435, n_4436, n_4437;
  wire n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445;
  wire n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453;
  wire n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461;
  wire n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4469, n_4470;
  wire n_4471, n_4472, n_4473, n_4474, n_4475, n_4476, n_4477, n_4478;
  wire n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485, n_4486;
  wire n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493, n_4494;
  wire n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501, n_4502;
  wire n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509, n_4510;
  wire n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518;
  wire n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526;
  wire n_4527, n_4528, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535;
  wire n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543;
  wire n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551;
  wire n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559;
  wire n_4560, n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567;
  wire n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575;
  wire n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583;
  wire n_4584, n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591;
  wire n_4592, n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599;
  wire n_4600, n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607;
  wire n_4608, n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615;
  wire n_4616, n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623;
  wire n_4624, n_4625, n_4626, n_4627, n_4628, n_4629, n_4630, n_4631;
  wire n_4632, n_4633, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640;
  wire n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4649;
  wire n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657;
  wire n_4658, n_4660, n_4661, n_4663, n_4664, n_4665, n_4666, n_4667;
  wire n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4675;
  wire n_4676, n_4677, n_4678, n_4679, n_4680, n_4681, n_4682, n_4683;
  wire n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, n_4690, n_4691;
  wire n_4692, n_4693, n_4694, n_4696, n_4698, n_4699, n_4700, n_4701;
  wire n_4703, n_4704, n_4705, n_4706, n_4707, n_4708, n_4709, n_4710;
  wire n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, n_4717, n_4718;
  wire n_4719, n_4720, n_4721, n_4722, n_4723, n_4724, n_4725, n_4726;
  wire n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734;
  wire n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742;
  wire n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750;
  wire n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758;
  wire n_4759, n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766;
  wire n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774;
  wire n_4775, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783;
  wire n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791;
  wire n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799;
  wire n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807;
  wire n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815;
  wire n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823;
  wire n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831;
  wire n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839;
  wire n_4840, n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847;
  wire n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855;
  wire n_4856, n_4857, n_4858, n_4860, n_4861, n_4862, n_4863, n_4864;
  wire n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872;
  wire n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, n_4880;
  wire n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888;
  wire n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4897;
  wire n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905;
  wire n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913;
  wire n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921;
  wire n_4922, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929;
  wire n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937;
  wire n_4940, n_4941, n_4943, n_4944, n_4945, n_4946, n_4947, n_4948;
  wire n_4949, n_4950, n_4951, n_4952, n_4953, n_4954, n_4955, n_4956;
  wire n_4957, n_4958, n_4959, n_4960, n_4961, n_4962, n_4963, n_4964;
  wire n_4965, n_4966, n_4967, n_4968, n_4969, n_4970, n_4971, n_4972;
  wire n_4973, n_4974, n_4975, n_4976, n_4977, n_4978, n_4979, n_4980;
  wire n_4981, n_4982, n_4983, n_4984, n_4985, n_4986, n_4987, n_4988;
  wire n_4989, n_4990, n_4991, n_4992, n_4993, n_4994, n_4995, n_4996;
  wire n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004;
  wire n_5005, n_5006, n_5008, n_5009, n_5010, n_5011, n_5013, n_5014;
  wire n_5015, n_5016, n_5017, n_5018, n_5019, n_5020, n_5021, n_5022;
  wire n_5023, n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031;
  wire n_5032, n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039;
  wire n_5040, n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047;
  wire n_5048, n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055;
  wire n_5056, n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063;
  wire n_5064, n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071;
  wire n_5072, n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079;
  wire n_5080, n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087;
  wire n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095;
  wire n_5096, n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103;
  wire n_5104, n_5105, n_5106, n_5107, n_5108, n_5109, n_5110, n_5111;
  wire n_5112, n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119;
  wire n_5120, n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127;
  wire n_5128, n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135;
  wire n_5136, n_5137, n_5138, n_5139, n_5140, n_5141, n_5142, n_5143;
  wire n_5144, n_5145, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151;
  wire n_5152, n_5153, n_5154, n_5155, n_5156, n_5157, n_5158, n_5159;
  wire n_5160, n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167;
  wire n_5168, n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175;
  wire n_5176, n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183;
  wire n_5184, n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191;
  wire n_5192, n_5193, n_5194, n_5195, n_5196, n_5197, n_5198, n_5199;
  wire n_5200, n_5201, n_5202, n_5203, n_5204, n_5205, n_5206, n_5207;
  wire n_5208, n_5209, n_5210, n_5211, n_5212, n_5213, n_5214, n_5215;
  wire n_5216, n_5217, n_5218, n_5219, n_5220, n_5221, n_5222, n_5223;
  wire n_5224, n_5225, n_5226, n_5227, n_5228, n_5229, n_5230, n_5231;
  wire n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240;
  wire n_5241, n_5242, n_5243, n_5245, n_5246, n_5247, n_5248, n_5249;
  wire n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256, n_5257;
  wire n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5265;
  wire n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272, n_5273;
  wire n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280, n_5281;
  wire n_5283, n_5284, n_5285, n_5286, n_5287, n_5289, n_5290, n_5291;
  wire n_5292, n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299;
  wire n_5300, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307;
  wire n_5308, n_5309, n_5310, n_5311, n_5312, n_5313, n_5314, n_5315;
  wire n_5316, n_5317, n_5323, n_5324, n_5326, n_5327, n_5328, n_5329;
  wire n_5331, n_5332, n_5333, n_5338, n_5340, n_5341, n_5342, n_5343;
  wire n_5344, n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351;
  wire n_5352, n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359;
  wire n_5360, n_5361, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367;
  wire n_5368, n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375;
  wire n_5376, n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383;
  wire n_5384, n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391;
  wire n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399;
  wire n_5400, n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407;
  wire n_5408, n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415;
  wire n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423;
  wire n_5424, n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431;
  wire n_5432, n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439;
  wire n_5440, n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447;
  wire n_5448, n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455;
  wire n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463;
  wire n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471;
  wire n_5472, n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479;
  wire n_5480, n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487;
  wire n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496;
  wire n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504;
  wire n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512;
  wire n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520;
  wire n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528;
  wire n_5529, n_5530, n_5531, n_5533, n_5534, n_5535, n_5536, n_5537;
  wire n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544, n_5545;
  wire n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552, n_5553;
  wire n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560, n_5561;
  wire n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568, n_5569;
  wire n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576, n_5577;
  wire n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584, n_5585;
  wire n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592, n_5593;
  wire n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600, n_5601;
  wire n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608, n_5609;
  wire n_5610, n_5611, n_5612, n_5613, n_5614, n_5615, n_5616, n_5617;
  wire n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5624, n_5625;
  wire n_5626, n_5627, n_5628, n_5629, n_5630, n_5631, n_5632, n_5633;
  wire n_5634, n_5635, n_5636, n_5637, n_5638, n_5639, n_5640, n_5641;
  wire n_5642, n_5643, n_5644, n_5645, n_5646, n_5647, n_5648, n_5649;
  wire n_5650, n_5651, n_5652, n_5653, n_5654, n_5655, n_5656, n_5657;
  wire n_5658, n_5659, n_5660, n_5661, n_5662, n_5663, n_5664, n_5665;
  wire n_5666, n_5667, n_5668, n_5669, n_5670, n_5671, n_5672, n_5673;
  wire n_5674, n_5675, n_5676, n_5677, n_5678, n_5679, n_5680, n_5681;
  wire n_5682, n_5683, n_5684, n_5685, n_5686, n_5687, n_5688, n_5689;
  wire n_5690, n_5691, n_5692, n_5693, n_5694, n_5695, n_5696, n_5697;
  wire n_5698, n_5699, n_5700, n_5701, n_5702, n_5703, n_5704, n_5705;
  wire n_5706, n_5707, n_5708, n_5709, n_5710, n_5711, n_5712, n_5713;
  wire n_5714, n_5715, n_5716, n_5717, n_5718, n_5719, n_5720, n_5721;
  wire n_5722, n_5723, n_5724, n_5725, n_5726, n_5727, n_5728, n_5729;
  wire n_5730, n_5731, n_5732, n_5733, n_5735, n_5736, n_5737, n_5739;
  wire n_5740, n_5741, n_5742, n_5743, n_5744, n_5745, n_5746, n_5747;
  wire n_5748, n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755;
  wire n_5756, n_5757, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763;
  wire n_5764, n_5765, n_5766, n_5767, n_5768, n_5769, n_5770, n_5771;
  wire n_5772, n_5773, n_5774, n_5775, n_5776, n_5777, n_5778, n_5779;
  wire n_5780, n_5781, n_5782, n_5783, n_5784, n_5785, n_5786, n_5787;
  wire n_5788, n_5789, n_5790, n_5791, n_5792, n_5793, n_5794, n_5795;
  wire n_5796, n_5797, n_5798, n_5799, n_5800, n_5801, n_5802, n_5803;
  wire n_5804, n_5805, n_5806, n_5807, n_5808, n_5809, n_5810, n_5811;
  wire n_5812, n_5813, n_5814, n_5815, n_5816, n_5817, n_5818, n_5819;
  wire n_5820, n_5821, n_5822, n_5823, n_5824, n_5825, n_5826, n_5827;
  wire n_5828, n_5829, n_5830, n_5831, n_5832, n_5833, n_5834, n_5835;
  wire n_5836, n_5837, n_5838, n_5839, n_5840, n_5841, n_5842, n_5843;
  wire n_5844, n_5845, n_5847, n_5848, n_5849, n_5851, n_5853, n_5854;
  wire n_5855, n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5864;
  wire n_5865, n_5867, n_5869, n_5870, n_5871, n_5872, n_5873, n_5874;
  wire n_5875, n_5877, n_5878, n_5879, n_5880, n_5881, n_5882, n_5883;
  wire n_5884, n_5885, n_5886, n_5887, n_5888, n_5889, n_5890, n_5891;
  wire n_5892, n_5893, n_5894, n_5895, n_5896, n_5897, n_5898, n_5899;
  wire n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907;
  wire n_5908, n_5909, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915;
  wire n_5916, n_5917, n_5918, n_5920, n_5921, n_5922, n_5923, n_5924;
  wire n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932;
  wire n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940;
  wire n_5941, n_5942, n_5944, n_5945, n_5946, n_5947, n_5948, n_5949;
  wire n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956, n_5957;
  wire n_5958, n_5959, n_5960, n_5961, n_5962, n_5963, n_5965, n_5966;
  wire n_5967, n_5968, n_5969, n_5970, n_5971, n_5972, n_5973, n_5974;
  wire n_5975, n_5976, n_5977, n_5978, n_5979, n_5980, n_5981, n_5982;
  wire n_5983, n_5984, n_5986, n_5987, n_5988, n_5989, n_5990, n_5991;
  wire n_5992, n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999;
  wire n_6000, n_6001, n_6002, n_6003, n_6004, n_6005, n_6007, n_6008;
  wire n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015, n_6016;
  wire n_6017, n_6018, n_6019, n_6020, n_6021, n_6022, n_6023, n_6025;
  wire n_6026, n_6027, n_6028, n_6029, n_6030, n_6031, n_6032, n_6033;
  wire n_6034, n_6035, n_6036, n_6037, n_6038, n_6039, n_6040, n_6041;
  wire n_6042, n_6043, n_6044, n_6045, n_6046, n_6047, n_6048, n_6049;
  wire n_6050, n_6051, n_6052, n_6053, n_6054, n_6058, n_6061, n_6062;
  wire n_6063, n_6064, n_6065, n_6066, n_6067, n_6068, n_6069, n_6070;
  wire n_6071, n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078;
  wire n_6080, n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087;
  wire n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095;
  wire n_6096, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103, n_6104;
  wire n_6105, n_6106, n_6107, n_6108, n_6109, n_6110, n_6111, n_6112;
  wire n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120;
  wire n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128;
  wire n_6129, n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136;
  wire n_6137, n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144;
  wire n_6145, n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6152;
  wire n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6159, n_6160;
  wire n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167, n_6168;
  wire n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175, n_6176;
  wire n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184;
  wire n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192;
  wire n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6203;
  wire n_6212, n_6216, n_6217, n_6218, n_6219, n_6220, n_6221, n_6222;
  wire n_6223, n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230;
  wire n_6231, n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238;
  wire n_6239, n_6240, n_6241, n_6242, n_6243, n_6244, n_6245, n_6246;
  wire n_6247, n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254;
  wire n_6255, n_6256, n_6257, n_6258, n_6259, n_6260, n_6261, n_6262;
  wire n_6263, n_6264, n_6265, n_6266, n_6267, n_6268, n_6269, n_6270;
  wire n_6271, n_6272, n_6273, n_6274, n_6275, n_6276, n_6277, n_6278;
  wire n_6279, n_6280, n_6281, n_6282, n_6283, n_6284, n_6285, n_6286;
  wire n_6287, n_6288, n_6289, n_6290, n_6291, n_6292, n_6293, n_6294;
  wire n_6295, n_6296, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303;
  wire n_6304, n_6305, n_6306, n_6307, n_6308, n_6309, n_6310, n_6311;
  wire n_6312, n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319;
  wire n_6320, n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327;
  wire n_6328, n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335;
  wire n_6336, n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343;
  wire n_6344, n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351;
  wire n_6352, n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6359;
  wire n_6360, n_6361, n_6362, n_6363, n_6364, n_6365, n_6366, n_6367;
  wire n_6368, n_6369, n_6370, n_6371, n_6372, n_6373, n_6374, n_6375;
  wire n_6376, n_6377, n_6378, n_6379, n_6380, n_6381, n_6382, n_6383;
  wire n_6384, n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391;
  wire n_6392, n_6394, n_6396, n_6397, n_6398, n_6399, n_6400, n_6401;
  wire n_6402, n_6403, n_6404, n_6405, n_6406, n_6407, n_6408, n_6409;
  wire n_6410, n_6411, n_6412, n_6413, n_6414, n_6415, n_6416, n_6417;
  wire n_6419, n_6421, n_6422, n_6423, n_6424, n_6425, n_6426, n_6427;
  wire n_6428, n_6429, n_6430, n_6431, n_6432, n_6433, n_6434, n_6435;
  wire n_6436, n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443;
  wire n_6444, n_6445, n_6446, n_6447, n_6448, n_6449, n_6450, n_6451;
  wire n_6453, n_6454, n_6455, n_6456, n_6457, n_6458, n_6459, n_6460;
  wire n_6461, n_6462, n_6463, n_6464, n_6465, n_6466, n_6467, n_6468;
  wire n_6469, n_6470, n_6471, n_6472, n_6473, n_6474, n_6475, n_6476;
  wire n_6477, n_6478, n_6479, n_6482, n_6483, n_6484, n_6485, n_6486;
  wire n_6487, n_6488, n_6489, n_6490, n_6492, n_6493, n_6494, n_6496;
  wire n_6497, n_6498, n_6499, n_6500, n_6501, n_6502, n_6503, n_6504;
  wire n_6505, n_6506, n_6507, n_6508, n_6509, n_6510, n_6511, n_6512;
  wire n_6513, n_6514, n_6515, n_6516, n_6517, n_6518, n_6519, n_6520;
  wire n_6521, n_6522, n_6523, n_6524, n_6525, n_6526, n_6527, n_6528;
  wire n_6529, n_6530, n_6531, n_6532, n_6533, n_6534, n_6535, n_6536;
  wire n_6537, n_6538, n_6539, n_6540, n_6541, n_6542, n_6543, n_6544;
  wire n_6545, n_6546, n_6547, n_6548, n_6549, n_6550, n_6551, n_6552;
  wire n_6553, n_6554, n_6555, n_6556, n_6557, n_6558, n_6559, n_6560;
  wire n_6561, n_6562, n_6563, n_6564, n_6565, n_6566, n_6567, n_6568;
  wire n_6569, n_6570, n_6571, n_6572, n_6573, n_6574, n_6575, n_6576;
  wire n_6577, n_6578, n_6579, n_6580, n_6581, n_6582, n_6583, n_6584;
  wire n_6585, n_6586, n_6587, n_6588, n_6589, n_6590, n_6591, n_6592;
  wire n_6593, n_6594, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600;
  wire n_6601, n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608;
  wire n_6609, n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616;
  wire n_6617, n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624;
  wire n_6625, n_6626, n_6627, n_6628, n_6629, n_6630, n_6631, n_6632;
  wire n_6633, n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640;
  wire n_6641, n_6642, n_6643, n_6644, n_6645, n_6646, n_6647, n_6648;
  wire n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655, n_6656;
  wire n_6657, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663, n_6664;
  wire n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671, n_6672;
  wire n_6673, n_6674, n_6675, n_6676, n_6677, n_6678, n_6679, n_6680;
  wire n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687, n_6688;
  wire n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695, n_6696;
  wire n_6697, n_6698, n_6699, n_6700, n_6701, n_6702, n_6703, n_6704;
  wire n_6705, n_6706, n_6707, n_6708, n_6709, n_6710, n_6711, n_6712;
  wire n_6713, n_6714, n_6715, n_6716, n_6717, n_6718, n_6719, n_6720;
  wire n_6721, n_6722, n_6723, n_6724, n_6725, n_6726, n_6727, n_6728;
  wire n_6729, n_6730, n_6731, n_6732, n_6733, n_6734, n_6735, n_6736;
  wire n_6737, n_6738, n_6739, n_6740, n_6746, n_6747, n_6748, n_6749;
  wire n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756, n_6757;
  wire n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764, n_6765;
  wire n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772, n_6773;
  wire n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780, n_6781;
  wire n_6782, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788, n_6789;
  wire n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796, n_6797;
  wire n_6798, n_6799, n_6800, n_6801, n_6802, n_6803, n_6804, n_6805;
  wire n_6806, n_6807, n_6808, n_6809, n_6810, n_6811, n_6812, n_6813;
  wire n_6814, n_6815, n_6816, n_6817, n_6818, n_6819, n_6820, n_6821;
  wire n_6822, n_6823, n_6824, n_6825, n_6826, n_6827, n_6828, n_6829;
  wire n_6830, n_6831, n_6832, n_6833, n_6834, n_6835, n_6836, n_6837;
  wire n_6838, n_6839, n_6840, n_6841, n_6843, n_6844, n_6845, n_6846;
  wire n_6847, n_6848, n_6849, n_6850, n_6851, n_6852, n_6853, n_6854;
  wire n_6855, n_6856, n_6857, n_6858, n_6859, n_6860, n_6861, n_6862;
  wire n_6863, n_6864, n_6865, n_6866, n_6868, n_6869, n_6870, n_6871;
  wire n_6872, n_6873, n_6874, n_6875, n_6877, n_6878, n_6879, n_6880;
  wire n_6881, n_6882, n_6883, n_6884, n_6885, n_6886, n_6887, n_6888;
  wire n_6889, n_6890, n_6891, n_6892, n_6893, n_6894, n_6895, n_6896;
  wire n_6897, n_6898, n_6899, n_6900, n_6901, n_6902, n_6903, n_6904;
  wire n_6905, n_6906, n_6907, n_6908, n_6909, n_6910, n_6911, n_6912;
  wire n_6913, n_6914, n_6915, n_6916, n_6917, n_6918, n_6919, n_6920;
  wire n_6921, n_6922, n_6923, n_6924, n_6925, n_6926, n_6927, n_6928;
  wire n_6929, n_6930, n_6931, n_6932, n_6933, n_6935, n_6936, n_6937;
  wire n_6938, n_6939, n_6940, n_6941, n_6942, n_6943, n_6944, n_6946;
  wire n_6947, n_6949, n_6950, n_6954, n_6958, n_6960, n_6961, n_6962;
  wire n_6963, n_6964, n_6965, n_6966, n_6973, n_6974, n_6975, n_6976;
  wire n_6977, n_6978, n_6979, n_6980, n_6981, n_6982, n_6983, n_6984;
  wire n_6985, n_6986, n_6987, n_6988, n_6989, n_6990, n_6991, n_6992;
  wire n_6993, n_6994, n_6995, n_6996, n_6997, n_6998, n_6999, n_7000;
  wire n_7001, n_7002, n_7003, n_7004, n_7005, n_7006, n_7007, n_7008;
  wire n_7009, n_7010, n_7011, n_7012, n_7013, n_7014, n_7015, n_7016;
  wire n_7017, n_7018, n_7019, n_7020, n_7021, n_7022, n_7023, n_7024;
  wire n_7025, n_7026, n_7027, n_7028, n_7029, n_7030, n_7031, n_7032;
  wire n_7034, n_7035, n_7036, n_7037, n_7038, n_7039, n_7040, n_7041;
  wire n_7042, n_7043, n_7044, n_7045, n_7046, n_7047, n_7048, n_7049;
  wire n_7050, n_7051, n_7052, n_7053, n_7054, n_7055, n_7056, n_7057;
  wire n_7058, n_7059, n_7060, n_7061, n_7062, n_7063, n_7064, n_7065;
  wire n_7066, n_7067, n_7068, n_7069, n_7070, n_7071, n_7072, n_7073;
  wire n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081;
  wire n_7082, n_7083, n_7084, n_7085, n_7086, n_7087, n_7088, n_7089;
  wire n_7090, n_7091, n_7092, n_7093, n_7094, n_7095, n_7096, n_7097;
  wire n_7098, n_7099, n_7100, n_7103, n_7104, n_7105, n_7106, n_7107;
  wire n_7108, n_7109, n_7110, n_7111, n_7112, n_7113, n_7114, n_7115;
  wire n_7116, n_7117, n_7118, n_7119, n_7120, n_7121, n_7122, n_7123;
  wire n_7124, n_7125, n_7126, n_7127, n_7128, n_7129, n_7130, n_7131;
  wire n_7132, n_7133, n_7134, n_7135, n_7136, n_7137, n_7138, n_7142;
  wire n_7143, n_7144, n_7145, n_7146, n_7147, n_7148, n_7149, n_7150;
  wire n_7151, n_7153, n_7154, n_7155, n_7156, n_7157, n_7158, n_7159;
  wire n_7160, n_7161, n_7162, n_7163, n_7164, n_7165, n_7166, n_7167;
  wire n_7168, n_7169, n_7170, n_7171, n_7172, n_7173, n_7174, n_7175;
  wire n_7176, n_7177, n_7178, n_7179, n_7180, n_7181, n_7182, n_7183;
  wire n_7184, n_7185, n_7186, n_7187, n_7188, n_7189, n_7190, n_7191;
  wire n_7192, n_7193, n_7194, n_7195, n_7196, n_7197, n_7198, n_7199;
  wire n_7200, n_7201, n_7202, n_7203, n_7204, n_7205, n_7206, n_7208;
  wire n_7215, n_7216, n_7217, n_7218, n_7219, n_7221, n_7222, n_7223;
  wire n_7224, n_7225, n_7227, n_7228, n_7229, n_7230, n_7231, n_7232;
  wire n_7233, n_7234, n_7235, n_7236, n_7237, n_7238, n_7239, n_7241;
  wire n_7242, n_7243, n_7244, n_7245, n_7246, n_7247, n_7248, n_7249;
  wire n_7250, n_7251, n_7252, n_7253, n_7254, n_7255, n_7256, n_7257;
  wire n_7258, n_7259, n_7260, n_7261, n_7262, n_7263, n_7264, n_7265;
  wire n_7266, n_7267, n_7268, n_7269, n_7270, n_7271, n_7272, n_7273;
  wire n_7274, n_7275, n_7276, n_7277, n_7278, n_7279, n_7280, n_7281;
  wire n_7282, n_7283, n_7284, n_7285, n_7286, n_7287, n_7288, n_7289;
  wire n_7290, n_7291, n_7292, n_7293, n_7295, n_7297, n_7298, n_7299;
  wire n_7300, n_7301, n_7302, n_7303, n_7304, n_7305, n_7306, n_7307;
  wire n_7308, n_7309, n_7310, n_7311, n_7312, n_7313, n_7314, n_7315;
  wire n_7316, n_7317, n_7318, n_7319, n_7320, n_7321, n_7322, n_7323;
  wire n_7324, n_7325, n_7326, n_7327, n_7328, n_7329, n_7330, n_7331;
  wire n_7332, n_7333, n_7334, n_7335, n_7336, n_7337, n_7338, n_7339;
  wire n_7340, n_7341, n_7342, n_7343, n_7344, n_7345, n_7346, n_7347;
  wire n_7348, n_7349, n_7350, n_7351, n_7352, n_7353, n_7354, n_7355;
  wire n_7356, n_7362, n_7363, n_7364, n_7365, n_7366, n_7367, n_7368;
  wire n_7369, n_7370, n_7371, n_7372, n_7373, n_7374, n_7375, n_7376;
  wire n_7377, n_7378, n_7379, n_7380, n_7381, n_7382, n_7383, n_7384;
  wire n_7385, n_7386, n_7387, n_7388, n_7389, n_7390, n_7391, n_7392;
  wire n_7393, n_7394, n_7395, n_7396, n_7397, n_7398, n_7399, n_7400;
  wire n_7401, n_7402, n_7403, n_7404, n_7407, n_7408, n_7409, n_7410;
  wire n_7411, n_7412, n_7413, n_7414, n_7415, n_7416, n_7417, n_7418;
  wire n_7419, n_7420, n_7421, n_7422, n_7423, n_7424, n_7425, n_7427;
  wire n_7428, n_7429, n_7430, n_7431, n_7432, n_7433, n_7434, n_7435;
  wire n_7436, n_7437, n_7438, n_7439, n_7440, n_7441, n_7442, n_7443;
  wire n_7444, n_7445, n_7446, n_7447, n_7448, n_7449, n_7450, n_7451;
  wire n_7452, n_7453, n_7454, n_7455, n_7457, n_7458, n_7459, n_7460;
  wire n_7461, n_7462, n_7463, n_7464, n_7465, n_7466, n_7467, n_7468;
  wire n_7469, n_7470, n_7471, n_7472, n_7473, n_7474, n_7475, n_7476;
  wire n_7477, n_7478, n_7479, n_7480, n_7481, n_7482, n_7483, n_7484;
  wire n_7485, n_7486, n_7487, n_7489, n_7490, n_7491, n_7493, n_7494;
  wire n_7495, n_7496, n_7497, n_7498, n_7499, n_7500, n_7501, n_7502;
  wire n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509, n_7510;
  wire n_7511, n_7512, n_7513, n_7514, n_7515, n_7516, n_7517, n_7518;
  wire n_7519, n_7520, n_7521, n_7522, n_7523, n_7524, n_7525, n_7527;
  wire n_7528, n_7529, n_7530, n_7531, n_7532, n_7533, n_7534, n_7535;
  wire n_7536, n_7537, n_7538, n_7539, n_7540, n_7541, n_7542, n_7543;
  wire n_7544, n_7545, n_7546, n_7547, n_7548, n_7549, n_7550, n_7552;
  wire n_7555, n_7556, n_7557, n_7558, n_7560, n_7561, n_7563, n_7564;
  wire n_7565, n_7566, n_7568, n_7569, n_7570, n_7571, n_7572, n_7574;
  wire n_7575, n_7576, n_7577, n_7578, n_7579, n_7580, n_7581, n_7582;
  wire n_7583, n_7584, n_7585, n_7586, n_7587, n_7588, n_7589, n_7590;
  wire n_7591, n_7592, n_7593, n_7594, n_7595, n_7597, n_7598, n_7599;
  wire n_7600, n_7601, n_7602, n_7603, n_7604, n_7606, n_7607, n_7608;
  wire n_7609, n_7611, n_7612, n_7613, n_7614, n_7615, n_7616, n_7617;
  wire n_7618, n_7619, n_7620, n_7621, n_7622, n_7623, n_7624, n_7625;
  wire n_7626, n_7627, n_7628, n_7629, n_7630, n_7632, n_7633, n_7634;
  wire n_7635, n_7636, n_7637, n_7638, n_7639, n_7640, n_7641, n_7642;
  wire n_7643, n_7644, n_7645, n_7646, n_7647, n_7648, n_7649, n_7650;
  wire n_7651, n_7652, n_7654, n_7655, n_7656, n_7657, n_7658, n_7659;
  wire n_7660, n_7661, n_7662, n_7663, n_7665, n_7666, n_7667, n_7668;
  wire n_7669, n_7670, n_7671, n_7672, n_7673, n_7674, n_7676, n_7677;
  wire n_7678, n_7679, n_7680, n_7681, n_7682, n_7683, n_7684, n_7685;
  wire n_7686, n_7687, n_7688, n_7689, n_7690, n_7691, n_7692, n_7693;
  wire n_7694, n_7695, n_7697, n_7699, n_7700, n_7701, n_7702, n_7703;
  wire n_7704, n_7705, n_7706, n_7707, n_7708, n_7710, n_7711, n_7712;
  wire n_7713, n_7714, n_7715, n_7716, n_7717, n_7719, n_7720, n_7721;
  wire n_7722, n_7723, n_7724, n_7725, n_7726, n_7727, n_7728, n_7729;
  wire n_7730, n_7731, n_7732, n_7733, n_7734, n_7735, n_7737, n_7738;
  wire n_7740, n_7741, n_7742, n_7743, n_7744, n_7745, n_7746, n_7747;
  wire n_7748, n_7749, n_7750, n_7751, n_7752, n_7755, n_7756, n_7757;
  wire n_7758, n_7759, n_7760, n_7761, n_7762, n_7763, n_7764, n_7765;
  wire n_7766, n_7767, n_7768, n_7769, n_7770, n_7771, n_7772, n_7773;
  wire n_7774, n_7775, n_7776, n_7777, n_7778, n_7779, n_7780, n_7781;
  wire n_7782, n_7783, n_7785, n_7786, n_7787, n_7788, n_7789, n_7791;
  wire n_7792, n_7793, n_7794, n_7795, n_7796, n_7797, n_7798, n_7799;
  wire n_7800, n_7801, n_7802, n_7803, n_7804, n_7805, n_7808, n_7809;
  wire n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816, n_7817;
  wire n_7818, n_7819, n_7820, n_7821, n_7822, n_7823, n_7824, n_7825;
  wire n_7826, n_7828, n_7829, n_7830, n_7831, n_7832, n_7833, n_7834;
  wire n_7835, n_7836, n_7837, n_7838, n_7839, n_7840, n_7841, n_7842;
  wire n_7843, n_7844, n_7845, n_7846, n_7847, n_7848, n_7849, n_7850;
  wire n_7851, n_7852, n_7853, n_7855, n_7856, n_7857, n_7858, n_7860;
  wire n_7861, n_7862, n_7864, n_7865, n_7866, n_7867, n_7868, n_7869;
  wire n_7870, n_7871, n_7872, n_7873, n_7874, n_7875, n_7876, n_7877;
  wire n_7878, n_7879, n_7881, n_7882, n_7883, n_7884, n_7885, n_7886;
  wire n_7887, n_7888, n_7889, n_7890, n_7891, n_7892, n_7893, n_7894;
  wire n_7895, n_7897, n_7898, n_7900, n_7901, n_7902, n_7903, n_7904;
  wire n_7905, n_7906, n_7907, n_7909, n_7910, n_7911, n_7912, n_7913;
  wire n_7914, n_7915, n_7916, n_7917, n_7918, n_7919, n_7920, n_7921;
  wire n_7922, n_7923, n_7924, n_7925, n_7926, n_7927, n_7928, n_7930;
  wire n_7932, n_7933, n_7935, n_7936, n_7937, n_7938, n_7939, n_7940;
  wire n_7941, n_7942, n_7943, n_7944, n_7946, n_7947, n_7950, n_7952;
  wire n_7953, n_7954, n_7955, n_7956, n_7957, n_7958, n_7959, n_7960;
  wire n_7962, n_7963, n_7964, n_7965, n_7966, n_7967, n_7968, n_7970;
  wire n_7971, n_7972, n_7973, n_7974, n_7977, n_7978, n_7979, n_7980;
  wire n_7981, n_7984, n_7985, n_7986, n_7987, n_7988, n_7989, n_7990;
  wire n_7991, n_7992, n_7993, n_7994, n_7995, n_7996, n_7997, n_7998;
  wire n_7999, n_8000, n_8001, n_8003, n_8004, n_8005, n_8007, n_8008;
  wire n_8009, n_8010, n_8011, n_8012, n_8013, n_8014, n_8015, n_8016;
  wire n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8023, n_8025;
  wire n_8026, n_8027, n_8029, n_8031, n_8032, n_8033, n_8034, n_8035;
  wire n_8036, n_8037, n_8038, n_8039, n_8040, n_8041, n_8042, n_8043;
  wire n_8044, n_8046, n_8048, n_8049, n_8050, n_8051, n_8052, n_8053;
  wire n_8054, n_8056, n_8057, n_8058, n_8059, n_8060, n_8061, n_8062;
  wire n_8066, n_8067, n_8068, n_8069, n_8070, n_8071, n_8072, n_8073;
  wire n_8074, n_8075, n_8076, n_8077, n_8078, n_8079, n_8080, n_8081;
  wire n_8082, n_8083, n_8084, n_8085, n_8086, n_8088, n_8089, n_8090;
  wire n_8091, n_8092, n_8093, n_8094, n_8096, n_8098, n_8099, n_8100;
  wire n_8101, n_8105, n_8106, n_8107, n_8108, n_8109, n_8110, n_8111;
  wire n_8112, n_8113, n_8114, n_8115, n_8116, n_8117, n_8118, n_8119;
  wire n_8120, n_8121, n_8122, n_8123, n_8124, n_8125, n_8126, n_8127;
  wire n_8128, n_8129, n_8130, n_8131, n_8132, n_8133, n_8134, n_8135;
  wire n_8136, n_8137, n_8138, n_8139, n_8140, n_8141, n_8142, n_8144;
  wire n_8145, n_8146, n_8147, n_8148, n_8151, n_8152, n_8153, n_8154;
  wire n_8155, n_8156, n_8157, n_8158, n_8159, n_8160, n_8161, n_8162;
  wire n_8163, n_8164, n_8165, n_8166, n_8167, n_8168, n_8169, n_8170;
  wire n_8171, n_8174, n_8175, n_8177, n_8178, n_8179, n_8180, n_8181;
  wire n_8182, n_8183, n_8184, n_8185, n_8186, n_8187, n_8190, n_8192;
  wire n_8193, n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200;
  wire n_8202, n_8204, n_8205, n_8206, n_8207, n_8208, n_8209, n_8210;
  wire n_8211, n_8212, n_8213, n_8214, n_8215, n_8216, n_8217, n_8218;
  wire n_8219, n_8220, n_8221, n_8222, n_8223, n_8225, n_8226, n_8227;
  wire n_8228, n_8229, n_8230, n_8233, n_8234, n_8235, n_8236, n_8237;
  wire n_8239, n_8240, n_8241, n_8242, n_8243, n_8244, n_8245, n_8246;
  wire n_8247, n_8251, n_8252, n_8253, n_8254, n_8255, n_8257, n_8258;
  wire n_8259, n_8260, n_8261, n_8262, n_8263, n_8264, n_8265, n_8266;
  wire n_8267, n_8268, n_8269, n_8270, n_8271, n_8272, n_8273, n_8274;
  wire n_8275, n_8276, n_8277, n_8278, n_8279, n_8280, n_8281, n_8282;
  wire n_8283, n_8284, n_8285, n_8286, n_8288, n_8289, n_8290, n_8291;
  wire n_8292, n_8293, n_8294, n_8295, n_8296, n_8297, n_8299, n_8300;
  wire n_8301, n_8302, n_8303, n_8304, n_8305, n_8306, n_8307, n_8308;
  wire n_8309, n_8310, n_8311, n_8312, n_8313, n_8314, n_8315, n_8316;
  wire n_8317, n_8318, n_8319, n_8320, n_8321, n_8322, n_8323, n_8324;
  wire n_8325, n_8326, n_8327, n_8329, n_8330, n_8331, n_8332, n_8333;
  wire n_8335, n_8336, n_8337, n_8338, n_8339, n_8340, n_8341, n_8342;
  wire n_8343, n_8344, n_8345, n_8346, n_8347, n_8348, n_8349, n_8350;
  wire n_8351, n_8352, n_8353, n_8354, n_8355, n_8356, n_8357, n_8358;
  wire n_8359, n_8360, n_8361, n_8362, n_8363, n_8364, n_8365, n_8366;
  wire n_8367, n_8368, n_8369, n_8370, n_8371, n_8372, n_8373, n_8374;
  wire n_8375, n_8376, n_8377, n_8378, n_8379, n_8380, n_8381, n_8382;
  wire n_8383, n_8384, n_8385, n_8386, n_8387, n_8388, n_8389, n_8391;
  wire n_8392, n_8393, n_8394, n_8395, n_8396, n_8397, n_8398, n_8399;
  wire n_8400, n_8401, n_8402, n_8403, n_8405, n_8406, n_8407, n_8408;
  wire n_8409, n_8410, n_8411, n_8412, n_8413, n_8414, n_8415, n_8416;
  wire n_8417, n_8418, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424;
  wire n_8425, n_8426, n_8427, n_8428, n_8429, n_8430, n_8431, n_8432;
  wire n_8433, n_8434, n_8435, n_8436, n_8437, n_8438, n_8439, n_8440;
  wire n_8441, n_8442, n_8443, n_8444, n_8445, n_8446, n_8447, n_8448;
  wire n_8449, n_8450, n_8451, n_8452, n_8453, n_8454, n_8455, n_8456;
  wire n_8457, n_8458, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464;
  wire n_8465, n_8466, n_8467, n_8468, n_8469, n_8470, n_8471, n_8472;
  wire n_8473, n_8474, n_8475, n_8476, n_8477, n_8479, n_8480, n_8481;
  wire n_8482, n_8483, n_8484, n_8485, n_8486, n_8487, n_8488, n_8489;
  wire n_8490, n_8491, n_8492, n_8493, n_8494, n_8495, n_8496, n_8497;
  wire n_8498, n_8499, n_8500, n_8501, n_8504, n_8505, n_8506, n_8508;
  wire n_8509, n_8510, n_8511, n_8512, n_8513, n_8514, n_8515, n_8516;
  wire n_8517, n_8518, n_8519, n_8520, n_8521, n_8522, n_8523, n_8524;
  wire n_8525, n_8526, n_8527, n_8528, n_8529, n_8530, n_8531, n_8532;
  wire n_8533, n_8535, n_8536, n_8538, n_8540, n_8541, n_8542, n_8543;
  wire n_8544, n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551;
  wire n_8552, n_8553, n_8554, n_8555, n_8556, n_8557, n_8558, n_8559;
  wire n_8560, n_8561, n_8562, n_8563, n_8564, n_8565, n_8566, n_8567;
  wire n_8568, n_8569, n_8570, n_8571, n_8572, n_8573, n_8574, n_8575;
  wire n_8576, n_8577, n_8578, n_8579, n_8580, n_8581, n_8582, n_8583;
  wire n_8584, n_8585, n_8586, n_8587, n_8588, n_8589, n_8590, n_8591;
  wire n_8592, n_8593, n_8594, n_8595, n_8596, n_8597, n_8598, n_8599;
  wire n_8600, n_8601, n_8602, n_8603, n_8604, n_8605, n_8606, n_8607;
  wire n_8608, n_8609, n_8610, n_8612, n_8614, n_8616, n_8617, n_8618;
  wire n_8619, n_8620, n_8621, n_8622, n_8626, n_8627, n_8628, n_8629;
  wire n_8630, n_8631, n_8632, n_8633, n_8634, n_8635, n_8636, n_8637;
  wire n_8638, n_8639, n_8640, n_8641, n_8642, n_8643, n_8644, n_8645;
  wire n_8646, n_8647, n_8648, n_8649, n_8650, n_8651, n_8652, n_8653;
  wire n_8654, n_8655, n_8657, n_8658, n_8659, n_8660, n_8661, n_8662;
  wire n_8663, n_8664, n_8665, n_8666, n_8667, n_8668, n_8669, n_8670;
  wire n_8671, n_8672, n_8673, n_8674, n_8675, n_8676, n_8677, n_8678;
  wire n_8679, n_8680, n_8681, n_8682, n_8683, n_8684, n_8685, n_8686;
  wire n_8687, n_8688, n_8689, n_8690, n_8691, n_8692, n_8693, n_8694;
  wire n_8695, n_8696, n_8698, n_8699, n_8700, n_8701, n_8702, n_8703;
  wire n_8704, n_8705, n_8706, n_8707, n_8708, n_8709, n_8710, n_8711;
  wire n_8712, n_8713, n_8714, n_8715, n_8716, n_8717, n_8718, n_8719;
  wire n_8720, n_8721, n_8722, n_8723, n_8724, n_8725, n_8726, n_8727;
  wire n_8728, n_8729, n_8730, n_8731, n_8732, n_8733, n_8734, n_8735;
  wire n_8739, n_8740, n_8741, n_8742, n_8743, n_8744, n_8745, n_8746;
  wire n_8747, n_8748, n_8749, n_8750, n_8751, n_8752, n_8753, n_8754;
  wire n_8755, n_8756, n_8757, n_8758, n_8759, n_8760, n_8761, n_8762;
  wire n_8763, n_8764, n_8765, n_8766, n_8767, n_8768, n_8769, n_8770;
  wire n_8771, n_8772, n_8773, n_8774, n_8775, n_8776, n_8777, n_8778;
  wire n_8779, n_8780, n_8781, n_8782, n_8783, n_8784, n_8785, n_8786;
  wire n_8787, n_8788, n_8789, n_8790, n_8791, n_8792, n_8793, n_8794;
  wire n_8795, n_8796, n_8797, n_8798, n_8799, n_8800, n_8801, n_8802;
  wire n_8803, n_8804, n_8805, n_8806, n_8807, n_8808, n_8809, n_8810;
  wire n_8811, n_8812, n_8813, n_8814, n_8815, n_8816, n_8817, n_8818;
  wire n_8819, n_8820, n_8821, n_8822, n_8823, n_8824, n_8825, n_8826;
  wire n_8827, n_8828, n_8829, n_8830, n_8831, n_8832, n_8833, n_8834;
  wire n_8835, n_8836, n_8837, n_8838, n_8839, n_8840, n_8841, n_8845;
  wire n_8846, n_8847, n_8848, n_8849, n_8850, n_8851, n_8852, n_8853;
  wire n_8854, n_8855, n_8856, n_8857, n_8858, n_8859, n_8860, n_8861;
  wire n_8862, n_8863, n_8864, n_8865, n_8866, n_8867, n_8868, n_8869;
  wire n_8870, n_8871, n_8872, n_8873, n_8874, n_8875, n_8876, n_8878;
  wire n_8880, n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888;
  wire n_8889, n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896;
  wire n_8897, n_8898, n_8899, n_8900, n_8901, n_8902, n_8903, n_8904;
  wire n_8905, n_8906, n_8907, n_8908, n_8909, n_8910, n_8911, n_8912;
  wire n_8913, n_8914, n_8915, n_8916, n_8917, n_8918, n_8919, n_8920;
  wire n_8921, n_8922, n_8923, n_8924, n_8925, n_8926, n_8927, n_8928;
  wire n_8929, n_8930, n_8931, n_8932, n_8933, n_8934, n_8935, n_8936;
  wire n_8937, n_8938, n_8939, n_8941, n_8942, n_8943, n_8944, n_8945;
  wire n_8946, n_8947, n_8948, n_8950, n_8951, n_8952, n_8953, n_8954;
  wire n_8955, n_8956, n_8957, n_8958, n_8960, n_8961, n_8962, n_8963;
  wire n_8964, n_8965, n_8966, n_8967, n_8968, n_8969, n_8970, n_8971;
  wire n_8972, n_8973, n_8974, n_8975, n_8976, n_8977, n_8978, n_8979;
  wire n_8980, n_8981, n_8982, n_8983, n_8984, n_8985, n_8986, n_8988;
  wire n_8989, n_8990, n_8991, n_8992, n_8993, n_8995, n_8997, n_8999;
  wire n_9000, n_9001, n_9002, n_9004, n_9005, n_9006, n_9007, n_9008;
  wire n_9009, n_9010, n_9011, n_9012, n_9013, n_9014, n_9015, n_9016;
  wire n_9017, n_9018, n_9019, n_9020, n_9021, n_9022, n_9023, n_9024;
  wire n_9025, n_9026, n_9027, n_9029, n_9030, n_9031, n_9032, n_9033;
  wire n_9034, n_9035, n_9036, n_9038, n_9042, n_9044, n_9045, n_9046;
  wire n_9047, n_9048, n_9049, n_9050, n_9051, n_9052, n_9053, n_9054;
  wire n_9055, n_9056, n_9057, n_9058, n_9059, n_9062, n_9063, n_9064;
  wire n_9065, n_9066, n_9067, n_9068, n_9069, n_9070, n_9071, n_9072;
  wire n_9073, n_9075, n_9076, n_9077, n_9078, n_9079, n_9080, n_9081;
  wire n_9082, n_9084, n_9085, n_9086, n_9087, n_9088, n_9089, n_9090;
  wire n_9091, n_9092, n_9093, n_9094, n_9095, n_9096, n_9097, n_9098;
  wire n_9099, n_9100, n_9101, n_9102, n_9103, n_9104, n_9105, n_9106;
  wire n_9107, n_9108, n_9109, n_9110, n_9111, n_9112, n_9113, n_9114;
  wire n_9115, n_9116, n_9117, n_9118, n_9119, n_9120, n_9121, n_9122;
  wire n_9123, n_9124, n_9125, n_9126, n_9127, n_9128, n_9129, n_9130;
  wire n_9131, n_9132, n_9133, n_9134, n_9135, n_9136, n_9137, n_9138;
  wire n_9139, n_9141, n_9145, n_9147, n_9148, n_9149, n_9150, n_9151;
  wire n_9152, n_9153, n_9154, n_9155, n_9156, n_9157, n_9158, n_9159;
  wire n_9160, n_9161, n_9162, n_9163, n_9164, n_9165, n_9166, n_9167;
  wire n_9168, n_9169, n_9170, n_9171, n_9172, n_9173, n_9174, n_9175;
  wire n_9176, n_9177, n_9181, n_9183, n_9185, n_9186, n_9187, n_9188;
  wire n_9189, n_9190, n_9191, n_9192, n_9193, n_9194, n_9195, n_9196;
  wire n_9197, n_9199, n_9203, n_9205, n_9206, n_9207, n_9208, n_9209;
  wire n_9210, n_9211, n_9212, n_9213, n_9214, n_9215, n_9216, n_9217;
  wire n_9218, n_9219, n_9220, n_9223, n_9227, n_9228, n_9229, n_9230;
  wire n_9231, n_9232, n_9233, n_9234, n_9235, n_9236, n_9237, n_9238;
  wire n_9239, n_9240, n_9241, n_9242, n_9243, n_9244, n_9245, n_9246;
  wire n_9247, n_9248, n_9249, n_9250, n_9251, n_9252, n_9253, n_9254;
  wire n_9255, n_9256, n_9257, n_9258, n_9259, n_9260, n_9261, n_9262;
  wire n_9263, n_9264, n_9265, n_9266, n_9267, n_9270, n_9271, n_9272;
  wire n_9273, n_9274, n_9275, n_9276, n_9277, n_9278, n_9279, n_9280;
  wire n_9281, n_9282, n_9283, n_9284, n_9285, n_9286, n_9287, n_9288;
  wire n_9289, n_9290, n_9291, n_9292, n_9293, n_9295, n_9296, n_10109;
  wire n_10110, n_10111, n_10112, n_10113, n_10114, n_10115, n_10116,
       n_10117;
  wire n_10118, n_10119, n_10120, n_10121, n_10122, n_10123, n_10124,
       n_10125;
  wire n_10126, n_10127, n_10128, n_10129, n_10131, n_10133, n_10134,
       n_10135;
  wire n_10137, n_10138, n_10141, n_10142, n_10143, n_10144, n_10145,
       n_10146;
  wire n_10147, n_10148, n_10149, n_10150, n_10151, n_10152, n_10153,
       n_10154;
  wire n_10155, n_10156, n_10157, n_10158, n_10159, n_10160, n_10161,
       n_10162;
  wire n_10163, n_10164, n_10165, n_10167, n_10169, n_10171, n_10173,
       n_10175;
  wire n_10177, n_10179, n_10181, n_10183, n_10185, n_10186, n_10187,
       n_10188;
  wire n_10189, n_10190, n_10191, n_10192, n_10193, n_10194, n_10195,
       n_10196;
  wire n_10197, n_10198, n_10199, n_10200, n_10201, n_10202, n_10203,
       n_10204;
  wire n_10205, n_10206, n_10207, n_10208, n_10209, n_10211, n_10212,
       n_10213;
  wire n_10215, n_10216, n_10217, n_10218, n_10219, n_10220, n_10221,
       n_10222;
  wire n_10223, n_10227, n_10228, n_10229, n_10231, n_10232, n_10233,
       n_10235;
  wire n_10237, n_10238, n_10239, n_10240, n_10241, n_10242, n_10243,
       n_10244;
  wire n_10245, n_10247, n_10249, n_10250, n_10251, n_10252, n_10253,
       n_10254;
  wire n_10255, n_10256, n_10257, n_10258, n_10260, n_10261, n_10262,
       n_10264;
  wire n_10265, n_10267, n_10268, n_10270, n_10271, n_10273, n_10274,
       n_10276;
  wire n_10277, n_10279, n_10280, n_10282, n_10283, n_10285, n_10286,
       n_10287;
  wire n_10288, n_10289, n_10290, n_10291, n_10292, n_10294, n_10295,
       n_10296;
  wire n_10297, n_10298, n_10299, n_10300, n_10301, n_10302, n_10303,
       n_10304;
  wire n_10305, n_10306, n_10307, n_10308, n_10309, n_10310, n_10311,
       n_10312;
  wire n_10313, n_10314, n_10316, n_10317, n_10318, n_10319, n_10320,
       n_10321;
  wire n_10322, n_10323, n_10325, n_10326, n_10327, n_10328, n_10329,
       n_10331;
  wire n_10332, n_10334, n_10335, n_10336, n_10337, n_10338, n_10339,
       n_10340;
  wire n_10341, n_10342, n_10343, n_10344, n_10346, n_10347, n_10349,
       n_10350;
  wire n_10351, n_10352, n_10353, n_10354, n_10355, n_10356, n_10357,
       n_10358;
  wire n_10359, n_10360, n_10361, n_10362, n_10363, n_10364, n_10365,
       n_10366;
  wire n_10367, n_10368, n_10369, n_10370, n_10371, n_10373, n_10374,
       n_10375;
  wire n_10376, n_10377, n_10378, n_10379, n_10380, n_10381, n_10382,
       n_10383;
  wire n_10384, n_10386, n_10387, n_10388, n_10389, n_10390, n_10391,
       n_10392;
  wire n_10393, n_10394, n_10395, n_10396, n_10397, n_10398, n_10399,
       n_10400;
  wire n_10401, n_10402, n_10403, n_10404, n_10405, n_10406, n_10407,
       n_10408;
  wire n_10409, n_10410, n_10411, n_10412, n_10413, n_10414, n_10415,
       n_10416;
  wire n_10417, n_10418, n_10419, n_10420, n_10421, n_10422, n_10423,
       n_10424;
  wire n_10425, n_10426, n_10427, n_10428, n_10429, n_10430, n_10431,
       n_10432;
  wire n_10433, n_10434, n_10435, n_10436, n_10437, n_10438, n_10439,
       n_10440;
  wire n_10441, n_10442, n_10443, n_10444, n_10445, n_10446, n_10447,
       n_10448;
  wire n_10449, n_10450, n_10451, n_10452, n_10453, new_g6821_,
       new_g6832_, new_g6856_;
  wire new_g6875_, new_g6888_, new_g6905_, new_g6928_, new_g6946_,
       new_g6961_, new_g7004_, new_g7028_;
  wire new_g7051_, new_g7074_, new_g7097_, new_g7121_, new_g7558_,
       new_g7586_, new_g7704_, new_g7717_;
  wire new_g7738_, new_g7753_, new_g7766_, new_g7791_, new_g7812_,
       new_g8038_, new_g8703_, new_g8880_;
  wire new_g10233_, new_g10295_, new_g10323_, new_g10354_, new_g10366_,
       new_g10371_, new_g10375_, new_g10383_;
  wire new_g10401_, new_g10405_, new_g10409_, new_g10413_, new_g10795_,
       new_g12440_, new_g12875_;
  assign g34972 = 1'b1;
  assign g34956 = g34839;
  assign g34927 = 1'b1;
  assign g34925 = 1'b1;
  assign g34923 = 1'b1;
  assign g34921 = 1'b1;
  assign g34919 = 1'b1;
  assign g34917 = 1'b1;
  assign g34915 = 1'b1;
  assign g34913 = 1'b1;
  assign g34788 = g33894;
  assign g34597 = 1'b0;
  assign g34437 = 1'b1;
  assign g34436 = 1'b1;
  assign g34435 = g31521;
  assign g34425 = 1'b1;
  assign g34383 = 1'b1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g34221 = 1'b1;
  assign g34201 = 1'b1;
  assign g33959 = g28753;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g33935 = 1'b1;
  assign g33874 = 1'b1;
  assign g33659 = 1'b1;
  assign g33636 = 1'b1;
  assign g33533 = g27831;
  assign g32975 = g26801;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g31863 = g25167;
  assign g31862 = g25259;
  assign g31861 = g25219;
  assign g31860 = g25114;
  assign g31665 = 1'b1;
  assign g31656 = 1'b1;
  assign g30332 = g23683;
  assign g30331 = g23759;
  assign g30330 = g23652;
  assign g30329 = g23612;
  assign g30327 = g23002;
  assign g29221 = g21292;
  assign g29220 = g21245;
  assign g29219 = g20654;
  assign g29218 = g18881;
  assign g29217 = g21270;
  assign g29216 = g21176;
  assign g29215 = g20901;
  assign g29214 = g20652;
  assign g29213 = g20557;
  assign g29212 = g20899;
  assign g29211 = g20763;
  assign g29210 = g20049;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g23190 = 1'b1;
  assign g21698 = g36;
  assign g18101 = g6746;
  assign g18100 = g6751;
  assign g18099 = g6745;
  assign g18098 = g6744;
  assign g18097 = g6747;
  assign g18096 = g6750;
  assign g18095 = g6749;
  assign g18094 = g6748;
  assign g18092 = g6753;
  assign g12368 = 1'b0;
  assign g9048 = 1'b0;
  assign g8403 = 1'b0;
  assign g8353 = 1'b0;
  assign g8283 = 1'b0;
  assign g8235 = 1'b0;
  assign g8178 = 1'b0;
  assign g8132 = 1'b0;
  fflopd g2955_reg(.CK (clock), .D (n_9296), .Q (g2955));
  nand g173601__2398 (n_9296, n_1169, n_9295);
  nand g173603__5107 (n_9295, g35, n_9293);
  nand g173602__6260 (g31793, n_9285, n_9292);
  nand g173604__4319 (n_9293, n_631, n_9291);
  nor g173605__8428 (n_9292, n_9282, n_9290);
  nor g173607__5526 (n_9291, g2946, n_9287);
  nand g173608__6783 (n_9290, n_9283, n_9289);
  fflopd g2864_reg(.CK (clock), .D (n_9288), .Q (g2864));
  nand g173611__3680 (n_9289, n_2876, n_9284);
  nand g173609__1617 (n_9288, n_2059, n_9286);
  nand g173610__2802 (n_9287, n_9286, n_7048);
  nor g173612__1705 (n_9286, n_3320, n_9285);
  nand g173613__5122 (n_9284, n_9273, n_9281);
  nand g173615__8246 (n_9283, n_1967, n_9280);
  nor g173614__7098 (n_9282, n_1966, n_9279);
  nand g173616__6131 (n_9281, n_487, n_9276);
  not g173618 (n_9280, n_9278);
  nand g173617__1881 (n_9285, n_3736, n_9275);
  nand g173619__5115 (n_9279, n_1699, n_9277);
  nand g173620__7482 (n_9278, n_1698, n_9277);
  nand g173622__4733 (n_9276, n_9274, n_9272);
  nor g173621__6161 (n_9275, n_2875, n_9274);
  nor g173625__9315 (n_9277, n_9270, n_9273);
  nand g173623__9945 (n_9274, n_9271, n_2878);
  nand g173624__2883 (n_9272, n_9271, n_4068);
  not g173626 (n_9270, n_9271);
  nand g173627__2346 (n_9271, g35, n_10110);
  fflopd g4420_reg(.CK (clock), .D (n_9267), .Q (g4420));
  wire w, w0, w1, w2;
  nand g173631__7410 (n_9267, w0, w2);
  nand g5 (w2, w1, g4534);
  not g1 (w1, n_4105);
  nand g0 (w0, w, n_4105);
  not g (w, g4534);
  fflopd g4534_reg(.CK (clock), .D (n_9266), .Q (g4534));
  nand g173633__6417 (n_9266, n_1845, n_9265);
  nand g173634__5477 (n_9265, g4564, n_9264);
  fflopd g4564_reg(.CK (clock), .D (n_9263), .Q (g4564));
  nand g173636__2398 (n_9264, g35, n_9262);
  nand g173637__5107 (n_9263, n_1773, n_9261);
  nand g173638__6260 (n_9262, g4561, n_9259);
  nand g173639__4319 (n_9261, g4561, n_9257);
  fflopd g4561_reg(.CK (clock), .D (n_9260), .Q (g4561));
  nand g173641__8428 (n_9260, n_1775, n_9258);
  not g173643 (n_9259, n_9256);
  nand g173642__5526 (n_9258, g4558, n_9257);
  nand g173644__6783 (n_9256, g4558, g4555);
  fflopd g4515_reg(.CK (clock), .D (n_9255), .Q (g4515));
  fflopd g4558_reg(.CK (clock), .D (n_9254), .Q (g4558));
  fflopd g4527_reg(.CK (clock), .D (n_9253), .Q (g4527));
  nand g173649__3680 (n_9255, n_9252, n_9251);
  nand g173650__1617 (n_9254, n_1881, n_9250);
  nand g173655__2802 (n_9253, n_9239, n_9249);
  fflopd g4483_reg(.CK (clock), .D (g_5902), .Q (g4483));
  nand g173653__1705 (n_9252, g4527, n_9248);
  nand g173654__5122 (n_9251, g35, n_9247);
  fflopd g4520_reg(.CK (clock), .D (g4519), .Q (g_5902));
  nand g173652__8246 (n_9250, g4555, n_9257);
  nand g173658__7098 (n_9249, g35, n_9246);
  nand g173659__6131 (n_9248, g35, n_9245);
  nand g173660__1881 (n_9247, n_9240, n_9244);
  fflopd g4519_reg(.CK (clock), .D (n_9241), .Q (g4519));
  not g173664 (n_9246, n_9242);
  fflopd g4555_reg(.CK (clock), .D (g_5903), .Q (g4555));
  nand g173662__5115 (n_9245, n_9243, n_3364);
  nand g173663__7482 (n_9244, n_9243, n_2977);
  nand g173667__4733 (n_9242, n_9243, n_5267);
  fflopd g4571_reg(.CK (clock), .D (g4570), .Q (g_5903));
  nand g173665__6161 (n_9241, n_1271, n_9238);
  nand g173666__9315 (n_9240, g4515, g4521);
  nand g173668__9945 (n_9239, g4521, n_3854);
  not g173669 (n_9243, g4521);
  fflopd g4521_reg(.CK (clock), .D (n_9237), .Q (g4521));
  fflopd g4570_reg(.CK (clock), .D (n_9235), .Q (g4570));
  nand g173672__2883 (n_9238, g35, n_9236);
  fflopd g2799_reg(.CK (clock), .D (n_9234), .Q (g2799));
  nand g173675__2346 (n_9237, n_9232, n_7915);
  nand g173676__1666 (n_9236, n_8154, n_9233);
  nand g173677__7410 (n_9235, n_9231, n_8303);
  nand g173678__6417 (n_9234, n_8435, n_9230);
  nand g173679__5477 (n_9233, g4512, n_3677);
  nand g173680__2398 (n_9232, g4512, n_9257);
  nand g173682__5107 (n_9231, g4552, n_9193);
  fflopd g2661_reg(.CK (clock), .D (n_9227), .Q (g2661));
  fflopd g1834_reg(.CK (clock), .D (n_10438), .Q (g1834));
  fflopd g1700_reg(.CK (clock), .D (n_10435), .Q (g1700));
  fflopd g2527_reg(.CK (clock), .D (n_10444), .Q (g2527));
  not g173685 (n_9230, n_9229);
  fflopd g2102_reg(.CK (clock), .D (n_9223), .Q (g2102));
  fflopd g2393_reg(.CK (clock), .D (n_9228), .Q (g2393));
  fflopd g1968_reg(.CK (clock), .D (n_10441), .Q (g1968));
  fflopd g2259_reg(.CK (clock), .D (n_10447), .Q (g2259));
  fflopd g1724_reg(.CK (clock), .D (n_9216), .Q (g1724));
  fflopd g1858_reg(.CK (clock), .D (n_9215), .Q (g1858));
  fflopd g2685_reg(.CK (clock), .D (n_9220), .Q (g2685));
  fflopd g2417_reg(.CK (clock), .D (n_9218), .Q (g2417));
  fflopd g2551_reg(.CK (clock), .D (n_9219), .Q (g2551));
  fflopd g4552_reg(.CK (clock), .D (n_9210), .Q (g4552));
  nand g173686__6260 (n_9229, n_9217, n_8524);
  fflopd g1992_reg(.CK (clock), .D (n_9214), .Q (g1992));
  fflopd g2126_reg(.CK (clock), .D (n_9212), .Q (g2126));
  fflopd g4512_reg(.CK (clock), .D (n_9213), .Q (g4512));
  fflopd g2283_reg(.CK (clock), .D (n_9211), .Q (g2283));
  nand g173762__4319 (n_9228, n_9099, n_9197);
  nand g173756__8428 (n_9227, n_9106, n_9209);
  nand g173760__1617 (n_9223, n_9102, n_9199);
  fflopd g4300_reg(.CK (clock), .D (n_9196), .Q (g4300));
  fflopd g2036_reg(.CK (clock), .D (n_9207), .Q (g2036));
  fflopd g2327_reg(.CK (clock), .D (n_9205), .Q (g2327));
  fflopd g2193_reg(.CK (clock), .D (n_9206), .Q (g2193));
  fflopd g2595_reg(.CK (clock), .D (n_9203), .Q (g2595));
  fflopd g1768_reg(.CK (clock), .D (n_9208), .Q (g1768));
  nand g173761__5122 (n_9220, n_540, n_9189);
  nand g173724__8246 (n_9219, n_709, n_9190);
  nand g173725__7098 (n_9218, n_1045, n_9191);
  nand g173689__6131 (n_9217, g20654, n_9257);
  nand g173750__1881 (n_9216, n_1131, n_9195);
  fflopd g1902_reg(.CK (clock), .D (n_9183), .Q (g1902));
  nand g173751__5115 (n_9215, n_1404, n_9187);
  nand g173752__7482 (n_9214, n_1061, n_9186);
  nand g173690__4733 (n_9213, n_9194, n_8164);
  nand g173753__6161 (n_9212, n_557, n_9185);
  nand g173754__9315 (n_9211, n_691, n_9192);
  nand g173691__9945 (n_9210, n_9188, n_8304);
  not g173821 (n_9209, n_9181);
  nand g173768__2883 (n_9208, n_1222, n_9163);
  nand g173770__2346 (n_9207, n_738, n_9158);
  nand g173771__1666 (n_9206, n_1063, n_9155);
  nand g173772__7410 (n_9205, n_637, n_9151);
  nand g173764__6417 (n_9203, n_757, n_9159);
  not g173830 (n_9199, n_9177);
  not g173834 (n_9197, n_9176);
  nand g173681__5477 (n_9196, n_1371, n_9154);
  fflopd g2657_reg(.CK (clock), .D (n_9173), .Q (g2657));
  fflopd g1830_reg(.CK (clock), .D (n_9174), .Q (g1830));
  fflopd g2461_reg(.CK (clock), .D (n_9175), .Q (g2461));
  fflopd g2413_reg(.CK (clock), .D (n_9172), .Q (g2413));
  fflopd g2681_reg(.CK (clock), .D (n_9167), .Q (g2681));
  fflopd g1854_reg(.CK (clock), .D (n_9162), .Q (g1854));
  fflopd g2279_reg(.CK (clock), .D (n_9153), .Q (g2279));
  fflopd g1720_reg(.CK (clock), .D (n_9165), .Q (g1720));
  fflopd g1988_reg(.CK (clock), .D (n_9160), .Q (g1988));
  fflopd g2122_reg(.CK (clock), .D (n_9157), .Q (g2122));
  fflopd g2547_reg(.CK (clock), .D (n_9170), .Q (g2547));
  not g173825 (n_9195, n_9164);
  nand g173710__2398 (n_9194, g4504, n_9193);
  not g173833 (n_9192, n_9152);
  not g173818 (n_9191, n_9169);
  not g173820 (n_9190, n_9171);
  not g173822 (n_9189, n_9166);
  nand g173708__5107 (n_9188, g4549, n_9193);
  not g173827 (n_9187, n_9161);
  not g173829 (n_9186, n_9168);
  not g173831 (n_9185, n_9156);
  fflopd g117_reg(.CK (clock), .D (n_9150), .Q (g21270));
  fflopd g121_reg(.CK (clock), .D (n_9149), .Q (g20654));
  nand g173840__4319 (n_9183, n_9098, n_9147);
  nand g173850__5526 (n_9181, n_1316, n_9145);
  nand g173868__2802 (n_9177, n_681, n_9141);
  nand g173877__1705 (n_9176, n_1147, n_9139);
  fflopd g807_reg(.CK (clock), .D (n_9148), .Q (g807));
  fflopd g2652_reg(.CK (clock), .D (n_9136), .Q (g2652));
  fflopd g1825_reg(.CK (clock), .D (n_9137), .Q (g1825));
  fflopd g2093_reg(.CK (clock), .D (n_9138), .Q (g2093));
  nand g173763__5122 (n_9175, n_1189, n_9084);
  nand g173777__8246 (n_9174, n_1334, n_9109);
  nand g173779__7098 (n_9173, n_1151, n_9110);
  nand g173835__6131 (n_9172, n_9089, n_9047);
  nand g173846__1881 (n_9171, n_9019, n_9116);
  nand g173845__5115 (n_9170, n_9115, n_9059);
  nand g173841__7482 (n_9169, n_9017, n_9085);
  fflopd g554_reg(.CK (clock), .D (n_9113), .Q (g554));
  fflopd g1964_reg(.CK (clock), .D (n_9112), .Q (g1964));
  fflopd g2523_reg(.CK (clock), .D (n_9111), .Q (g2523));
  fflopd g2098_reg(.CK (clock), .D (n_9097), .Q (g2098));
  fflopd g1811_reg(.CK (clock), .D (n_9124), .Q (g1811));
  fflopd g2079_reg(.CK (clock), .D (n_9131), .Q (g2079));
  fflopd g2638_reg(.CK (clock), .D (n_9117), .Q (g2638));
  fflopd g1792_reg(.CK (clock), .D (n_9086), .Q (g1792));
  fflopd g2060_reg(.CK (clock), .D (n_9108), .Q (g2060));
  fflopd g2619_reg(.CK (clock), .D (n_9087), .Q (g2619));
  nand g173865__4733 (n_9168, n_9014, n_9130);
  nand g173851__6161 (n_9167, n_9135, n_9056);
  nand g173852__9315 (n_9166, n_9016, n_9120);
  nand g173855__9945 (n_9165, n_9122, n_9055);
  nand g173856__2883 (n_9164, n_9018, n_9123);
  nand g173857__2346 (n_9163, g35, n_9095);
  nand g173860__1666 (n_9162, n_9126, n_9052);
  nand g173861__7410 (n_9161, n_9015, n_9127);
  nand g173864__6417 (n_9160, n_9129, n_9051);
  nand g173848__5477 (n_9159, g35, n_9096);
  nand g173866__2398 (n_9158, g35, n_9093);
  nand g173869__5107 (n_9157, n_9133, n_9049);
  nand g173870__6260 (n_9156, n_9013, n_9134);
  nand g173871__4319 (n_9155, g35, n_9092);
  nand g173687__8428 (n_9154, g35, n_10112);
  nand g173873__5526 (n_9153, n_9090, n_9048);
  nand g173874__6783 (n_9152, n_9012, n_9118);
  nand g173876__3680 (n_9151, g35, n_9104);
  nand g173766__1617 (n_9150, n_9046, n_8792);
  nand g173767__2802 (n_9149, n_9057, n_8794);
  nand g174367__1705 (n_9148, n_9031, n_9073);
  not g173953 (n_9147, n_9094);
  nand g173977__8246 (n_9145, g35, n_9042);
  nand g173987__5115 (n_9141, g35, n_9038);
  nand g173991__4733 (n_9139, g35, n_9036);
  fflopd g4549_reg(.CK (clock), .D (n_9034), .Q (g4549));
  fflopd g4504_reg(.CK (clock), .D (n_9077), .Q (g4504));
  fflopd g1632_reg(.CK (clock), .D (n_9062), .Q (g1632));
  fflopd g2389_reg(.CK (clock), .D (n_10418), .Q (g2389));
  fflopd g1959_reg(.CK (clock), .D (n_9035), .Q (g1959));
  fflopd g2518_reg(.CK (clock), .D (n_9044), .Q (g2518));
  fflopd g1691_reg(.CK (clock), .D (n_9075), .Q (g1691));
  fflopd g2384_reg(.CK (clock), .D (n_9076), .Q (g2384));
  nand g173867__6161 (n_9138, n_8975, n_9050);
  nand g173858__9315 (n_9137, n_8788, n_9053);
  nand g173849__9945 (n_9136, n_8803, n_9058);
  fflopd g2255_reg(.CK (clock), .D (n_10416), .Q (g2255));
  fflopd g1696_reg(.CK (clock), .D (n_10414), .Q (g1696));
  fflopd g2504_reg(.CK (clock), .D (n_9078), .Q (g2504));
  fflopd g1677_reg(.CK (clock), .D (n_9079), .Q (g1677));
  fflopd g1945_reg(.CK (clock), .D (n_9080), .Q (g1945));
  fflopd g2370_reg(.CK (clock), .D (n_9033), .Q (g2370));
  fflopd g2236_reg(.CK (clock), .D (n_9081), .Q (g2236));
  fflopd g2250_reg(.CK (clock), .D (n_9070), .Q (g2250));
  fflopd g1894_reg(.CK (clock), .D (n_9068), .Q (g1894));
  fflopd g2485_reg(.CK (clock), .D (n_9071), .Q (g2485));
  fflopd g1624_reg(.CK (clock), .D (n_9069), .Q (g1624));
  fflopd g2453_reg(.CK (clock), .D (n_9082), .Q (g2453));
  fflopd g2587_reg(.CK (clock), .D (n_9065), .Q (g2587));
  fflopd g1926_reg(.CK (clock), .D (n_9072), .Q (g1926));
  fflopd g1760_reg(.CK (clock), .D (n_9064), .Q (g1760));
  fflopd g2185_reg(.CK (clock), .D (n_9067), .Q (g2185));
  fflopd g2028_reg(.CK (clock), .D (n_9063), .Q (g2028));
  fflopd g2319_reg(.CK (clock), .D (n_9066), .Q (g2319));
  nand g173912__2883 (n_9135, g2681, n_9119);
  nand g173895__2346 (n_9134, g2126, n_9132);
  nand g173896__1666 (n_9133, g2122, n_9132);
  nand g173897__7410 (n_9131, n_1124, n_9023);
  nand g173898__6417 (n_9130, g1992, n_9128);
  nand g173899__5477 (n_9129, g1988, n_9128);
  nand g173901__2398 (n_9127, g1858, n_9125);
  nand g173902__5107 (n_9126, g1854, n_9125);
  nand g173903__6260 (n_9124, n_1223, n_9021);
  nand g173905__4319 (n_9123, g1724, n_9121);
  nand g173906__8428 (n_9122, g1720, n_9121);
  nand g173911__5526 (n_9120, g2685, n_9119);
  nand g173892__6783 (n_9118, g2283, n_9100);
  nand g173914__3680 (n_9117, n_767, n_9022);
  nand g173915__1617 (n_9116, g2551, n_9114);
  nand g173916__2802 (n_9115, g2547, n_9114);
  nand g174391__1705 (n_9113, n_5278, n_9026);
  nand g173776__5122 (n_9112, n_635, n_9029);
  nand g173780__8246 (n_9111, n_1314, n_9030);
  not g173951 (n_9110, n_9045);
  not g173952 (n_9109, n_9054);
  nand g173956__7098 (n_9108, n_8741, n_9008);
  nand g173957__6131 (n_9107, g2527, n_9114);
  nand g173958__1881 (n_9106, g2661, n_9119);
  nand g173959__5115 (n_9105, g1700, n_9121);
  nand g174018__7482 (n_9104, n_8988, n_8942);
  nand g173961__4733 (n_9103, g1968, n_9128);
  nand g173962__6161 (n_9102, g2102, n_9132);
  nand g173963__9315 (n_9101, g2259, n_9100);
  nand g173964__9945 (n_9099, g2393, n_9088);
  nand g173984__2883 (n_9098, g35, n_9032);
  nand g173986__2346 (n_9097, n_9007, n_8927);
  nand g173997__1666 (n_9096, n_8992, n_8948);
  nand g174005__7410 (n_9095, n_8991, n_8946);
  nand g174009__6417 (n_9094, n_730, n_9020);
  nand g174013__5477 (n_9093, n_8990, n_8944);
  nand g174016__2398 (n_9092, n_8989, n_8943);
  nand g173960__5107 (n_9091, g1834, n_9125);
  nand g173891__6260 (n_9090, g2279, n_9100);
  nand g173888__4319 (n_9089, g2413, n_9088);
  nand g173886__8428 (n_9087, n_8746, n_9010);
  nand g173885__5526 (n_9086, n_8727, n_9009);
  nand g173883__6783 (n_9085, g2417, n_9088);
  nand g173842__3680 (n_9084, g35, n_9024);
  fflopd g794_reg(.CK (clock), .D (n_9027), .Q (g794));
  fflopd g74_reg(.CK (clock), .D (n_8999), .Q (g20763));
  fflopd g1657_reg(.CK (clock), .D (n_9006), .Q (g1657));
  fflopd g2217_reg(.CK (clock), .D (n_9011), .Q (g2217));
  fflopd g2351_reg(.CK (clock), .D (n_9025), .Q (g2351));
  nand g173968__2802 (n_9082, n_8907, n_8966);
  nand g173894__1705 (n_9081, n_508, n_8963);
  nand g173900__5122 (n_9080, n_735, n_8964);
  nand g173907__8246 (n_9079, n_489, n_8961);
  nand g173917__7098 (n_9078, n_932, n_8965);
  nand g173774__6131 (n_9077, n_8937, n_9193);
  nand g173775__1881 (n_9076, n_8932, n_8968);
  nand g173778__5115 (n_9075, n_8925, n_8972);
  nand g174476__4733 (n_9073, n_8904, n_8969);
  nand g173965__6161 (n_9072, n_8702, n_8928);
  nand g173966__9315 (n_9071, n_8699, n_8967);
  nand g173893__9945 (n_9070, n_1383, n_8960);
  nand g173969__2883 (n_9069, n_8908, n_8923);
  nand g173970__2346 (n_9068, n_8909, n_8939);
  nand g173971__1666 (n_9067, n_8910, n_8930);
  nand g173972__7410 (n_9066, n_8911, n_8931);
  nand g173973__6417 (n_9065, n_8869, n_8924);
  nand g173974__5477 (n_9064, n_8883, n_8926);
  nand g173975__2398 (n_9063, n_8857, n_8929);
  nand g173980__5107 (n_9062, n_8922, n_8941);
  nand g173995__8428 (n_9059, g2541, n_8976);
  nand g173998__5526 (n_9058, g2638, n_8953);
  nand g173838__6783 (n_9057, g2831, n_9257);
  nand g174000__3680 (n_9056, g2675, n_8982);
  nand g174004__1617 (n_9055, g1714, n_8977);
  nand g174006__2802 (n_9054, n_8833, n_8957);
  nand g174007__1705 (n_9053, g1811, n_8951);
  nand g174008__5122 (n_9052, g1848, n_8979);
  nand g174012__8246 (n_9051, g1982, n_8978);
  nand g174014__7098 (n_9050, g2079, n_8947);
  nand g174015__6131 (n_9049, g2116, n_8980);
  nand g174017__1881 (n_9048, g2273, n_8983);
  nand g174020__5115 (n_9047, g2407, n_8981);
  nand g173837__7482 (n_9046, g2834, n_9257);
  nand g173999__4733 (n_9045, n_8834, n_8958);
  nand g173843__6161 (n_9044, n_8787, n_8974);
  not g174136 (n_9042, n_8985);
  not g174140 (n_9038, n_9001);
  not g174142 (n_9036, n_9005);
  nand g173862__9315 (n_9035, n_8786, n_8971);
  nand g173878__9945 (n_9034, n_8938, n_9193);
  nand g173890__2883 (n_9033, n_863, n_8962);
  not g174034 (n_9032, n_8945);
  nor g174458__2346 (n_9031, n_1665, n_8906);
  not g173950 (n_9030, n_8973);
  not g173954 (n_9029, n_8970);
  nand g174474__1666 (n_9027, n_8905, n_8830);
  nand g174532__7410 (n_9026, g807, n_8901);
  nand g173988__6417 (n_9025, n_8739, n_8878);
  nand g173992__5477 (n_9024, n_8892, n_8845);
  not g174024 (n_9023, n_8956);
  not g174026 (n_9022, n_8955);
  not g174027 (n_9021, n_8954);
  nand g174090__2398 (n_9020, n_7413, n_8921);
  nand g174073__5107 (n_9019, n_2236, n_8986);
  nand g174074__6260 (n_9018, n_2204, n_8993);
  nand g174077__4319 (n_9017, n_2223, n_9004);
  nand g174079__8428 (n_9016, n_2225, n_8984);
  nand g174081__5526 (n_9015, n_2257, n_8995);
  nand g174083__6783 (n_9014, n_2293, n_8997);
  nand g174085__3680 (n_9013, n_2122, n_9000);
  nand g174087__1617 (n_9012, n_2321, n_9002);
  not g173881 (g23652, g2834);
  not g173882 (g23759, g2831);
  fflopd g2803_reg(.CK (clock), .D (n_8873), .Q (g2803));
  fflopd g2771_reg(.CK (clock), .D (n_8874), .Q (g2771));
  fflopd g1783_reg(.CK (clock), .D (n_8868), .Q (g1783));
  fflopd g1917_reg(.CK (clock), .D (n_8866), .Q (g1917));
  fflopd g2208_reg(.CK (clock), .D (n_8861), .Q (g2208));
  fflopd g2342_reg(.CK (clock), .D (n_8859), .Q (g2342));
  fflopd g2051_reg(.CK (clock), .D (n_8863), .Q (g2051));
  nand g173884__2802 (n_9011, n_8740, n_8880);
  not g174111 (n_9010, n_8933);
  not g174121 (n_9009, n_8934);
  not g174125 (n_9008, n_8935);
  not g174126 (n_9007, n_8936);
  nand g173887__1705 (n_9006, n_8757, n_8882);
  nand g174217__5122 (n_9005, n_7260, n_9004);
  nand g174215__7098 (n_9001, n_7571, n_9000);
  nand g173749__6131 (n_8999, n_4890, n_8884);
  nand g174154__4733 (n_8992, n_1552, n_8856);
  nand g174180__6161 (n_8991, n_1803, n_8915);
  nand g174191__9315 (n_8990, n_1557, n_8917);
  nand g174196__9945 (n_8989, n_1763, n_8919);
  nand g174203__2883 (n_8988, n_1427, n_8913);
  nand g174210__1666 (n_8985, n_7263, n_8984);
  not g174146 (n_9100, n_8983);
  not g174149 (n_9119, n_8982);
  not g174148 (n_9088, n_8981);
  not g174147 (n_9132, n_8980);
  not g174150 (n_9125, n_8979);
  not g174145 (n_9128, n_8978);
  not g174144 (n_9121, n_8977);
  not g174143 (n_9114, n_8976);
  fflopd g1648_reg(.CK (clock), .D (n_8871), .Q (g1648));
  fflopd g2610_reg(.CK (clock), .D (n_8875), .Q (g2610));
  fflopd g2476_reg(.CK (clock), .D (n_8900), .Q (g2476));
  nand g174100__7410 (n_8975, g35, n_8840);
  nand g173993__6417 (n_8974, g2504, n_8813);
  nand g173994__5477 (n_8973, n_8681, n_8817);
  nand g174003__2398 (n_8972, g1677, n_8790);
  nand g174010__5107 (n_8971, g1945, n_8832);
  nand g174011__6260 (n_8970, n_8664, n_8816);
  not g174603 (n_8969, n_8903);
  nand g174019__4319 (n_8968, g2370, n_8804);
  not g174022 (n_8967, n_8899);
  not g174023 (n_8966, n_8898);
  not g174025 (n_8965, n_8897);
  not g174028 (n_8964, n_8896);
  not g174029 (n_8963, n_8895);
  not g174031 (n_8962, n_8893);
  not g174033 (n_8961, n_8891);
  not g174030 (n_8960, n_8894);
  nand g174041__5526 (n_8958, g2657, n_8952);
  nand g174051__6783 (n_8957, g1830, n_8950);
  nand g174057__3680 (n_8956, n_8780, n_8809);
  nand g174059__1617 (n_8955, n_8777, n_8810);
  nand g174060__2802 (n_8954, n_8775, n_8848);
  nand g174070__1705 (n_8953, n_8571, n_8952);
  nand g174071__5122 (n_8951, n_8574, n_8950);
  nand g174078__7098 (n_8948, g2595, n_8855);
  nand g174101__6131 (n_8947, g35, n_8839);
  nand g174080__1881 (n_8946, g1768, n_8914);
  nand g174082__5115 (n_8945, g1902, n_8920);
  nand g174084__7482 (n_8944, g2036, n_8916);
  nand g174086__4733 (n_8943, g2193, n_8918);
  nand g174088__6161 (n_8942, g2327, n_8912);
  nand g174098__9315 (n_8941, g35, n_8841);
  fflopd g4242_reg(.CK (clock), .D (n_8835), .Q (g4242));
  fflopd g2831_reg(.CK (clock), .D (n_8795), .Q (g2831));
  fflopd g2834_reg(.CK (clock), .D (n_8793), .Q (g2834));
  fflopd g2775_reg(.CK (clock), .D (n_8802), .Q (g2775));
  not g174122 (n_8939, n_8867);
  not g173880 (n_8938, g4546);
  not g173879 (n_8937, g4501);
  nand g174194__2883 (n_8936, n_1205, n_8850);
  nand g174193__2346 (n_8935, n_1369, n_8849);
  nand g174182__1666 (n_8934, n_1266, n_8837);
  nand g174156__7410 (n_8933, n_705, n_8807);
  not g174132 (n_8932, n_8858);
  not g174130 (n_8931, n_8860);
  not g174127 (n_8930, n_8862);
  not g174124 (n_8929, n_8864);
  not g174123 (n_8928, n_8865);
  nand g174102__6417 (n_8927, g35, n_8838);
  not g174120 (n_8926, n_8885);
  not g174117 (n_8925, n_8870);
  not g174110 (n_8924, n_8876);
  not g174115 (n_8923, n_8872);
  nand g174218__5477 (n_8976, g35, n_8854);
  fflopd g355_reg(.CK (clock), .D (n_8811), .Q (g355));
  nand g174225__2398 (n_8979, g35, n_8888);
  nand g174224__5107 (n_8982, g35, n_8853);
  nand g174223__6260 (n_8981, g35, n_8890);
  nand g174222__4319 (n_8980, g35, n_8886);
  nand g174221__8428 (n_8983, g35, n_8887);
  nand g174220__5526 (n_8978, g35, n_8889);
  nand g174219__6783 (n_8977, g35, n_8852);
  fflopd g2827_reg(.CK (clock), .D (n_8818), .Q (g2827));
  fflopd g2767_reg(.CK (clock), .D (n_8846), .Q (g2767));
  fflopd g2823_reg(.CK (clock), .D (n_8819), .Q (g2823));
  fflopd g2811_reg(.CK (clock), .D (n_8820), .Q (g2811));
  fflopd g2791_reg(.CK (clock), .D (n_8851), .Q (g2791));
  fflopd g2779_reg(.CK (clock), .D (n_8847), .Q (g2779));
  fflopd g2795_reg(.CK (clock), .D (n_8821), .Q (g2795));
  fflopd g790_reg(.CK (clock), .D (n_8831), .Q (g790));
  fflopd g2807_reg(.CK (clock), .D (n_8799), .Q (g2807));
  fflopd g2787_reg(.CK (clock), .D (n_8800), .Q (g2787));
  fflopd g2783_reg(.CK (clock), .D (n_8801), .Q (g2783));
  fflopd g2819_reg(.CK (clock), .D (n_8797), .Q (g2819));
  fflopd g2815_reg(.CK (clock), .D (n_8798), .Q (g2815));
  not g174032 (n_8922, n_8814);
  fflopd g4546_reg(.CK (clock), .D (n_8725), .Q (g4546));
  not g174338 (n_8921, n_8920);
  not g174339 (n_8919, n_8918);
  not g174340 (n_8917, n_8916);
  not g174341 (n_8915, n_8914);
  not g174342 (n_8913, n_8912);
  nand g174092__3680 (n_8911, n_8822, n_8721);
  nand g174091__1617 (n_8910, n_8824, n_8720);
  nand g174089__2802 (n_8909, n_8823, n_8719);
  nand g174076__1705 (n_8908, n_2109, n_8722);
  nand g174075__5122 (n_8907, n_2534, n_8718);
  nor g174582__8246 (n_8906, g807, n_8902);
  nand g174616__7098 (n_8905, n_8904, n_8743);
  nand g174619__6131 (n_8903, g807, n_8902);
  nand g174620__1881 (n_8901, g35, n_8902);
  fflopd g4501_reg(.CK (clock), .D (n_8726), .Q (g4501));
  nand g174036__5115 (n_8900, n_8745, n_8684);
  nand g174037__7482 (n_8899, n_679, n_8761);
  nand g174039__4733 (n_8898, n_722, n_8763);
  nand g174058__6161 (n_8897, n_8778, n_8660);
  nand g174061__9315 (n_8896, n_8774, n_8693);
  nand g174063__9945 (n_8895, n_8773, n_8712);
  nand g174064__2883 (n_8894, n_8772, n_8710);
  nand g174065__2346 (n_8893, n_8770, n_8709);
  nand g174066__1666 (n_8892, n_1867, n_8724);
  nand g174068__7410 (n_8891, n_8728, n_8704);
  not g174345 (n_9004, n_8890);
  not g174346 (n_8997, n_8889);
  not g174347 (n_8995, n_8888);
  not g174344 (n_9002, n_8887);
  not g174343 (n_9000, n_8886);
  nand g174179__6417 (n_8885, n_760, n_8765);
  not g173823 (n_8884, n_8796);
  nand g174094__5477 (n_8883, n_8826, n_8781);
  not g174116 (n_8882, n_8791);
  not g174128 (n_8880, n_8785);
  not g174131 (n_8878, n_8783);
  nand g174153__2398 (n_8876, n_560, n_8767);
  nand g174155__5107 (n_8875, n_8744, n_8680);
  nand g174159__6260 (n_8874, n_782, n_8734);
  nand g174163__4319 (n_8873, n_647, n_8733);
  nand g174172__8428 (n_8872, n_1391, n_8760);
  nand g174173__5526 (n_8871, n_8758, n_8670);
  nand g174176__6783 (n_8870, n_3174, n_8776);
  nand g174093__3680 (n_8869, n_8829, n_8782);
  nand g174181__1617 (n_8868, n_8735, n_8646);
  nand g174185__2802 (n_8867, n_891, n_8756);
  nand g174186__1705 (n_8866, n_8754, n_8667);
  nand g174187__5122 (n_8865, n_961, n_8742);
  nand g174190__8246 (n_8864, n_843, n_8753);
  nand g174192__7098 (n_8863, n_8751, n_8663);
  nand g174195__6131 (n_8862, n_1283, n_8750);
  nand g174197__1881 (n_8861, n_8749, n_8662);
  nand g174201__5115 (n_8860, n_867, n_8748);
  nand g174202__7482 (n_8859, n_8747, n_8686);
  nand g174206__4733 (n_8858, n_3087, n_8769);
  nand g174214__6161 (n_8857, n_8825, n_8779);
  not g174233 (n_8856, n_8855);
  not g174237 (n_8986, n_8854);
  not g174238 (n_8984, n_8853);
  not g174235 (n_8993, n_8852);
  nand g174044__9315 (n_8851, n_8432, n_8717);
  nand g174284__9945 (n_8850, n_2747, n_8640);
  nand g174296__2883 (n_8849, g2051, n_8808);
  nand g174254__2346 (n_8848, n_10200, n_8836);
  nand g174043__1666 (n_8847, n_8431, n_8694);
  nand g174042__7410 (n_8846, n_8430, n_8695);
  nand g174038__6417 (n_8845, g2461, n_8723);
  not g174330 (n_8841, n_8732);
  not g174333 (n_8840, n_8731);
  not g174334 (n_8839, n_8730);
  not g174335 (n_8838, n_8729);
  nand g174350__5477 (n_8837, g1783, n_8836);
  nand g173769__2398 (n_8835, n_8366, n_8638);
  nand g174379__5107 (n_8834, n_2804, n_8827);
  nand g174398__6260 (n_8833, n_2786, n_8828);
  nand g174035__4319 (n_8832, n_8575, n_8815);
  nand g174615__8428 (n_8831, n_8582, n_8637);
  nor g174581__5526 (n_8830, n_1472, n_8635);
  nand g174307__6783 (n_8855, n_8829, n_8642);
  nor g174418__3680 (n_8950, n_9257, n_8828);
  nor g174420__1617 (n_8952, n_9257, n_8827);
  nand g174423__2802 (n_8886, g2060, n_8655);
  nand g174424__1705 (n_8887, g2217, n_8650);
  nand g174425__5122 (n_8890, g2351, n_8648);
  nand g174426__8246 (n_8889, g1926, n_8653);
  nand g174427__7098 (n_8888, g1792, n_8669);
  nand g174416__6131 (n_8914, n_8826, n_8644);
  nand g174415__1881 (n_8916, n_8825, n_8654);
  nand g174414__5115 (n_8918, n_8824, n_8651);
  nand g174413__7482 (n_8920, n_8823, n_8647);
  nand g174314__4733 (n_8853, g2619, n_8641);
  nand g174312__6161 (n_8854, g2485, n_8643);
  nand g174310__9315 (n_8852, g1657, n_8652);
  nand g174417__9945 (n_8912, n_8822, n_8649);
  nand g174045__2883 (n_8821, n_8433, n_8688);
  nand g174047__2346 (n_8820, n_8436, n_8691);
  nand g174048__1666 (n_8819, n_8426, n_8690);
  nand g174049__7410 (n_8818, n_8425, n_8689);
  nand g174056__6417 (n_8817, g2523, n_8812);
  nand g174062__5477 (n_8816, g1964, n_8815);
  nand g174067__2398 (n_8814, n_1380, n_8705);
  nand g174069__5107 (n_8813, n_8570, n_8812);
  nand g173836__6260 (n_8811, n_4301, n_8632);
  nand g174253__4319 (n_8810, n_10198, n_8806);
  nand g174249__8428 (n_8809, n_10202, n_8808);
  nand g174246__5526 (n_8807, g2610, n_8806);
  nand g174207__6783 (n_8805, n_1176, n_8687);
  nand g174205__3680 (n_8804, g35, n_8714);
  nand g174157__1617 (n_8803, g2652, n_8679);
  nand g174160__2802 (n_8802, n_948, n_8677);
  nand g174161__1705 (n_8801, n_549, n_8676);
  nand g174162__5122 (n_8800, n_959, n_8675);
  nand g174164__8246 (n_8799, n_1292, n_8673);
  nand g174165__7098 (n_8798, n_789, n_8672);
  nand g174166__6131 (n_8797, n_1163, n_8671);
  nand g173853__1881 (n_8796, n_5311, n_8633);
  nand g174167__5115 (n_8795, n_1153, n_8794);
  nand g174168__7482 (n_8793, n_1248, n_8792);
  nand g174174__4733 (n_8791, n_669, n_8703);
  nand g174175__6161 (n_8790, g35, n_8707);
  nand g174177__9315 (n_8789, n_1226, n_8698);
  nand g174183__9945 (n_8788, g1825, n_8668);
  nand g174184__2883 (n_8787, g2518, n_8683);
  nand g174189__2346 (n_8786, g1959, n_8666);
  nand g174198__1666 (n_8785, n_1281, n_8701);
  nand g174199__7410 (n_8784, n_1322, n_8661);
  nand g174204__6417 (n_8783, n_1289, n_8700);
  fflopd g5808_reg(.CK (clock), .D (n_10116), .Q (g5808));
  fflopd g5462_reg(.CK (clock), .D (n_10114), .Q (g5462));
  fflopd g194_reg(.CK (clock), .D (n_8685), .Q (g8358));
  fflopd g5115_reg(.CK (clock), .D (n_8674), .Q (g5115));
  fflopd g6154_reg(.CK (clock), .D (n_8696), .Q (g6154));
  nor g174256__5477 (n_8782, n_8577, n_8630);
  nor g174257__2398 (n_8781, n_8579, n_8629);
  nand g174265__5107 (n_8780, g2079, n_8752);
  nor g174267__6260 (n_8779, n_8568, n_8631);
  nand g174272__4319 (n_8778, g2504, n_8762);
  nand g174273__8428 (n_8777, g2638, n_8766);
  nand g174275__5526 (n_8776, g1691, n_8759);
  nand g174276__6783 (n_8775, g1811, n_8764);
  nand g174277__3680 (n_8774, g1945, n_8755);
  nand g174278__1617 (n_8773, g2236, n_8771);
  nand g174279__2802 (n_8772, g2250, n_8771);
  nand g174280__1705 (n_8770, g2370, n_8768);
  nand g174281__5122 (n_8769, g2384, n_8768);
  nand g174282__8246 (n_8767, g2587, n_8766);
  nand g174283__7098 (n_8765, g1760, n_8764);
  nand g174285__6131 (n_8763, g2453, n_8762);
  nand g174286__1881 (n_8761, g2485, n_8762);
  nand g174287__5115 (n_8760, g1624, n_8759);
  nand g174288__7482 (n_8758, g1648, n_8759);
  nand g174289__4733 (n_8757, g1657, n_8759);
  nand g174291__6161 (n_8756, g1894, n_8755);
  nand g174292__9315 (n_8754, g1917, n_8755);
  nand g174294__9945 (n_8753, g2028, n_8752);
  nand g174295__2883 (n_8751, g2051, n_8752);
  nand g174297__2346 (n_8750, g2185, n_8771);
  nand g174298__1666 (n_8749, g2208, n_8771);
  nand g174300__7410 (n_8748, g2319, n_8768);
  nand g174301__6417 (n_8747, g2342, n_8768);
  nand g174303__5477 (n_8746, g2619, n_8766);
  nand g174304__2398 (n_8745, g2476, n_8762);
  nand g174306__5107 (n_8744, g2610, n_8766);
  not g174672 (n_8743, n_8636);
  nand g174352__6260 (n_8742, g1926, n_8755);
  nand g174354__4319 (n_8741, g2060, n_8752);
  nand g174356__8428 (n_8740, g2217, n_8771);
  nand g174358__5526 (n_8739, g2351, n_8768);
  nand g174380__2802 (n_8735, g1783, n_8764);
  nand g174381__1705 (n_8734, g35, n_8605);
  nand g174385__5122 (n_8733, g35, n_8604);
  nand g174392__8246 (n_8732, g1632, n_8573);
  nand g174405__7098 (n_8731, g2093, n_8608);
  nand g174406__6131 (n_8730, n_2114, n_8576);
  nand g174407__1881 (n_8729, g2098, n_8639);
  nand g174239__5115 (n_8728, g1677, n_8759);
  nand g174349__7482 (n_8727, g1792, n_8764);
  nand g174095__4733 (n_8726, n_8586, n_9193);
  nand g174096__6161 (n_8725, n_8585, n_9193);
  not g174234 (n_8724, n_8723);
  not g174231 (n_8722, n_8708);
  not g174230 (n_8721, n_8715);
  not g174229 (n_8720, n_8716);
  not g174228 (n_8719, n_8658);
  not g174227 (n_8718, n_8657);
  nand g174665__9315 (n_8902, g794, n_8584);
  fflopd g1141_reg(.CK (clock), .D (n_8589), .Q (g1141));
  fflopd g344_reg(.CK (clock), .D (n_8581), .Q (g7540));
  fflopd g785_reg(.CK (clock), .D (n_8583), .Q (g785));
  fflopd g3106_reg(.CK (clock), .D (n_10120), .Q (g3106));
  fflopd g6500_reg(.CK (clock), .D (n_10122), .Q (g6500));
  fflopd g3808_reg(.CK (clock), .D (n_10118), .Q (g3808));
  not g174321 (n_8717, n_8620);
  nand g174258__9945 (n_8716, n_8551, n_8711);
  nand g174259__2883 (n_8715, n_8548, n_8713);
  nand g174260__2346 (n_8714, n_2601, n_8713);
  nand g174261__1666 (n_8712, n_10206, n_8711);
  nand g174262__7410 (n_8710, n_2916, n_8711);
  nand g174263__6417 (n_8709, n_10208, n_8713);
  nand g174268__5477 (n_8708, n_8550, n_8706);
  nand g174269__2398 (n_8707, n_2593, n_8706);
  nand g174270__5107 (n_8705, n_2125, n_8706);
  nand g174271__6260 (n_8704, n_10382, n_8706);
  nand g174290__4319 (n_8703, g1648, n_8706);
  nand g174293__8428 (n_8702, g1917, n_8692);
  nand g174299__5526 (n_8701, g2208, n_8711);
  nand g174302__6783 (n_8700, g2342, n_8713);
  nand g174305__3680 (n_8699, g2476, n_8659);
  nand g174394__1617 (n_8698, n_2772, n_8612);
  nand g173765__1705 (n_8696, n_567, n_8540);
  not g174319 (n_8695, n_8622);
  not g174320 (n_8694, n_8621);
  nand g174255__5122 (n_8693, n_10204, n_8692);
  not g174323 (n_8691, n_8618);
  not g174324 (n_8690, n_8617);
  not g174325 (n_8689, n_8616);
  not g174322 (n_8688, n_8619);
  nand g174355__8246 (n_8687, n_2803, n_8610);
  nand g174357__7098 (n_8686, g2319, n_8564);
  nand g174359__6131 (n_8685, n_8556, n_4861);
  nand g174373__1881 (n_8684, g2453, n_8682);
  nand g174375__5115 (n_8683, n_2964, n_8682);
  nand g174376__7482 (n_8681, n_2884, n_8627);
  nand g174377__4733 (n_8680, g2587, n_8678);
  nand g174378__6161 (n_8679, n_2660, n_8678);
  nand g174382__9315 (n_8677, g35, n_8563);
  nand g174383__9945 (n_8676, g35, n_8555);
  nand g174384__2883 (n_8675, g35, n_8554);
  nand g173773__2346 (n_8674, n_1001, n_8541);
  nand g174386__1666 (n_8673, g35, n_8553);
  nand g174387__7410 (n_8672, g35, n_8552);
  nand g174388__6417 (n_8671, g35, n_8557);
  nand g174393__5477 (n_8670, g1624, n_8566);
  nand g174308__2398 (n_8723, g2476, n_8559);
  not g174438 (n_8669, n_8593);
  nand g174397__5107 (n_8668, n_2659, n_8645);
  nand g174400__6260 (n_8667, g1894, n_8665);
  nand g174401__4319 (n_8666, n_2962, n_8665);
  nand g174402__8428 (n_8664, n_2793, n_8628);
  nand g174403__5526 (n_8663, g2028, n_8567);
  nand g174409__6783 (n_8662, g2185, n_8565);
  nand g174411__3680 (n_8661, n_2731, n_8614);
  nand g174252__1617 (n_8660, n_10196, n_8659);
  nand g174251__2802 (n_8658, n_8549, n_8692);
  nand g174250__1705 (n_8657, n_8546, n_8659);
  not g174428 (n_8655, n_8609);
  not g174429 (n_8654, n_8606);
  not g174431 (n_8653, n_8603);
  not g174432 (n_8652, n_8602);
  not g174433 (n_8651, n_8601);
  not g174434 (n_8650, n_8600);
  not g174435 (n_8649, n_8598);
  not g174436 (n_8648, n_8597);
  not g174437 (n_8647, n_8595);
  nand g174396__8246 (n_8646, g1760, n_8645);
  not g174439 (n_8644, n_8592);
  not g174440 (n_8643, n_8590);
  not g174441 (n_8642, n_8626);
  not g174442 (n_8641, n_8588);
  not g174502 (n_8640, n_8639);
  nand g173839__7098 (n_8638, g35, n_8535);
  nand g174693__6131 (n_8637, n_8904, n_8536);
  nand g174687__1881 (n_8636, g794, n_8634);
  nor g174658__5115 (n_8635, g794, n_8634);
  nand g173979__7482 (n_8633, g35, n_8538);
  nand g173978__4733 (n_8632, n_5310, n_10124);
  not g174509 (n_8808, n_8631);
  not g174508 (n_8806, n_8630);
  not g174507 (n_8836, n_8629);
  nor g174412__6161 (n_8815, n_9257, n_8628);
  not g174506 (n_8828, n_8580);
  not g174503 (n_8827, n_8578);
  nor g174422__9315 (n_8794, n_8531, n_8561);
  nor g174421__9945 (n_8792, n_8532, n_8562);
  nor g174419__2883 (n_8812, n_9257, n_8627);
  fflopd g2902_reg(.CK (clock), .D (n_8558), .Q (g2902));
  nand g174486__2346 (n_8626, g2610, n_8587);
  nand g174360__5477 (n_8622, n_8511, n_8529);
  nand g174361__2398 (n_8621, n_504, n_8527);
  nand g174362__5107 (n_8620, n_1240, n_8526);
  nand g174363__6260 (n_8619, n_1255, n_8525);
  nand g174364__4319 (n_8618, n_825, n_8523);
  nand g174365__8428 (n_8617, n_578, n_8533);
  nand g174366__5526 (n_8616, n_1114, n_8522);
  nand g174448__6783 (n_8609, g2028, n_8607);
  nand g174449__3680 (n_8608, n_1957, n_8607);
  nand g174450__1617 (n_8606, g2051, n_8607);
  nand g174460__2802 (n_8605, n_8519, n_8481);
  nand g174461__1705 (n_8604, n_8518, n_8482);
  nand g174472__5122 (n_8603, g1894, n_8594);
  nand g174477__8246 (n_8602, g1624, n_8572);
  nand g174478__7098 (n_8601, g2208, n_8599);
  nand g174479__6131 (n_8600, g2185, n_8599);
  nand g174480__1881 (n_8598, g2342, n_8596);
  nand g174481__5115 (n_8597, g2319, n_8596);
  nand g174482__7482 (n_8595, g1917, n_8594);
  nand g174483__4733 (n_8593, g1760, n_8591);
  nand g174484__6161 (n_8592, g1783, n_8591);
  nand g174485__9315 (n_8590, g2453, n_8569);
  nand g174266__9945 (n_8589, n_8439, n_8521);
  nand g174487__2883 (n_8588, g2587, n_8587);
  not g174232 (n_8586, g4498);
  not g174226 (n_8585, g4567);
  not g174710 (n_8584, n_8634);
  nand g174691__2346 (n_8583, n_8516, n_8469);
  nor g174657__1666 (n_8582, n_1450, n_8508);
  nand g174001__7410 (n_8581, n_8504, n_2049);
  nand g174552__6417 (n_8580, n_8579, n_8591);
  nand g174549__5477 (n_8578, n_8577, n_8587);
  nand g174521__2398 (n_8576, n_1047, n_8607);
  nand g174522__5107 (n_8575, n_1079, n_8594);
  nand g174524__6260 (n_8574, n_1081, n_8591);
  nand g174525__4319 (n_8573, g25167, n_8572);
  nand g174526__8428 (n_8571, n_1083, n_8587);
  nand g174529__5526 (n_8570, n_1085, n_8569);
  fflopd g534_reg(.CK (clock), .D (n_8512), .Q (g534));
  nand g174553__6783 (n_8629, g35, n_8591);
  nand g174554__3680 (n_8630, g35, n_8587);
  nand g174557__1617 (n_8631, g35, n_8607);
  fflopd g4821_reg(.CK (clock), .D (n_8510), .Q (g4821));
  fflopd g4831_reg(.CK (clock), .D (n_8509), .Q (g4831));
  nand g174548__2802 (n_8639, n_8568, n_8607);
  not g174514 (n_8755, n_8665);
  not g174513 (n_8764, n_8645);
  fflopd g3457_reg(.CK (clock), .D (n_8520), .Q (g3457));
  not g174510 (n_8752, n_8567);
  not g174511 (n_8766, n_8678);
  not g174515 (n_8762, n_8682);
  not g174512 (n_8759, n_8566);
  not g174516 (n_8771, n_8565);
  not g174517 (n_8768, n_8564);
  nand g174540__1705 (n_8563, n_8467, n_8491);
  nor g174527__5122 (n_8562, n_4825, n_8560);
  nor g174528__8246 (n_8561, n_4852, n_8560);
  nor g174530__7098 (n_8559, g2485, n_8547);
  nand g174537__6131 (n_8558, n_693, n_8483);
  nand g174539__1881 (n_8557, n_8466, n_8492);
  nand g174523__5115 (n_8556, g222, n_9257);
  nand g174541__7482 (n_8555, n_8463, n_8498);
  nand g174542__4733 (n_8554, n_8462, n_8489);
  nand g174543__6161 (n_8553, n_8459, n_8487);
  nand g174544__9315 (n_8552, n_8457, n_8485);
  fflopd g4498_reg(.CK (clock), .D (n_8490), .Q (g4498));
  nand g174561__9945 (n_8567, g35, n_8499);
  nor g174489__2883 (n_8614, n_8551, n_8543);
  nor g174490__2346 (n_8612, n_8550, n_8542);
  nor g174491__1666 (n_8628, n_8549, n_8545);
  nor g174492__7410 (n_8610, n_8548, n_8544);
  nor g174495__6417 (n_8627, n_8546, n_8547);
  nor g174556__5477 (n_8692, n_9257, n_8545);
  nor g174555__2398 (n_8659, n_9257, n_8547);
  nor g174559__5107 (n_8713, n_9257, n_8544);
  nor g174558__6260 (n_8711, n_9257, n_8543);
  nor g174560__4319 (n_8706, n_9257, n_8542);
  fflopd g4567_reg(.CK (clock), .D (n_8497), .Q (g4567));
  nand g173875__8428 (n_8541, g35, n_8496);
  nand g173847__5526 (n_8540, g35, n_8493);
  not g174113 (n_8538, n_8514);
  not g174738 (n_8536, n_8506);
  wire w3, w4, w5, w6;
  nand g174021__6783 (n_8535, w4, w6);
  nand g9 (w6, w5, n_6474);
  not g8 (w5, n_8460);
  nand g7 (w4, w3, n_8460);
  not g6 (w3, n_6474);
  nand g174563__1617 (n_8566, g35, n_8542);
  fflopd g4035_reg(.CK (clock), .D (n_8471), .Q (g4035));
  fflopd g5011_reg(.CK (clock), .D (n_8479), .Q (g5011));
  fflopd g3333_reg(.CK (clock), .D (n_8472), .Q (g3333));
  nand g174568__2802 (n_8564, g35, n_8544);
  nand g174567__1705 (n_8565, g35, n_8543);
  nand g174564__5122 (n_8645, g35, n_8501);
  fflopd g4375_reg(.CK (clock), .D (n_8477), .Q (g4375));
  nand g174566__8246 (n_8682, g35, n_8547);
  nand g174565__7098 (n_8665, g35, n_8545);
  nand g174724__6131 (n_8634, g790, n_8473);
  nand g174562__1881 (n_8678, g35, n_8500);
  fflopd g781_reg(.CK (clock), .D (n_8470), .Q (g781));
  fflopd g1094_reg(.CK (clock), .D (n_8495), .Q (g1094));
  nand g174471__5115 (n_8533, n_68, n_8528);
  nor g174455__7482 (n_8532, n_4824, n_8530);
  nor g174456__4733 (n_8531, n_4826, n_8530);
  nand g174465__6161 (n_8529, n_122, n_8528);
  nand g174466__9315 (n_8527, n_1, n_8528);
  nand g174467__9945 (n_8526, n_53, n_8528);
  nand g174468__2883 (n_8525, n_71, n_8528);
  nand g174469__2346 (n_8524, n_126, n_8528);
  nand g174470__1666 (n_8523, n_241, n_8528);
  nand g174447__7410 (n_8522, n_233, n_8528);
  not g174498 (n_8521, n_8494);
  nand g174002__6417 (n_8520, n_1311, n_8450);
  nand g174586__5477 (n_8519, n_2, n_8517);
  nand g174587__2398 (n_8518, n_26, n_8517);
  not g174607 (n_8569, n_8547);
  not g174606 (n_8596, n_8544);
  not g174605 (n_8599, n_8543);
  not g174604 (n_8572, n_8542);
  nand g174755__5107 (n_8516, n_8904, n_8451);
  nand g174208__6260 (n_8515, n_8452, n_8446);
  nand g174169__4319 (n_8514, g333, g351);
  nand g174151__8428 (n_8513, n_8453, n_8444);
  nand g174621__5526 (n_8512, n_1204, n_8454);
  nand g174625__6783 (n_8511, g2763, n_9257);
  nand g174053__3680 (n_8510, n_5444, n_8465);
  nand g174054__1617 (n_8509, n_5446, n_8464);
  nor g174754__2802 (n_8508, g790, n_8505);
  nand g174763__1705 (n_8506, g790, n_8505);
  nand g174097__5122 (n_8504, g333, n_9257);
  fflopd g4826_reg(.CK (clock), .D (n_8455), .Q (g4826));
  not g174610 (n_8594, n_8545);
  not g174609 (n_8591, n_8501);
  not g174608 (n_8587, n_8500);
  not g174611 (n_8607, n_8499);
  nand g174592__8246 (n_8498, g2783, n_8484);
  nand g174475__7098 (n_8497, n_8441, n_9193);
  nand g173967__6131 (n_8496, n_8380, n_8414);
  nand g174534__1881 (n_8495, n_8001, n_8438);
  nand g174538__5115 (n_8494, n_657, n_8437);
  nand g173996__7482 (n_8493, n_8356, n_8417);
  fflopd g222_reg(.CK (clock), .D (n_8423), .Q (g222));
  nand g174584__4733 (n_8492, g2819, n_8488);
  nand g174591__6161 (n_8491, g2775, n_8486);
  nand g174473__9315 (n_8490, n_8449, n_9193);
  nand g174593__9945 (n_8489, g2787, n_8488);
  nand g174594__2883 (n_8487, g2807, n_8486);
  nand g174595__2346 (n_8485, g2815, n_8484);
  nand g174622__1666 (n_8483, g35, n_8424);
  nand g174623__7410 (n_8482, g2803, n_8480);
  nand g174624__6417 (n_8481, g2771, n_8480);
  nand g174630__5477 (n_8560, g35, n_8421);
  nand g174634__2398 (n_8542, n_7519, n_8468);
  nand g174055__5107 (n_8479, n_5453, n_8447);
  nand g174188__6260 (n_8477, n_4597, n_8445);
  nand g174178__4319 (n_8476, n_8408, n_8427);
  nand g174170__8428 (n_8475, n_8410, n_8422);
  nand g174158__5526 (n_8474, n_8411, n_8419);
  not g174770 (n_8473, n_8505);
  nand g174050__6783 (n_8472, n_5438, n_8440);
  nand g174052__3680 (n_8471, n_5441, n_8448);
  nand g174742__1617 (n_8470, n_8388, n_8418);
  nor g174712__2802 (n_8469, n_1491, n_8429);
  nand g174639__1705 (n_8501, n_7523, n_8468);
  nand g174638__5122 (n_8500, n_7524, n_8468);
  nand g174641__8246 (n_8499, n_7521, n_8468);
  nand g174636__7098 (n_8544, n_7520, n_8468);
  nand g174635__6131 (n_8543, n_7517, n_8468);
  nand g174640__1881 (n_8545, n_7522, n_8468);
  fflopd g128_reg(.CK (clock), .D (n_8428), .Q (g21245));
  nand g174637__5115 (n_8547, n_7525, n_8468);
  nand g174583__7482 (n_8467, n_152, n_8458);
  nand g174614__4733 (n_8466, n_61, n_8461);
  not g174332 (n_8465, n_8443);
  not g174336 (n_8464, n_8442);
  nand g174571__6161 (n_8463, n_41, n_8456);
  nand g174573__9315 (n_8462, n_193, n_8461);
  nand g174309__9945 (n_8460, n_8398, n_8395);
  nand g174612__2883 (n_8459, n_12, n_8458);
  nand g174613__2346 (n_8457, n_207, n_8456);
  nand g174632__1666 (n_8530, g35, n_8420);
  fflopd g333_reg(.CK (clock), .D (n_8403), .Q (g333));
  fflopd g1124_reg(.CK (clock), .D (n_8397), .Q (g1124));
  nand g174247__7410 (n_8455, n_5388, n_8412);
  fflopd g2763_reg(.CK (clock), .D (n_8389), .Q (g2763));
  nand g174694__6417 (n_8454, g35, n_10126);
  nand g174241__5477 (n_8453, n_8384, n_8400);
  nand g174248__2398 (n_8452, n_8382, n_8402);
  not g174804 (n_8451, n_8416);
  nand g174171__5107 (n_8450, g35, n_8405);
  not g174679 (n_8517, n_8480);
  nand g174794__6260 (n_8505, g785, n_8393);
  fflopd g1111_reg(.CK (clock), .D (n_8396), .Q (g1111));
  fflopd g776_reg(.CK (clock), .D (n_8391), .Q (g776));
  nor g174642__4319 (n_8528, n_9257, n_8392);
  not g174570 (n_8449, g4495);
  not g174331 (n_8448, n_8407);
  not g174337 (n_8447, n_8406);
  nand g174353__8428 (n_8446, g35, n_8383);
  nand g174372__5526 (n_8445, g4427, n_9257);
  nand g174374__6783 (n_8444, g35, n_8385);
  nand g174404__3680 (n_8443, n_927, n_8401);
  nand g174408__1617 (n_8442, n_1034, n_8399);
  not g174569 (n_8441, g4543);
  not g174329 (n_8440, n_8409);
  nand g174590__2802 (n_8439, n_7851, n_8368);
  not g174602 (n_8438, n_8394);
  nand g174627__1705 (n_8437, g1141, n_8369);
  nand g174648__5122 (n_8436, g2811, n_8434);
  nand g174649__8246 (n_8435, g2799, n_8434);
  nand g174650__7098 (n_8433, g2795, n_8434);
  nand g174652__6131 (n_8432, g2791, n_8434);
  nand g174654__1881 (n_8431, g2779, n_8434);
  nand g174659__5115 (n_8430, g2767, n_8434);
  nor g174775__7482 (n_8429, g785, n_8415);
  nand g174245__4733 (n_8428, n_5393, n_8378);
  nand g174244__6161 (n_8427, n_8357, n_8377);
  nand g174681__9315 (n_8426, g2823, n_8434);
  nand g174682__9945 (n_8425, g2827, n_8434);
  nand g174683__2883 (n_8424, n_8367, n_2717);
  nand g174698__2346 (n_8423, n_8363, n_8185);
  nand g174243__1666 (n_8422, n_8359, n_8375);
  not g174676 (n_8421, n_8420);
  nand g174242__7410 (n_8419, n_8351, n_8373);
  nand g174818__6417 (n_8418, n_8904, n_8365);
  nand g174152__5477 (n_8417, g6154, n_8386);
  nand g174827__2398 (n_8416, g785, n_8415);
  nand g174200__5107 (n_8414, g5115, n_8379);
  not g174680 (n_8486, n_8458);
  not g174678 (n_8488, n_8461);
  not g174677 (n_8484, n_8456);
  nand g174705__6260 (n_8480, n_8413, n_8370);
  nand g174707__4319 (n_8468, n_8413, n_8364);
  not g174430 (n_8412, n_8381);
  nand g174348__8428 (n_8411, g35, n_8352);
  nand g174389__5526 (n_8410, g35, n_8360);
  nand g174390__6783 (n_8409, n_1293, n_8374);
  nand g174395__3680 (n_8408, g35, n_8358);
  nand g174399__1617 (n_8407, n_1407, n_8376);
  nand g174410__2802 (n_8406, n_1199, n_8372);
  nand g174264__1705 (n_8405, n_8317, n_8353);
  nand g174451__5122 (n_8403, n_8121, n_8348);
  not g174500 (n_8402, n_8401);
  not g174501 (n_8400, n_8399);
  wire w7, w8, w9, w10;
  nand g174519__8246 (n_8398, w8, w10);
  nand g13 (w10, w9, g4235);
  not g12 (w9, n_8152);
  nand g11 (w8, w7, n_8152);
  not g10 (w7, g4235);
  nand g174535__7098 (n_8397, n_946, n_8349);
  nand g174536__6131 (n_8396, n_1133, n_8350);
  fflopd g4543_reg(.CK (clock), .D (n_8340), .Q (g4543));
  nand g174579__1881 (n_8395, n_8361, n_8336);
  nand g174618__5115 (n_8394, n_763, n_8342);
  not g174837 (n_8393, n_8415);
  nand g174684__7482 (n_8392, n_8319, n_8387);
  nand g174817__4733 (n_8391, n_8333, n_8322);
  fflopd g4495_reg(.CK (clock), .D (n_8341), .Q (g4495));
  nand g174757__9315 (n_8389, n_9257, n_8335);
  nor g174776__9945 (n_8388, n_1448, n_8332);
  nand g174702__2883 (n_8420, n_8413, n_8338);
  fflopd g3684_reg(.CK (clock), .D (n_8347), .Q (g3684));
  nor g174706__2346 (n_8458, n_6485, n_8387);
  nor g174703__1666 (n_8456, n_6248, n_8387);
  nor g174704__7410 (n_8461, n_6250, n_8387);
  nand g174368__6417 (n_8386, n_8355, n_8329);
  nor g174452__5477 (n_8385, n_8384, n_8362);
  nor g174459__2398 (n_8383, n_8382, n_8371);
  nand g174462__5107 (n_8381, n_1227, n_8330);
  nand g174464__6260 (n_8380, g28753, n_8327);
  nand g174351__4319 (n_8379, g28753, n_8326);
  not g174497 (n_8378, n_8354);
  not g174499 (n_8377, n_8376);
  not g174504 (n_8375, n_8374);
  not g174505 (n_8373, n_8372);
  fflopd g4427_reg(.CK (clock), .D (n_10286), .Q (g4427));
  nand g174546__8428 (n_8401, n_5270, n_8371);
  not g174740 (n_8370, n_8387);
  nand g174660__5526 (n_8369, n_7919, n_8324);
  not g174673 (n_8368, n_8339);
  nor g174719__6783 (n_8367, g301, g2902);
  nand g174626__3680 (n_8366, g4235, n_9257);
  not g174882 (n_8365, n_8337);
  nand g174750__1617 (n_8364, n_7882, n_8320);
  nand g174756__2802 (n_8363, g301, n_9257);
  nand g174547__1705 (n_8399, n_5023, n_8362);
  fflopd g160_reg(.CK (clock), .D (n_8321), .Q (g160));
  nand g174860__5122 (n_8415, g781, n_8325);
  fflopd g772_reg(.CK (clock), .D (n_8318), .Q (g772));
  not g174741 (n_8434, n_8343);
  not g174644 (n_8361, g4235);
  nor g174454__8246 (n_8360, n_8359, n_8345);
  nor g174457__7098 (n_8358, n_8357, n_8344);
  nand g174463__6131 (n_8356, n_8355, n_8308);
  nand g174531__1881 (n_8354, n_761, n_8316);
  nand g174533__5115 (n_8353, g3457, n_8313);
  nor g174453__7482 (n_8352, n_8351, n_8346);
  nand g174629__4733 (n_8350, g35, n_8310);
  nand g174628__6161 (n_8349, g35, n_8311);
  nor g174576__9315 (n_8348, n_8306, n_8125);
  nand g174577__9945 (n_8347, n_5394, n_8305);
  nand g174551__2883 (n_8372, n_5240, n_8346);
  nand g174550__2346 (n_8374, n_5011, n_8345);
  nand g174545__1666 (n_8376, n_5251, n_8344);
  nand g174766__7410 (n_8343, g35, n_8293);
  nand g174686__6417 (n_8342, n_8008, n_8300);
  nand g174690__5477 (n_8341, n_8314, n_9193);
  nand g174692__2398 (n_8340, n_8294, n_9193);
  nand g174697__5107 (n_8339, n_7848, n_8323);
  nor g174751__6260 (n_8338, new_g7558_, n_8295);
  nand g174910__4319 (n_8337, g781, n_8331);
  nor g174655__8428 (n_8336, g8920, n_8299);
  not g174767 (n_8335, g2759);
  nand g174886__5526 (n_8333, n_8904, n_8301);
  nor g174851__6783 (n_8332, g781, n_8331);
  fflopd g5084_reg(.CK (clock), .D (n_8309), .Q (g5084));
  nand g174765__3680 (n_8387, new_g7558_, n_8297);
  fflopd g1157_reg(.CK (clock), .D (n_10450), .Q (g7916));
  nand g174589__1617 (n_8330, n_5110, n_8289);
  wire w11, w12, w13, w14;
  nand g174520__2802 (n_8329, w12, w14);
  nand g17 (w14, w13, n_4289);
  not g16 (w13, n_8307);
  nand g15 (w12, w11, n_8307);
  not g14 (w11, n_4289);
  nor g174585__5122 (n_8327, g5115, n_8290);
  wire w15, w16, w17, w18;
  nand g174518__8246 (n_8326, w16, w18);
  nand g21 (w18, w17, n_4691);
  not g20 (w17, n_8315);
  nand g19 (w16, w15, n_8315);
  not g18 (w15, n_4691);
  nand g174597__7098 (n_8371, n_7281, n_8288);
  nand g174596__6131 (n_8362, n_7279, n_8291);
  fflopd g4235_reg(.CK (clock), .D (g8920), .Q (g4235));
  not g174924 (n_8325, n_8331);
  fflopd g2759_reg(.CK (clock), .D (n_8282), .Q (g2759));
  not g174739 (n_8324, n_8323);
  nor g174852__1881 (n_8322, n_1680, n_8281);
  nand g174814__5115 (n_8321, n_8258, n_8277);
  nor g174824__7482 (n_8320, n_8296, n_8319);
  nand g174839__4733 (n_8318, n_8257, n_8279);
  fflopd g301_reg(.CK (clock), .D (n_8278), .Q (g301));
  fflopd g106_reg(.CK (clock), .D (n_8284), .Q (g21176));
  nand g174664__6161 (n_8317, n_8312, n_8268);
  nand g174588__9315 (n_8316, n_5243, n_8315);
  not g174708 (n_8314, g4480);
  nand g174617__9945 (n_8313, n_8312, n_8269);
  nand g174696__2883 (n_8311, n_7731, n_8259);
  nand g174695__2346 (n_8310, n_7732, n_8276);
  nand g174663__1666 (n_8309, n_8117, n_8270);
  nor g174575__7410 (n_8308, g6154, n_8307);
  not g174674 (n_8306, n_8285);
  not g174675 (n_8305, n_8283);
  nand g174688__6417 (n_8304, g4578, n_8302);
  nand g174689__5477 (n_8303, g4575, n_8302);
  nand g174633__2398 (n_8345, n_6561, n_8274);
  nand g174631__5107 (n_8346, n_6581, n_8272);
  nand g174598__6260 (n_8344, n_7283, n_8273);
  not g174977 (n_8301, n_8286);
  nand g174753__4319 (n_8300, n_8262, n_8235);
  nand g174713__8428 (n_8299, n_8266, n_8251);
  nor g174780__6783 (n_8297, n_8296, n_8254);
  nand g174784__3680 (n_8295, n_8296, n_8292);
  not g174709 (n_8294, g4540);
  nand g174822__1617 (n_8293, new_g7558_, n_8292);
  nand g174764__2802 (n_8323, n_8263, n_8234);
  nand g174956__1705 (n_8331, g776, n_8275);
  fflopd g1036_reg(.CK (clock), .D (n_8260), .Q (g1036));
  fflopd g157_reg(.CK (clock), .D (n_8267), .Q (g157));
  fflopd g142_reg(.CK (clock), .D (n_8264), .Q (g142));
  fflopd g767_reg(.CK (clock), .D (n_8265), .Q (g767));
  fflopd g1061_reg(.CK (clock), .D (n_8271), .Q (g1061));
  nor g174661__5122 (n_8291, n_6990, n_10290);
  not g174643 (n_8290, n_8315);
  not g174645 (n_8289, n_8307);
  nor g174646__8246 (n_8288, n_6993, n_10288);
  nand g175024__6131 (n_8286, g776, n_8280);
  nand g174699__1881 (n_8285, g35, n_8244);
  nand g174700__5115 (n_8284, n_827, n_8243);
  nand g174701__7482 (n_8283, n_852, n_8247);
  fflopd g4480_reg(.CK (clock), .D (n_8245), .Q (g4480));
  fflopd g4540_reg(.CK (clock), .D (n_8242), .Q (g4540));
  nand g174894__4733 (n_8282, n_9257, n_8239);
  nor g174938__6161 (n_8281, g776, n_8280);
  nand g175006__9315 (n_8279, n_8904, n_8252);
  not g174881 (n_8278, n_8255);
  nand g174842__9945 (n_8277, n_8214, n_8240);
  not g174838 (n_8319, n_8292);
  fflopd g1105_reg(.CK (clock), .D (n_8236), .Q (g1105));
  fflopd g4232_reg(.CK (clock), .D (g8919), .Q (g8920));
  fflopd g1379_reg(.CK (clock), .D (n_8237), .Q (g1379));
  fflopd g1129_reg(.CK (clock), .D (n_10258), .Q (g1129));
  fflopd g1135_reg(.CK (clock), .D (n_10256), .Q (g1135));
  nand g174758__2883 (n_8276, n_8209, n_8007);
  not g175035 (n_8275, n_8280);
  nor g174651__2346 (n_8274, n_5299, n_8223);
  nor g174653__1666 (n_8273, n_6998, n_10128);
  nor g174662__7410 (n_8272, n_5487, n_8221);
  nand g174748__6417 (n_8271, n_8193, n_8210);
  not g174736 (n_8270, n_8253);
  wire w19, w20, w21, w22;
  nand g174685__5477 (n_8269, w20, w22);
  nand g25 (w22, w21, n_4692);
  not g24 (w21, n_8246);
  nand g23 (w20, w19, n_8246);
  not g22 (w19, n_4692);
  fflopd g4578_reg(.CK (clock), .D (n_8211), .Q (g4578));
  nor g174717__2398 (n_8268, g3457, n_8218);
  fflopd g4575_reg(.CK (clock), .D (n_8212), .Q (g4575));
  nor g174669__5107 (n_8307, n_7867, n_8222);
  nand g174667__6260 (n_8315, n_6563, n_8225);
  fflopd g1570_reg(.CK (clock), .D (n_8213), .Q (g12923));
  nand g174843__4319 (n_8267, n_8215, n_8180);
  not g174769 (n_8266, g8919);
  nand g175005__8428 (n_8265, n_8228, n_8199);
  nand g174805__5526 (n_8264, n_8204, n_8192);
  nand g174812__6783 (n_8263, n_3256, n_8261);
  nand g174816__3680 (n_8262, n_8074, n_8261);
  nand g174820__1617 (n_8260, n_7964, n_8206);
  nand g174759__2802 (n_8259, n_8015, n_8208);
  nor g174845__1705 (n_8258, n_1451, n_8205);
  nor g174927__5122 (n_8257, n_1447, n_8229);
  nand g174905__8246 (n_8255, g160, n_8217);
  nand g174906__7098 (n_8254, new_g6856_, new_g7586_);
  nor g174869__6131 (n_8292, new_g6856_, new_g7586_);
  fflopd g4950_reg(.CK (clock), .D (n_8220), .Q (g4950));
  nand g174749__1881 (n_8253, n_7735, n_8194);
  not g175122 (n_8252, n_8227);
  nor g174778__5115 (n_8251, g8918, n_10301);
  nand g174747__6161 (n_8247, n_8166, n_8246);
  nand g174777__9315 (n_8245, n_2299, n_8241);
  nor g174752__9945 (n_8244, g311, n_8196);
  nand g174761__2883 (n_8243, g35, n_8200);
  nand g174773__2346 (n_8242, n_4482, n_8241);
  fflopd g4430_reg(.CK (clock), .D (n_8195), .Q (g4430));
  fflopd g4229_reg(.CK (clock), .D (g8918), .Q (g8919));
  nand g175096__1666 (n_8280, g772, n_8202);
  fflopd g1052_reg(.CK (clock), .D (n_8197), .Q (g1052));
  not g174983 (n_8240, n_8230);
  not g174925 (n_8239, new_g6856_);
  nand g174895__6417 (n_8237, n_8139, n_8177);
  nand g174819__5477 (n_8236, n_8160, n_8190);
  nand g174815__2398 (n_8235, g1135, n_8233);
  nand g174811__5107 (n_8234, g956, n_8233);
  fflopd g1874_reg(.CK (clock), .D (n_8178), .Q (g1874));
  fflopd g1978_reg(.CK (clock), .D (n_8179), .Q (g1978));
  fflopd g1146_reg(.CK (clock), .D (n_8187), .Q (g1146));
  fflopd g153_reg(.CK (clock), .D (n_8186), .Q (g153));
  fflopd g763_reg(.CK (clock), .D (n_8198), .Q (g763));
  fflopd g298_reg(.CK (clock), .D (n_8183), .Q (g298));
  fflopd g890_reg(.CK (clock), .D (n_8184), .Q (g890));
  nand g175031__8428 (n_8230, g160, n_8216);
  nor g175044__5526 (n_8229, g772, n_8226);
  nand g175160__6783 (n_8228, n_8904, n_8174);
  nand g175194__3680 (n_8227, g772, n_8226);
  nor g174714__1617 (n_8225, n_7940, n_10297);
  nand g174718__1705 (n_8223, n_4771, n_10295);
  nand g174744__5122 (n_8222, n_7072, n_8168);
  nand g174746__8246 (n_8221, n_4678, n_10299);
  nand g174760__7098 (n_8220, n_5387, n_8167);
  nand g174762__6131 (n_8219, g35, n_8165);
  not g174771 (n_8218, n_8246);
  nand g175016__1881 (n_8217, g35, n_8216);
  fflopd g1373_reg(.CK (clock), .D (n_8147), .Q (g1373));
  nand g174998__5115 (n_8215, n_8214, n_8170);
  nand g174823__7482 (n_8213, n_8155, n_786);
  nand g174828__4733 (n_8212, n_8162, n_8011);
  nand g174829__6161 (n_8211, n_8161, n_8009);
  nand g174832__9315 (n_8210, g1061, n_8163);
  wire w23, w24, w25, w26;
  nand g174834__9945 (n_8209, w24, w26);
  nand g29 (w26, w25, g1105);
  not g28 (w25, n_8207);
  nand g27 (w24, w23, n_8207);
  not g26 (w23, g1105);
  wire w27, w28, w29, w30;
  nand g174835__2883 (n_8208, w28, w30);
  nand g33 (w30, w29, g1129);
  not g32 (w29, n_8207);
  nand g31 (w28, w27, n_8207);
  not g30 (w27, g1129);
  not g174883 (n_8206, n_8182);
  nor g174988__2346 (n_8205, g160, n_8216);
  nand g174898__1666 (n_8204, n_8107, n_8148);
  not g174885 (n_8261, n_8181);
  fflopd g2756_reg(.CK (clock), .D (n_8175), .Q (new_g6856_));
  fflopd g1982_reg(.CK (clock), .D (n_8151), .Q (g1982));
  fflopd g1030_reg(.CK (clock), .D (n_8169), .Q (g1030));
  not g175216 (n_8202, n_8226);
  nor g174782__5477 (n_8200, n_8123, n_5175);
  nor g175047__2398 (n_8199, n_1475, n_8134);
  nand g175159__5107 (n_8198, n_8080, n_8133);
  nand g174808__6260 (n_8197, n_10134, n_8119);
  nand g174813__4319 (n_8196, n_2163, n_8124);
  nand g174826__8428 (n_8195, n_378, n_8118);
  nand g174830__5526 (n_8194, n_7502, n_8130);
  nand g174831__6783 (n_8193, g1052, n_8120);
  fflopd g1882_reg(.CK (clock), .D (n_8137), .Q (g1882));
  fflopd g1878_reg(.CK (clock), .D (n_8138), .Q (g1878));
  fflopd g1710_reg(.CK (clock), .D (n_8112), .Q (g1710));
  fflopd g4704_reg(.CK (clock), .D (n_8128), .Q (g4704));
  nand g174797__3680 (n_8246, n_7284, n_8122);
  fflopd g4939_reg(.CK (clock), .D (n_8114), .Q (g4939));
  fflopd g4961_reg(.CK (clock), .D (n_8113), .Q (g4961));
  fflopd g1604_reg(.CK (clock), .D (n_8111), .Q (g1604));
  nor g174850__1617 (n_8192, n_1479, n_8106);
  not g174876 (n_8190, n_8159);
  not g174879 (n_8187, n_8156);
  nand g174997__1705 (n_8186, n_8096, n_8140);
  nand g174892__5122 (n_8185, g35, n_8110);
  nand g174896__8246 (n_8184, n_2026, n_8105);
  nand g174897__7098 (n_8183, n_8066, n_8108);
  nand g174920__6131 (n_8182, n_702, n_8145);
  nand g174922__1881 (n_8181, g35, n_8207);
  nor g174987__5115 (n_8180, n_1521, n_8144);
  nand g174931__7482 (n_8179, n_1263, n_8141);
  nand g174940__4733 (n_8178, n_7780, n_8142);
  not g174975 (n_8177, n_8171);
  not g174884 (n_8241, n_8153);
  nor g174923__6161 (n_8233, n_9257, n_8207);
  fflopd g4226_reg(.CK (clock), .D (g8870), .Q (g8918));
  fflopd g956_reg(.CK (clock), .D (n_8127), .Q (g956));
  nand g175163__9315 (n_8175, n_9257, n_8082);
  not g175360 (n_8174, n_8132);
  nand g175017__2346 (n_8171, n_550, n_8091);
  not g175127 (n_8170, n_8136);
  nand g175286__1666 (n_8226, g767, n_8078);
  fflopd g4894_reg(.CK (clock), .D (n_8057), .Q (g4894));
  fflopd g4760_reg(.CK (clock), .D (n_8077), .Q (g4760));
  fflopd g4771_reg(.CK (clock), .D (n_8059), .Q (g4771));
  fflopd g4749_reg(.CK (clock), .D (n_8061), .Q (g4749));
  nand g175079__7410 (n_8216, g157, n_8081);
  fflopd g1870_reg(.CK (clock), .D (n_10420), .Q (g1870));
  fflopd g1886_reg(.CK (clock), .D (n_8090), .Q (g1886));
  fflopd g1152_reg(.CK (clock), .D (n_8100), .Q (g1152));
  fflopd g1955_reg(.CK (clock), .D (n_8085), .Q (g1955));
  fflopd g1974_reg(.CK (clock), .D (n_8084), .Q (g1974));
  fflopd g150_reg(.CK (clock), .D (n_8089), .Q (g150));
  fflopd g758_reg(.CK (clock), .D (n_8079), .Q (g758));
  fflopd g1099_reg(.CK (clock), .D (n_8088), .Q (g1099));
  fflopd g1714_reg(.CK (clock), .D (n_8060), .Q (g1714));
  nand g175010__6417 (n_8169, n_7965, n_8092);
  nor g174821__5477 (n_8168, n_5892, n_8058);
  nand g174833__2398 (n_8167, n_8062, n_8166);
  wire w31, w32, w33, w34;
  nand g174836__5107 (n_8165, w32, w34);
  nand g40 (w34, w33, g4434);
  not g39 (w33, g4401);
  nand g38 (w32, w31, g4401);
  not g34 (w31, g4434);
  nand g174840__6260 (n_8164, g4572, n_8302);
  nand g174841__4319 (n_8163, n_1998, n_8068);
  nand g174889__8428 (n_8162, g20049, n_9257);
  nand g174890__5526 (n_8161, g4572, n_9257);
  nand g174893__6783 (n_8160, g35, n_8072);
  nand g174900__3680 (n_8159, n_819, n_8071);
  nand g174901__1617 (n_8158, n_1250, n_8073);
  nand g174902__2802 (n_8157, n_1193, n_8075);
  nand g174903__1705 (n_8156, g35, n_8101);
  nand g174907__5122 (n_8155, g35, g496);
  nand g174911__8246 (n_8154, g20049, new_g10233_);
  nand g174921__7098 (n_8153, n_8099, n_9193);
  not g174926 (n_8152, g8870);
  nand g174929__6131 (n_8151, n_7987, n_8093);
  not g174980 (n_8148, n_8146);
  nand g175009__7482 (n_8147, n_7988, n_8094);
  fflopd g294_reg(.CK (clock), .D (n_8076), .Q (g294));
  nand g175027__4733 (n_8146, g142, n_8109);
  nand g175032__6161 (n_8145, n_7889, n_8035);
  nor g175037__9315 (n_8144, g157, n_8135);
  not g175121 (n_8142, n_8086);
  not g175123 (n_8141, n_8083);
  nand g175153__9945 (n_8140, n_8214, n_8053);
  nand g175165__2883 (n_8139, g35, n_8032);
  nand g175170__2346 (n_8138, n_8033, n_7944);
  nand g175171__1666 (n_8137, n_8052, n_7968);
  nand g175203__7410 (n_8136, g157, n_8135);
  nor g175237__6417 (n_8134, g767, n_8131);
  nand g175410__5477 (n_8133, n_8904, n_8031);
  nand g175473__2398 (n_8132, g767, n_8131);
  nor g174844__5107 (n_8130, g5080, n_8116);
  nand g174825__6260 (n_8129, n_4813, n_8025);
  fflopd g2112_reg(.CK (clock), .D (n_8054), .Q (g2112));
  fflopd g1950_reg(.CK (clock), .D (n_8034), .Q (g1950));
  fflopd g164_reg(.CK (clock), .D (n_10422), .Q (g164));
  fflopd g1024_reg(.CK (clock), .D (n_8039), .Q (g1024));
  fflopd g1608_reg(.CK (clock), .D (n_8056), .Q (g1608));
  fflopd g1612_reg(.CK (clock), .D (n_8040), .Q (g1612));
  fflopd g1367_reg(.CK (clock), .D (n_8042), .Q (g1367));
  fflopd g1906_reg(.CK (clock), .D (n_8026), .Q (g1906));
  nand g174912__4319 (n_8128, n_5391, n_10304);
  nand g174848__8428 (n_8127, n_8041, n_8048);
  nand g174849__5526 (n_8126, n_7639, n_8021);
  nor g174853__6783 (n_8125, n_8023, n_5695);
  nor g174854__3680 (n_8124, g329, g319);
  nand g174856__1617 (n_8123, g329, n_7768);
  nor g174857__2802 (n_8122, n_7942, n_10309);
  nand g174888__1705 (n_8121, g329, n_9257);
  nand g174891__5122 (n_8120, g35, n_8029);
  nand g174899__8246 (n_8119, g35, n_8067);
  nand g174908__7098 (n_8118, g4434, n_6995);
  nand g174909__6131 (n_8117, g5080, n_8116);
  nand g174847__1881 (n_8115, n_7636, n_8022);
  nand g174918__5115 (n_8114, n_5449, n_10307);
  nand g174919__7482 (n_8113, n_5451, n_8027);
  nand g174930__4733 (n_8112, n_916, n_8049);
  nand g174934__6161 (n_8111, n_7591, n_8050);
  nor g174937__9315 (n_8110, n_63, n_8109);
  nand g175012__9945 (n_8108, n_8107, n_8051);
  nor g175004__2883 (n_8106, g142, n_8109);
  not g174979 (n_8105, n_8098);
  fflopd g4222_reg(.CK (clock), .D (g8917), .Q (g8870));
  nor g174974__7410 (n_8207, g976, n_2502);
  nand g175014__5477 (n_8101, n_7811, n_7999);
  nand g175015__2398 (n_8100, n_7918, n_8004);
  nand g175023__5107 (n_8099, g35, new_g8880_);
  nand g175026__6260 (n_8098, n_1256, n_8017);
  nor g175038__4319 (n_8096, n_1466, n_7985);
  not g175116 (n_8094, n_8038);
  not g175124 (n_8093, n_8037);
  not g175128 (n_8092, n_8036);
  nand g175136__5526 (n_8091, n_7901, n_7986);
  nand g175137__6783 (n_8090, n_6919, n_7977);
  nand g175152__3680 (n_8089, n_7974, n_7907);
  nand g175013__1617 (n_8088, n_7920, n_8005);
  nand g175191__1705 (n_8086, n_1230, n_7973);
  nand g175193__5122 (n_8085, n_7893, n_7972);
  nand g175195__8246 (n_8084, n_7892, n_7971);
  nand g175196__7098 (n_8083, n_7796, n_7979);
  not g175213 (n_8082, new_g7586_);
  not g175214 (n_8081, n_8135);
  nor g175238__6131 (n_8080, n_1641, n_7956);
  nand g175409__1881 (n_8079, n_7954, n_7881);
  not g175513 (n_8078, n_8131);
  fflopd g1748_reg(.CK (clock), .D (n_8016), .Q (g1748));
  fflopd g1687_reg(.CK (clock), .D (n_7993), .Q (g1687));
  fflopd g1706_reg(.CK (clock), .D (n_7992), .Q (g1706));
  fflopd g1227_reg(.CK (clock), .D (n_7998), .Q (g12919));
  nand g174914__5115 (n_8077, n_5443, n_10321);
  nand g175011__7482 (n_8076, n_8000, n_7936);
  nand g175002__4733 (n_8075, n_8074, n_8046);
  nand g175001__6161 (n_8073, n_5368, n_8044);
  nor g174996__9315 (n_8072, n_8069, n_8070);
  nand g174995__9945 (n_8071, n_8069, n_8070);
  not g174984 (n_8068, n_8067);
  nor g174936__2883 (n_8066, n_1469, n_8014);
  fflopd g496_reg(.CK (clock), .D (n_7995), .Q (g496));
  nor g174887__6417 (n_8062, n_3376, n_7947);
  nand g174913__5477 (n_8061, n_5442, n_10312);
  nand g174928__2398 (n_8060, n_7835, n_8013);
  nand g174915__5107 (n_8059, n_5390, n_7950);
  nand g174916__6260 (n_8058, n_7280, n_7946);
  nand g174917__4319 (n_8057, n_5447, n_10318);
  fflopd g4572_reg(.CK (clock), .D (n_8010), .Q (g4572));
  fflopd g1752_reg(.CK (clock), .D (n_7981), .Q (g1752));
  fflopd g1600_reg(.CK (clock), .D (n_10424), .Q (g1600));
  fflopd g1744_reg(.CK (clock), .D (n_7980), .Q (g1744));
  fflopd g1736_reg(.CK (clock), .D (n_8020), .Q (g1736));
  fflopd g1890_reg(.CK (clock), .D (n_7967), .Q (g1890));
  fflopd g2016_reg(.CK (clock), .D (n_7966), .Q (g2016));
  fflopd g2084_reg(.CK (clock), .D (n_10138), .Q (g2084));
  fflopd g59_reg(.CK (clock), .D (n_8012), .Q (g20049));
  fflopd g2116_reg(.CK (clock), .D (n_7984), .Q (g2116));
  fflopd g5052_reg(.CK (clock), .D (n_7955), .Q (g5052));
  nand g175167__8428 (n_8056, n_7932, n_7826);
  fflopd g976_reg(.CK (clock), .D (n_10260), .Q (g976));
  nand g175042__6783 (n_8054, n_7575, n_7884);
  not g175364 (n_8053, n_7958);
  not g175358 (n_8052, n_7959);
  not g175115 (n_8051, n_7997);
  not g175117 (n_8050, n_7994);
  not g175118 (n_8049, n_7991);
  not g175125 (n_8048, n_7990);
  nand g175155__3680 (n_8043, n_10327, n_5916);
  nand g175164__1617 (n_8042, n_7719, n_7930);
  nand g175028__2802 (n_8041, g956, n_7914);
  nand g175168__1705 (n_8040, n_7943, n_7825);
  nand g175173__5122 (n_8039, n_7691, n_7903);
  nand g175182__8246 (n_8038, n_1058, n_7902);
  nand g175197__7098 (n_8037, n_658, n_7897);
  nand g175204__6131 (n_8036, n_662, n_7890);
  nand g175205__1881 (n_8035, n_1975, n_7888);
  nand g175223__5115 (n_8034, n_7548, n_7887);
  not g175357 (n_8033, n_7960);
  not g175349 (n_8032, n_7963);
  nor g175033__7482 (n_8067, g979, n_7923);
  fflopd g2748_reg(.CK (clock), .D (n_7883), .Q (new_g7586_));
  nand g175268__4733 (n_8135, g153, n_7886);
  nand g175058__6161 (n_8109, g298, n_7910);
  fflopd g4219_reg(.CK (clock), .D (g8916), .Q (g8917));
  not g175706 (n_8031, n_7953);
  nand g175003__9945 (n_8029, n_2503, n_7924);
  nand g174991__2346 (n_8027, n_7925, n_5338);
  nand g175434__1666 (n_8026, n_7549, n_7885);
  nor g174859__7410 (n_8025, n_7506, n_7941);
  nor g174935__5477 (n_8023, g319, n_4664);
  not g174981 (n_8022, n_8018);
  not g174978 (n_8021, n_8019);
  fflopd g4434_reg(.CK (clock), .D (n_7937), .Q (g4434));
  fflopd g5080_reg(.CK (clock), .D (n_7913), .Q (g5080));
  nand g175632__2398 (n_8131, g763, n_7912);
  fflopd g4446_reg(.CK (clock), .D (n_7938), .Q (g7245));
  fflopd g2403_reg(.CK (clock), .D (n_7928), .Q (g2403));
  fflopd g2671_reg(.CK (clock), .D (n_7935), .Q (g2671));
  fflopd g146_reg(.CK (clock), .D (n_7895), .Q (g146));
  fflopd g1682_reg(.CK (clock), .D (n_7909), .Q (g1682));
  fflopd g2008_reg(.CK (clock), .D (n_7900), .Q (g2008));
  fflopd g1844_reg(.CK (clock), .D (n_7906), .Q (g1844));
  fflopd g2004_reg(.CK (clock), .D (n_10426), .Q (g2004));
  fflopd g329_reg(.CK (clock), .D (g319), .Q (g329));
  fflopd g1740_reg(.CK (clock), .D (n_7911), .Q (g1740));
  fflopd g1756_reg(.CK (clock), .D (n_7905), .Q (g1756));
  fflopd g291_reg(.CK (clock), .D (n_7921), .Q (g291));
  fflopd g749_reg(.CK (clock), .D (n_7904), .Q (g749));
  fflopd g714_reg(.CK (clock), .D (n_7916), .Q (new_g10354_));
  fflopd g1636_reg(.CK (clock), .D (n_7898), .Q (g1636));
  nand g175429__5107 (n_8020, n_7714, n_7810);
  nand g175025__6260 (n_8019, n_4124, n_7871);
  nand g175029__4319 (n_8018, n_4123, n_7870);
  nand g175041__8428 (n_8017, n_1948, n_7858);
  fflopd g4372_reg(.CK (clock), .D (n_7862), .Q (new_g8880_));
  nand g175049__5526 (n_8016, n_7189, n_7856);
  nand g175051__6783 (n_8015, n_104, n_7843);
  nor g175053__3680 (n_8014, g298, n_7996);
  not g175119 (n_8013, n_7917);
  not g175130 (n_8012, n_8011);
  not g175131 (n_8010, n_8009);
  nand g175135__1617 (n_8008, n_216, n_7845);
  nand g175138__2802 (n_8007, n_199, n_7850);
  nand g175150__5122 (n_8005, g1099, n_8003);
  nand g175151__8246 (n_8004, g1152, n_8003);
  nand g175174__6131 (n_8001, g35, n_7855);
  nand g175176__1881 (n_8000, n_8107, n_7857);
  nand g175178__5115 (n_7999, g1146, n_7852);
  nand g175180__7482 (n_7998, n_7819, n_1202);
  nand g175181__4733 (n_7997, g298, n_7996);
  nand g175183__6161 (n_7995, n_330, n_7834);
  nand g175184 (n_7994, n_1306, n_7840);
  nand g175185 (n_7993, n_7728, n_7839);
  nand g175186 (n_7992, n_7727, n_7837);
  nand g175187 (n_7991, n_7587, n_7836);
  nand g175201 (n_7990, n_1273, n_7847);
  nand g175022 (n_7989, n_5354, n_7868);
  nand g175418 (n_7988, g35, n_7795);
  nand g175401 (n_7987, g1982, n_7978);
  nor g175225 (n_7986, g1379, n_7962);
  nor g175230 (n_7985, g153, n_7957);
  nand g175235 (n_7984, n_7239, n_7788);
  nand g175244 (n_7981, n_688, n_7808);
  nand g175245 (n_7980, n_547, n_7809);
  nand g175400 (n_7979, g1978, n_7978);
  not g175359 (n_7977, n_7894);
  nand g175386 (n_7974, n_8214, n_7787);
  nand g175397 (n_7973, g1874, n_7978);
  nand g175398 (n_7972, g1955, n_7978);
  nand g175399 (n_7971, g1974, n_7978);
  nor g175210 (n_8044, n_7970, n_7842);
  nor g175211 (n_8070, n_7970, n_7865);
  nor g175207 (n_8046, n_7970, n_7846);
  fflopd g2675_reg(.CK (clock), .D (n_7860), .Q (g2675));
  nand g175432 (n_7968, g35, n_7793);
  nand g175433 (n_7967, n_7686, n_7792);
  nand g175437 (n_7966, n_7694, n_7791);
  nand g175440 (n_7965, g35, n_7786);
  nand g175441 (n_7964, g35, n_7785);
  nand g175454 (n_7963, g1379, n_7962);
  nand g175469 (n_7960, n_698, n_7800);
  nand g175470 (n_7959, n_1128, n_7799);
  nand g175487 (n_7958, g153, n_7957);
  nor g175566 (n_7956, g763, n_7952);
  nand g175572 (n_7955, n_7328, n_7812);
  nand g175580 (n_7954, n_8904, n_7797);
  nand g175815 (n_7953, g763, n_7952);
  nand g174992 (n_7950, n_7873, n_5397);
  nor g174986 (n_7947, g4950, n_7879);
  nand g174985 (n_7946, n_4492, n_7872);
  nand g175431 (n_7944, g35, n_7794);
  fflopd g2429_reg(.CK (clock), .D (n_7833), .Q (g2429));
  fflopd g2307_reg(.CK (clock), .D (n_7820), .Q (g2307));
  fflopd g2575_reg(.CK (clock), .D (n_7832), .Q (g2575));
  fflopd g1620_reg(.CK (clock), .D (n_7823), .Q (g1620));
  fflopd g2441_reg(.CK (clock), .D (n_7877), .Q (g2441));
  fflopd g1437_reg(.CK (clock), .D (n_7830), .Q (g1437));
  fflopd g1454_reg(.CK (clock), .D (n_7829), .Q (g1454));
  fflopd g1018_reg(.CK (clock), .D (n_7821), .Q (g1018));
  fflopd g1616_reg(.CK (clock), .D (n_7824), .Q (g1616));
  fflopd g854_reg(.CK (clock), .D (n_7789), .Q (g854));
  fflopd g1816_reg(.CK (clock), .D (n_7804), .Q (g1816));
  fflopd g1467_reg(.CK (clock), .D (n_7828), .Q (g1467));
  fflopd g2161_reg(.CK (clock), .D (n_7822), .Q (g2161));
  fflopd g2173_reg(.CK (clock), .D (n_7878), .Q (g2173));
  fflopd g1728_reg(.CK (clock), .D (n_7805), .Q (g1728));
  fflopd g4593_reg(.CK (clock), .D (n_7782), .Q (g4593));
  fflopd g2643_reg(.CK (clock), .D (n_10142), .Q (g2643));
  fflopd g1862_reg(.CK (clock), .D (n_7802), .Q (g1862));
  fflopd g5057_reg(.CK (clock), .D (n_7803), .Q (g5057));
  fflopd g2375_reg(.CK (clock), .D (n_10144), .Q (g2375));
  fflopd g1592_reg(.CK (clock), .D (n_7817), .Q (g1592));
  fflopd g2407_reg(.CK (clock), .D (n_7864), .Q (g2407));
  fflopd g1361_reg(.CK (clock), .D (n_7831), .Q (g1361));
  fflopd g1848_reg(.CK (clock), .D (n_7861), .Q (g1848));
  fflopd g1936_reg(.CK (clock), .D (n_7777), .Q (g1936));
  fflopd g2040_reg(.CK (clock), .D (n_7781), .Q (g2040));
  fflopd g1772_reg(.CK (clock), .D (n_7801), .Q (g1772));
  not g175353 (n_7943, n_7815);
  nand g175019 (n_7942, n_6318, n_7771);
  nand g175020 (n_7941, n_7309, n_7770);
  nand g175021 (n_7940, n_3699, n_7772);
  nand g175030 (n_7939, n_4126, n_7773);
  nand g175043 (n_7938, n_5792, n_7752);
  nand g175046 (n_7937, n_1138, n_7766);
  nor g175052 (n_7936, n_1661, n_7761);
  nand g175054 (n_7935, n_7287, n_7755);
  nand g175018 (n_7933, n_4122, n_7769);
  not g175352 (n_7932, n_7816);
  not g175348 (n_7930, n_7818);
  nand g175134 (n_7928, n_7265, n_7751);
  nand g175139 (n_7927, n_206, n_7767);
  nand g175143 (n_7926, n_145, n_7740);
  nand g175144 (n_7925, n_214, n_7750);
  nor g175149 (n_7924, g1061, n_7922);
  nand g175172 (n_7923, g1052, n_7922);
  nand g175175 (n_7921, n_7661, n_7733);
  nand g175177 (n_7920, g1152, n_7919);
  nand g175179 (n_7918, g1146, n_7919);
  nand g175188 (n_7917, n_727, n_7738);
  nand g175189 (n_7916, n_7113, n_7724);
  nand g175198 (n_7915, g35, n_7723);
  nand g175200 (n_7914, n_7919, n_2782);
  nand g175206 (n_7913, n_7746, n_7269);
  not g175906 (n_7912, n_7952);
  nand g175246 (n_7911, n_6950, n_7702);
  not g175215 (n_7910, n_7996);
  nand g175224 (n_7909, n_7201, n_7703);
  nor g175232 (n_7907, n_535, n_7674);
  nand g175242 (n_7906, n_1221, n_7700);
  nand g175243 (n_7905, n_7583, n_7701);
  nand g175209 (n_8009, g35, n_7742);
  nand g175208 (n_8011, g35, n_7743);
  fflopd g319_reg(.CK (clock), .D (n_7762), .Q (g319));
  fflopd g2563_reg(.CK (clock), .D (n_10428), .Q (g2563));
  fflopd g2020_reg(.CK (clock), .D (n_7716), .Q (g2020));
  fflopd g2299_reg(.CK (clock), .D (n_7745), .Q (g2299));
  fflopd g4216_reg(.CK (clock), .D (g8915), .Q (g8916));
  nand g175603 (n_7904, n_7552, n_7672);
  not g175365 (n_7903, n_7813);
  nand g175380 (n_7902, n_7901, n_7711);
  nand g175385 (n_7900, n_6929, n_7699);
  nand g175427 (n_7898, n_7202, n_7704);
  nand g175435 (n_7897, g35, n_7757);
  nand g175836 (n_7895, n_1141, n_7774);
  nand g175471 (n_7894, n_743, n_7697);
  nand g175472 (n_7893, g1950, n_7891);
  nand g175476 (n_7892, g1968, n_7891);
  nand g175489 (n_7890, n_7889, n_7708);
  nand g175490 (n_7888, g1030, n_7710);
  not g175705 (n_7887, n_7783);
  not g175511 (n_7886, n_7957);
  not g175703 (n_7885, n_7778);
  not g175362 (n_7884, n_7853);
  nor g175538 (n_7883, g35, n_7882);
  nor g175565 (n_7881, n_1535, n_7706);
  fflopd g287_reg(.CK (clock), .D (n_7734), .Q (g287));
  fflopd g2449_reg(.CK (clock), .D (n_7776), .Q (g2449));
  fflopd g2567_reg(.CK (clock), .D (n_7747), .Q (g2567));
  fflopd g2169_reg(.CK (clock), .D (n_7763), .Q (g2169));
  fflopd g2181_reg(.CK (clock), .D (n_7741), .Q (g2181));
  fflopd g2433_reg(.CK (clock), .D (n_7749), .Q (g2433));
  fflopd g2295_reg(.CK (clock), .D (n_10430), .Q (g2295));
  fflopd g2437_reg(.CK (clock), .D (n_7758), .Q (g2437));
  fflopd g2537_reg(.CK (clock), .D (n_7760), .Q (g2537));
  fflopd g2165_reg(.CK (clock), .D (n_7748), .Q (g2165));
  fflopd g2269_reg(.CK (clock), .D (n_7765), .Q (g2269));
  fflopd g6163_reg(.CK (clock), .D (n_7720), .Q (g6163));
  fflopd g6177_reg(.CK (clock), .D (n_7721), .Q (g6177));
  fflopd g2012_reg(.CK (clock), .D (n_7695), .Q (g2012));
  fflopd g2024_reg(.CK (clock), .D (n_7692), .Q (g2024));
  fflopd g3466_reg(.CK (clock), .D (n_7737), .Q (g3466));
  fflopd g3480_reg(.CK (clock), .D (n_7756), .Q (g3480));
  fflopd g5124_reg(.CK (clock), .D (n_7715), .Q (g5124));
  fflopd g5138_reg(.CK (clock), .D (n_7717), .Q (g5138));
  fflopd g2445_reg(.CK (clock), .D (n_7759), .Q (g2445));
  fflopd g2177_reg(.CK (clock), .D (n_7764), .Q (g2177));
  fflopd g4616_reg(.CK (clock), .D (n_7684), .Q (new_g10383_));
  nand g175039 (n_7879, n_7324, n_7635);
  nand g175040 (n_7878, n_6763, n_7652);
  nand g175050 (n_7877, n_6788, n_7654);
  nand g175140 (n_7876, n_161, n_7665);
  nand g175141 (n_7875, n_148, n_7666);
  nand g175142 (n_7874, n_129, n_7667);
  nand g175145 (n_7873, n_44, n_7650);
  nand g175156 (n_7872, n_6508, n_7637);
  nand g175157 (n_7871, n_6359, n_7649);
  nand g175158 (n_7870, n_6357, n_7648);
  nand g175190 (n_7869, n_4179, n_7642);
  nand g175192 (n_7868, g25219, n_7633);
  nand g175199 (n_7867, n_4125, n_7638);
  nand g175202 (n_7866, g6727, n_7651);
  nand g175222 (n_7865, g1111, n_7849);
  nand g175226 (n_7864, n_6836, n_7595);
  nand g175239 (n_7862, n_7659, n_7183);
  nand g175241 (n_7861, n_7233, n_7658);
  nand g175247 (n_7860, n_6809, n_7604);
  nand g175481 (n_7858, g896, n_7574);
  not g175346 (n_7857, n_7730);
  not g175355 (n_7856, n_7725);
  not g175366 (n_7855, n_7722);
  nand g175479 (n_7853, n_7238, n_7572);
  nand g175378 (n_7852, g1152, n_7851);
  nand g175379 (n_7850, n_7848, n_7849);
  nand g175381 (n_7847, n_7851, n_2871);
  nand g175382 (n_7846, g1094, n_7844);
  nand g175383 (n_7845, n_7848, n_7844);
  nand g175390 (n_7843, n_7848, n_7841);
  nand g175391 (n_7842, g1124, n_7841);
  nand g175392 (n_7840, g1604, n_7838);
  nand g175393 (n_7839, g1687, n_7838);
  nand g175394 (n_7837, g1706, n_7838);
  nand g175395 (n_7836, g1710, n_7838);
  nand g175396 (n_7835, g1714, n_7838);
  nand g175413 (n_7834, g20901, n_9257);
  nand g175414 (n_7833, n_7491, n_7607);
  nand g175416 (n_7832, n_7494, n_7606);
  nand g175417 (n_7831, n_7392, n_7608);
  nand g175419 (n_7830, n_7497, n_7625);
  nand g175420 (n_7829, n_7498, n_7626);
  nand g175421 (n_7828, n_7499, n_7628);
  nand g175423 (n_7826, g35, n_7629);
  nand g175424 (n_7825, g35, n_7630);
  nand g175425 (n_7824, n_7500, n_7647);
  nand g175426 (n_7823, n_7501, n_7655);
  nand g175438 (n_7822, n_7457, n_7563);
  nand g175439 (n_7821, n_7386, n_7598);
  nand g175444 (n_7820, n_7454, n_7597);
  nand g175450 (n_7819, g35, g20901);
  nand g175453 (n_7818, n_531, n_7592);
  nand g175457 (n_7817, n_7327, n_7624);
  nand g175459 (n_7816, n_1022, n_7613);
  nand g175460 (n_7815, n_672, n_7612);
  nand g175467 (n_7814, n_826, n_7579);
  not g175370 (n_8003, n_7919);
  nand g175278 (n_7996, g294, n_7627);
  nand g175488 (n_7813, n_571, n_7614);
  not g176244 (n_7812, n_7775);
  nand g175494 (n_7811, n_88, n_7851);
  not g175499 (n_7810, n_7693);
  not g175500 (n_7809, n_7713);
  not g175501 (n_7808, n_7712);
  nand g175558 (n_7805, n_7081, n_7555);
  nand g175564 (n_7804, n_495, n_7570);
  nand g175573 (n_7803, n_7513, n_7560);
  nand g175585 (n_7802, n_7415, n_7662);
  nand g175587 (n_7801, n_6915, n_7556);
  nand g175597 (n_7800, n_7798, n_7669);
  nand g175598 (n_7799, n_7798, n_7569);
  not g176231 (n_7797, n_7744);
  nand g175816 (n_7796, n_2251, n_7779);
  not g175686 (n_7795, n_7690);
  not g175700 (n_7794, n_7688);
  not g175701 (n_7793, n_7687);
  not g175702 (n_7792, n_7685);
  not g175709 (n_7791, n_7683);
  not g175711 (n_7789, n_7681);
  not g175712 (n_7788, n_7680);
  not g175719 (n_7787, n_7679);
  not g175723 (n_7786, n_7678);
  not g175724 (n_7785, n_7677);
  nand g175814 (n_7783, n_1328, n_7565);
  nand g175735 (n_7782, n_5858, n_7557);
  nand g175740 (n_7781, n_6912, n_7558);
  nand g175806 (n_7780, n_7798, n_7779);
  nand g175811 (n_7778, n_1154, n_7564);
  nand g175812 (n_7777, n_7544, n_7657);
  nand g175625 (n_7962, n_5344, n_7566);
  fflopd g2108_reg(.CK (clock), .D (n_7576), .Q (g2108));
  fflopd g2241_reg(.CK (clock), .D (n_7617), .Q (g2241));
  fflopd g2509_reg(.CK (clock), .D (n_7620), .Q (g2509));
  nand g175630 (n_7957, g150, n_7561);
  nand g176104 (n_7952, g758, n_7670);
  fflopd g4449_reg(.CK (clock), .D (n_7640), .Q (g7260));
  fflopd g1413_reg(.CK (clock), .D (n_7619), .Q (g1413));
  fflopd g1002_reg(.CK (clock), .D (n_7594), .Q (g1002));
  fflopd g1345_reg(.CK (clock), .D (n_7623), .Q (g1345));
  fflopd g2153_reg(.CK (clock), .D (n_7618), .Q (g2153));
  fflopd g2421_reg(.CK (clock), .D (n_7621), .Q (g2421));
  fflopd g744_reg(.CK (clock), .D (n_7599), .Q (g744));
  fflopd g1821_reg(.CK (clock), .D (n_7582), .Q (g1821));
  fflopd g1840_reg(.CK (clock), .D (n_7581), .Q (g1840));
  fflopd g2089_reg(.CK (clock), .D (n_7577), .Q (g2089));
  fflopd g1668_reg(.CK (clock), .D (n_7589), .Q (g1668));
  not g175732 (n_7978, n_7891);
  fflopd g2541_reg(.CK (clock), .D (n_7660), .Q (g2541));
  fflopd g2273_reg(.CK (clock), .D (n_7663), .Q (g2273));
  fflopd g5142_reg(.CK (clock), .D (n_10342), .Q (g5142));
  fflopd g3484_reg(.CK (clock), .D (n_10339), .Q (g3484));
  fflopd g6181_reg(.CK (clock), .D (n_10336), .Q (g6181));
  fflopd g2599_reg(.CK (clock), .D (n_7622), .Q (g2599));
  fflopd g2331_reg(.CK (clock), .D (n_7593), .Q (g2331));
  fflopd g2197_reg(.CK (clock), .D (n_7615), .Q (g2197));
  fflopd g2465_reg(.CK (clock), .D (n_7616), .Q (g2465));
  nand g175402 (n_7776, n_7471, n_7305);
  nand g176494 (n_7775, n_6245, n_7514);
  nand g176507 (n_7774, n_5021, n_8214);
  nand g175133 (n_7773, n_6580, n_7512);
  nand g175147 (n_7772, n_6562, n_7509);
  nand g175148 (n_7771, n_6582, n_7511);
  nand g175161 (n_7770, n_6361, n_7504);
  nand g175162 (n_7769, n_6560, n_7510);
  not g175212 (n_7768, g341);
  nor g175220 (n_7767, n_7282, n_7429);
  nand g175221 (n_7766, g4430, n_7459);
  nand g175229 (n_7765, n_556, n_7461);
  nand g175233 (n_7764, n_572, n_7463);
  nand g175234 (n_7763, n_646, n_7464);
  nand g175248 (n_7762, n_6494, n_7466);
  nor g175250 (n_7761, g294, n_7729);
  nand g175254 (n_7760, n_778, n_7470);
  nand g175255 (n_7759, n_922, n_7472);
  nand g175256 (n_7758, n_1295, n_7473);
  nor g175557 (n_7757, g1982, n_7671);
  nand g175556 (n_7756, n_6903, n_7400);
  not g175347 (n_7755, n_7646);
  not g175361 (n_7752, n_7641);
  not g175367 (n_7751, n_7632);
  nor g175373 (n_7750, n_7427, n_7273);
  nand g175376 (n_7749, n_6428, n_7534);
  nand g175377 (n_7748, n_6430, n_7465);
  nand g175384 (n_7747, n_6379, n_7468);
  nand g175388 (n_7746, g5084, n_7503);
  nand g175389 (n_7745, n_6369, n_7460);
  nand g176458 (n_7744, g758, n_7705);
  nand g175403 (n_7743, n_2510, n_7527);
  nand g175404 (n_7742, n_1751, n_7528);
  nand g175405 (n_7741, n_7462, n_7304);
  nor g175406 (n_7740, n_7274, n_7428);
  nand g175428 (n_7738, g35, n_7476);
  nand g175555 (n_7737, n_6906, n_7396);
  nand g175443 (n_7735, g35, n_7475);
  nand g175445 (n_7734, n_7292, n_7469);
  nand g175446 (n_7733, n_8107, n_7467);
  nand g175447 (n_7732, g1111, n_7601);
  nand g175449 (n_7731, g1124, n_7602);
  nand g175451 (n_7730, g294, n_7729);
  nand g175462 (n_7728, g1682, n_7726);
  nand g175463 (n_7727, g1700, n_7726);
  nand g175464 (n_7725, n_1301, n_7439);
  nand g175466 (n_7724, g676, n_7438);
  nand g175477 (n_7723, g4531, new_g10233_);
  nand g175492 (n_7722, g1094, n_7603);
  nand g175547 (n_7721, n_6943, n_7398);
  nand g175545 (n_7720, n_6932, n_7399);
  nand g175524 (n_7719, g35, n_7397);
  nand g175517 (n_7717, n_6899, n_7417);
  fflopd g5831_reg(.CK (clock), .D (n_7486), .Q (g5831));
  nand g175497 (n_7922, g12919, n_7531);
  fflopd g5471_reg(.CK (clock), .D (n_7482), .Q (g5471));
  fflopd g4608_reg(.CK (clock), .D (n_7516), .Q (g4608));
  fflopd g225_reg(.CK (clock), .D (n_7490), .Q (g225));
  nand g175498 (n_7919, g35, n_7600);
  nand g175738 (n_7716, n_7407, n_7390);
  nand g175576 (n_7715, n_6893, n_7416);
  nand g175577 (n_7714, g35, n_7401);
  nand g175581 (n_7713, n_7410, n_7375);
  nand g175584 (n_7712, n_7412, n_7374);
  nor g175590 (n_7711, g1373, n_7689);
  nor g175591 (n_7710, g1036, n_7707);
  nor g175599 (n_7708, g1030, n_7707);
  nor g175962 (n_7706, g758, n_7705);
  not g175694 (n_7704, n_7590);
  not g175695 (n_7703, n_7588);
  not g175696 (n_7702, n_7585);
  not g175697 (n_7701, n_7584);
  not g175698 (n_7700, n_7580);
  not g175708 (n_7699, n_7578);
  nand g175733 (n_7697, g1886, n_7545);
  nand g175736 (n_7695, n_7403, n_7391);
  nand g175737 (n_7694, g35, n_7404);
  nand g175571 (n_7693, n_720, n_7421);
  nand g175739 (n_7692, n_7411, n_7388);
  nand g175743 (n_7691, g35, n_7536);
  nand g175777 (n_7690, g1373, n_7689);
  nand g175807 (n_7688, g1878, n_7668);
  nand g175808 (n_7687, g1882, n_7568);
  nand g175809 (n_7686, g35, n_7402);
  nand g175810 (n_7685, n_846, n_7424);
  nand g175819 (n_7684, n_6873, n_7541);
  nand g175820 (n_7683, n_1366, n_7532);
  nand g175825 (n_7682, n_1276, n_7538);
  nand g175826 (n_7681, g35, n_7425);
  nand g175831 (n_7680, n_515, n_7423);
  nand g175846 (n_7679, g150, n_7673);
  nand g175852 (n_7678, g1030, n_7707);
  nand g175853 (n_7677, g1036, n_7707);
  nand g175857 (n_7676, n_776, n_7419);
  nor g175569 (n_7674, g150, n_7673);
  nand g176319 (n_7672, n_8904, n_7518);
  not g175909 (n_7882, new_g7558_);
  not g175506 (g34839, n_7609);
  fflopd g5485_reg(.CK (clock), .D (n_7515), .Q (g5485));
  fflopd g5817_reg(.CK (clock), .D (n_7489), .Q (g5817));
  fflopd g3817_reg(.CK (clock), .D (n_7479), .Q (g3817));
  fflopd g2571_reg(.CK (clock), .D (n_7493), .Q (g2571));
  fflopd g2579_reg(.CK (clock), .D (n_7495), .Q (g2579));
  fflopd g2583_reg(.CK (clock), .D (n_7496), .Q (g2583));
  fflopd g6509_reg(.CK (clock), .D (n_7485), .Q (g6509));
  fflopd g6523_reg(.CK (clock), .D (n_7484), .Q (g6523));
  fflopd g3129_reg(.CK (clock), .D (n_7480), .Q (g3129));
  fflopd g2303_reg(.CK (clock), .D (n_7455), .Q (g2303));
  fflopd g2315_reg(.CK (clock), .D (n_7452), .Q (g2315));
  fflopd g4213_reg(.CK (clock), .D (g11770), .Q (g8915));
  nand g175885 (n_7891, g35, n_7671);
  fflopd g2311_reg(.CK (clock), .D (n_7453), .Q (g2311));
  fflopd g3115_reg(.CK (clock), .D (n_7481), .Q (g3115));
  fflopd g3831_reg(.CK (clock), .D (n_7478), .Q (g3831));
  fflopd g1542_reg(.CK (clock), .D (n_7550), .Q (g1542));
  fflopd g2070_reg(.CK (clock), .D (n_7539), .Q (g2070));
  fflopd g1802_reg(.CK (clock), .D (n_7546), .Q (g1802));
  fflopd g446_reg(.CK (clock), .D (n_7483), .Q (g446));
  fflopd g1996_reg(.CK (clock), .D (n_7529), .Q (g1996));
  fflopd g691_reg(.CK (clock), .D (n_7477), .Q (g691));
  not g176537 (n_7670, n_7705);
  not g175900 (n_7669, n_7668);
  nor g175217 (n_7667, n_7108, n_7252);
  nor g175218 (n_7666, n_7111, n_7257);
  nor g175219 (n_7665, n_7112, n_7258);
  nand g175228 (n_7663, n_6829, n_7295);
  nand g175922 (n_7662, g1862, n_7656);
  nor g175251 (n_7661, n_1188, n_7317);
  fflopd g341_reg(.CK (clock), .D (n_7286), .Q (g341));
  nand g175253 (n_7660, n_6848, n_7297);
  not g175704 (n_7659, n_7436);
  not g175699 (n_7658, n_7437);
  nand g175920 (n_7657, g1936, n_7656);
  not g175693 (n_7655, n_7440);
  not g175345 (n_7654, n_7508);
  not g175363 (n_7652, n_7505);
  nand g175371 (n_7651, n_5127, n_7251);
  nor g175374 (n_7650, n_7256, n_7110);
  nand g175411 (n_7649, n_6837, n_7322);
  nand g175412 (n_7648, n_6839, n_7312);
  not g175692 (n_7647, n_7441);
  nand g175452 (n_7646, n_6794, n_7264);
  nand g175456 (n_7645, g3338, n_7320);
  nand g175458 (n_7644, n_499, n_7285);
  nand g175461 (n_7643, g3689, n_7262);
  nand g175468 (n_7642, g25219, n_7321);
  nand g175474 (n_7641, n_972, n_7458);
  nand g175475 (n_7640, n_5599, n_7319);
  nand g175478 (n_7639, g5689, n_7255);
  nand g175480 (n_7638, g6381, n_7318);
  nor g175482 (n_7637, n_7254, n_5564);
  nand g175483 (n_7636, g6035, n_7253);
  nand g175485 (n_7635, n_6159, n_7310);
  nand g175486 (n_7634, g6727, n_7250);
  nand g175491 (n_7633, n_4615, n_7259);
  nand g175493 (n_7632, n_6835, n_7261);
  not g175691 (n_7630, n_7442);
  not g175690 (n_7629, n_7443);
  not g175689 (n_7628, n_7444);
  not g175512 (n_7627, n_7729);
  not g175688 (n_7626, n_7445);
  not g175687 (n_7625, n_7446);
  nand g175520 (n_7624, g35, n_7247);
  nand g175525 (n_7623, n_2658, n_7221);
  nand g175526 (n_7622, n_6345, n_7219);
  nand g175540 (n_7621, n_6506, n_7208);
  nand g175544 (n_7620, n_1396, n_7218);
  nand g175550 (n_7619, n_4822, n_7380);
  nand g175568 (n_7618, n_6507, n_7216);
  nand g175570 (n_7617, n_1269, n_7224);
  nand g175586 (n_7616, n_6343, n_7217);
  nand g175588 (n_7615, n_6340, n_7222);
  nand g175589 (n_7614, n_7535, n_7215);
  nand g175595 (n_7613, n_7611, n_7246);
  nand g175596 (n_7612, n_7611, n_7339);
  nand g175624 (n_7609, g4369, n_7242);
  not g175685 (n_7608, n_7447);
  not g175670 (n_7607, n_7451);
  not g175680 (n_7606, n_7450);
  not g175684 (n_7604, n_7448);
  not g175508 (n_7844, n_7603);
  not g175509 (n_7841, n_7602);
  not g175510 (n_7849, n_7601);
  fflopd g686_reg(.CK (clock), .D (n_7313), .Q (g686));
  not g175515 (n_7851, n_7600);
  fflopd g102_reg(.CK (clock), .D (n_7379), .Q (g20901));
  fflopd g3835_reg(.CK (clock), .D (n_10351), .Q (g3835));
  fflopd g6527_reg(.CK (clock), .D (n_10357), .Q (g6527));
  not g175516 (n_7838, n_7726);
  fflopd g5343_reg(.CK (clock), .D (n_7301), .Q (g25219));
  fflopd g6035_reg(.CK (clock), .D (n_7299), .Q (g6035));
  nand g176318 (n_7599, n_7346, n_7161);
  not g175720 (n_7598, n_7433);
  not g175728 (n_7597, n_7432);
  not g175730 (n_7595, n_7430);
  nand g175742 (n_7594, n_3753, n_7223);
  nand g175749 (n_7593, n_6338, n_7225);
  nand g175776 (n_7592, n_5492, n_7337);
  nand g175782 (n_7591, n_7611, n_7586);
  nand g175789 (n_7590, n_1046, n_7326);
  nand g175790 (n_7589, n_7191, n_7323);
  nand g175791 (n_7588, n_1106, n_7232);
  nand g175792 (n_7587, n_2328, n_7586);
  nand g175794 (n_7585, n_703, n_7227);
  nand g175797 (n_7584, n_1323, n_7373);
  nand g175798 (n_7583, g1802, n_7243);
  nand g175799 (n_7582, n_7188, n_7228);
  nand g175802 (n_7581, n_7186, n_7229);
  nand g175803 (n_7580, n_6947, n_7231);
  nand g175805 (n_7579, n_7798, n_7487);
  nand g175818 (n_7578, n_719, n_7234);
  nand g175827 (n_7577, n_7180, n_7235);
  nand g175829 (n_7576, n_7179, n_7236);
  nand g175830 (n_7575, g2108, n_7367);
  nand g175832 (n_7574, n_2931, n_7289);
  nand g175876 (n_7572, n_7571, n_7244);
  not g175895 (n_7570, n_7408);
  not g175899 (n_7569, n_7568);
  not g175908 (n_7566, n_7689);
  nand g175919 (n_7565, g1950, n_7656);
  nand g175921 (n_7564, g1906, n_7656);
  not g175713 (n_7563, n_7434);
  not g176257 (n_7561, n_7673);
  not g176245 (n_7560, n_7533);
  not g176237 (n_7558, n_7540);
  not g176232 (n_7557, n_7542);
  not g176229 (n_7556, n_7547);
  not g176184 (n_7555, n_7420);
  nor g175963 (n_7552, n_1646, n_7362);
  not g176259 (n_7779, n_7671);
  fflopd g4119_reg(.CK (clock), .D (n_7343), .Q (g4119));
  fflopd g4122_reg(.CK (clock), .D (n_7342), .Q (g4122));
  fflopd g1075_reg(.CK (clock), .D (n_7248), .Q (g17291));
  fflopd g2667_reg(.CK (clock), .D (n_7288), .Q (g2667));
  fflopd g676_reg(.CK (clock), .D (n_7314), .Q (g676));
  fflopd g283_reg(.CK (clock), .D (n_7293), .Q (g283));
  fflopd g2399_reg(.CK (clock), .D (n_7266), .Q (g2399));
  fflopd g336_reg(.CK (clock), .D (n_7393), .Q (g336));
  fflopd g2533_reg(.CK (clock), .D (n_7341), .Q (g2533));
  fflopd g2265_reg(.CK (clock), .D (n_7271), .Q (g2265));
  fflopd g1484_reg(.CK (clock), .D (n_7315), .Q (g1484));
  fflopd g2380_reg(.CK (clock), .D (n_7267), .Q (g2380));
  fflopd g2246_reg(.CK (clock), .D (n_7272), .Q (g2246));
  fflopd g2741_reg(.CK (clock), .D (n_7344), .Q (new_g7558_));
  fflopd g671_reg(.CK (clock), .D (n_7311), .Q (g671));
  fflopd g2514_reg(.CK (clock), .D (n_7340), .Q (g2514));
  fflopd g2648_reg(.CK (clock), .D (n_7389), .Q (g2648));
  fflopd g5835_reg(.CK (clock), .D (n_10360), .Q (g5835));
  fflopd g1183_reg(.CK (clock), .D (n_10146), .Q (g1183));
  fflopd g3133_reg(.CK (clock), .D (n_10354), .Q (g3133));
  fflopd g4709_reg(.CK (clock), .D (n_10148), .Q (g4709));
  fflopd g5489_reg(.CK (clock), .D (n_10363), .Q (g5489));
  fflopd g4601_reg(.CK (clock), .D (n_7241), .Q (g4601));
  fflopd g5046_reg(.CK (clock), .D (n_7363), .Q (g5046));
  fflopd g3338_reg(.CK (clock), .D (n_7303), .Q (g3338));
  fflopd g3689_reg(.CK (clock), .D (n_7306), .Q (g3689));
  fflopd g6727_reg(.CK (clock), .D (n_7302), .Q (g6727));
  fflopd g5689_reg(.CK (clock), .D (n_7300), .Q (g5689));
  fflopd g4040_reg(.CK (clock), .D (n_7307), .Q (g4040));
  fflopd g6381_reg(.CK (clock), .D (n_7308), .Q (g6381));
  nand g176361 (n_7550, n_4575, n_7137);
  nand g176365 (n_7549, g35, n_7395);
  nand g176366 (n_7548, g35, n_7138);
  nand g176446 (n_7547, n_721, n_7134);
  nand g176447 (n_7546, n_7132, n_6897);
  nand g176454 (n_7545, n_2041, n_7543);
  nand g176456 (n_7544, g1906, n_7543);
  nand g176462 (n_7542, n_731, n_7205);
  nand g176464 (n_7541, g4608, n_7136);
  nand g176469 (n_7540, n_1042, n_7145);
  nand g176470 (n_7539, n_7143, n_6895);
  nand g176471 (n_7538, n_4332, n_7422);
  nand g176472 (n_7537, n_7142, n_6944);
  nor g176492 (n_7536, n_7535, n_7394);
  not g175671 (n_7534, n_7291);
  nand g176495 (n_7533, n_773, n_7163);
  nand g176518 (n_7532, n_7046, n_7154);
  nand g175617 (n_7531, n_187, n_7530);
  nand g175615 (n_7529, n_7146, n_7083);
  nor g175610 (n_7528, n_1132, n_7181);
  nor g175608 (n_7527, n_2608, n_7197);
  not g176824 (n_7525, n_7355);
  not g176825 (n_7524, n_7354);
  not g176827 (n_7523, n_7353);
  not g176828 (n_7522, n_7352);
  not g176829 (n_7521, n_7350);
  not g176830 (n_7520, n_7348);
  not g176842 (n_7519, n_7335);
  not g176847 (n_7518, n_7334);
  not g176858 (n_7517, n_7332);
  nand g175583 (n_7516, n_700, n_7043);
  nand g175579 (n_7515, n_6341, n_7052);
  nand g177128 (n_7514, g5046, n_7121);
  nand g177129 (n_7513, g5057, n_7120);
  nand g175372 (n_7512, n_6702, n_7126);
  nand g175375 (n_7511, n_6754, n_7127);
  nand g175407 (n_7510, n_7104, n_6578);
  nand g175408 (n_7509, n_7103, n_6577);
  nand g175448 (n_7508, n_1329, n_7118);
  nand g175455 (n_7507, g3338, n_7105);
  nand g175465 (n_7506, n_7114, n_3999);
  nand g175484 (n_7505, n_791, n_7109);
  nand g175495 (n_7504, n_5790, n_7122);
  not g175507 (n_7503, n_7502);
  nand g175518 (n_7501, g35, n_7069);
  nand g175519 (n_7500, g35, n_7067);
  nand g175521 (n_7499, g35, n_7064);
  nand g175522 (n_7498, g35, n_7051);
  nand g175523 (n_7497, g35, n_7063);
  nand g175527 (n_7496, n_7059, n_7027);
  nand g175528 (n_7495, n_7060, n_7028);
  fflopd g4531_reg(.CK (clock), .D (n_7182), .Q (g4531));
  nand g175532 (n_7494, g35, n_7058);
  nand g175533 (n_7493, n_7057, n_7029);
  nand g175535 (n_7491, g35, n_7053);
  nand g175541 (n_7490, n_2952, n_7054);
  nand g175542 (n_7489, n_6329, n_7055);
  nand g175543 (n_7486, n_6327, n_7056);
  nand g175548 (n_7485, n_6386, n_7061);
  nand g175549 (n_7484, n_6325, n_7062);
  nand g175551 (n_7483, n_3263, n_7068);
  nand g175578 (n_7482, n_6334, n_7078);
  nand g175552 (n_7481, n_6323, n_7065);
  nand g175553 (n_7480, n_6321, n_7066);
  nand g175560 (n_7479, n_6316, n_7070);
  nand g175561 (n_7478, n_6314, n_7071);
  nand g175563 (n_7477, n_538, n_7099);
  nor g175567 (n_7476, g1714, n_7474);
  nor g175575 (n_7475, g5073, n_7082);
  nand g175627 (n_7603, g13259, n_2131);
  not g176255 (g33894, n_7364);
  nand g175650 (n_7600, g13259, n_4291);
  nand g175629 (n_7601, g13259, n_4319);
  nand g175628 (n_7602, g13259, n_4343);
  nand g176526 (n_7673, g164, n_7418);
  fflopd g4049_reg(.CK (clock), .D (n_7150), .Q (g4049));
  nand g176528 (n_7671, n_1317, n_7414);
  nand g175664 (n_7726, g35, n_7474);
  nand g175631 (n_7729, g291, n_7079);
  nand g176768 (n_7705, g749, n_7129);
  fflopd g2629_reg(.CK (clock), .D (n_7195), .Q (g2629));
  fflopd g2287_reg(.CK (clock), .D (n_7123), .Q (g2287));
  not g176884 (n_8214, n_7330);
  fflopd g246_reg(.CK (clock), .D (n_7050), .Q (g246));
  not g175672 (n_7473, n_7290);
  not g175673 (n_7472, n_7298);
  not g175674 (n_7471, n_7329);
  not g175675 (n_7470, n_7345);
  not g175678 (n_7469, n_7356);
  not g175679 (n_7468, n_7384);
  not g175681 (n_7467, n_7385);
  not g175683 (n_7466, n_7249);
  not g175714 (n_7465, n_7278);
  not g175715 (n_7464, n_7277);
  not g175716 (n_7463, n_7276);
  not g175717 (n_7462, n_7275);
  not g175721 (n_7461, n_7270);
  not g175726 (n_7460, n_7268);
  not g175731 (n_7459, n_7458);
  nand g175741 (n_7457, g35, n_7073);
  nand g175745 (n_7455, n_7074, n_7025);
  nand g175746 (n_7454, g35, n_7075);
  nand g175747 (n_7453, n_7076, n_7024);
  nand g175748 (n_7452, n_7077, n_7023);
  nand g175753 (n_7451, n_673, n_7169);
  nand g175766 (n_7450, n_1274, n_7168);
  nand g175768 (n_7449, n_1405, n_7194);
  nand g175773 (n_7448, n_1192, n_7087);
  nand g175775 (n_7447, n_680, n_7049);
  nand g175778 (n_7446, n_636, n_7166);
  nand g175779 (n_7445, n_645, n_7044);
  nand g175780 (n_7444, n_889, n_7080);
  nand g175784 (n_7443, g1608, n_7245);
  nand g175785 (n_7442, g1612, n_7338);
  nand g175786 (n_7441, n_644, n_7090);
  nand g175787 (n_7440, n_729, n_7091);
  nand g175796 (n_7439, g1748, n_7190);
  nand g175801 (n_7438, g35, n_7187);
  nand g175804 (n_7437, n_1235, n_7184);
  nand g175813 (n_7436, n_7203, n_3898);
  nand g175817 (n_7435, n_704, n_7047);
  nand g175835 (n_7434, n_890, n_7167);
  nand g175848 (n_7433, n_641, n_7042);
  nand g175858 (n_7432, n_1175, n_7092);
  nand g175859 (n_7431, n_991, n_7171);
  nand g175863 (n_7430, n_920, n_7089);
  nand g175871 (n_7429, n_7093, n_2082);
  nand g175880 (n_7428, n_7147, n_2080);
  nand g175881 (n_7427, n_7204, n_2104);
  nand g176338 (n_7425, n_2895, n_7160);
  nand g176335 (n_7424, n_7798, n_7158);
  nand g176329 (n_7423, n_132, n_7422);
  nand g176324 (n_7421, n_6949, n_7156);
  nand g176322 (n_7420, n_7135, n_6922);
  nand g176320 (n_7419, n_534, n_7418);
  not g176249 (n_7417, n_7365);
  not g176248 (n_7416, n_7366);
  nand g175945 (n_7415, n_7413, n_7414);
  nand g175947 (n_7412, n_1480, n_7409);
  not g176236 (n_7411, n_7368);
  nand g175953 (n_7410, n_1490, n_7409);
  nand g175954 (n_7408, n_7131, n_6960);
  not g176235 (n_7407, n_7369);
  nand g176337 (g33435, n_6925, n_7149);
  nand g176487 (g33079, n_6924, n_7148);
  not g176234 (n_7404, n_7370);
  not g176233 (n_7403, n_7371);
  not g176230 (n_7402, n_7372);
  not g176225 (n_7401, n_7376);
  not g176222 (n_7400, n_7377);
  not g176199 (n_7399, n_7383);
  not g176202 (n_7398, n_7382);
  not g176210 (n_7397, n_7381);
  not g176221 (n_7396, n_7378);
  nand g175984 (n_7668, g1906, n_7414);
  nand g175980 (n_7568, g1936, n_7395);
  fflopd g723_reg(.CK (clock), .D (n_7119), .Q (g723));
  fflopd g4185_reg(.CK (clock), .D (n_7130), .Q (g11770));
  nand g176112 (n_7689, n_5493, n_7165);
  fflopd g1070_reg(.CK (clock), .D (n_7045), .Q (g1070));
  fflopd g3347_reg(.CK (clock), .D (n_7128), .Q (g3347));
  fflopd g5352_reg(.CK (clock), .D (n_7100), .Q (g5352));
  nand g176154 (n_7707, n_5370, n_7394);
  fflopd g5037_reg(.CK (clock), .D (n_7162), .Q (g5037));
  fflopd g2555_reg(.CK (clock), .D (n_7124), .Q (g2555));
  fflopd g2227_reg(.CK (clock), .D (n_7176), .Q (g2227));
  fflopd g2495_reg(.CK (clock), .D (n_7199), .Q (g2495));
  fflopd g2361_reg(.CK (clock), .D (n_7172), .Q (g2361));
  fflopd g979_reg(.CK (clock), .D (g13259), .Q (g979));
  nand g176359 (n_7393, n_5794, n_6939);
  nand g176360 (n_7392, g35, n_6938);
  nand g176368 (n_7391, g35, n_6937);
  nand g176369 (n_7390, g35, n_6936);
  nand g175769 (n_7389, n_6779, n_6851);
  nand g176370 (n_7388, g35, n_6935);
  nand g176371 (n_7387, g35, n_6965);
  nand g176372 (n_7386, g35, n_6892);
  nand g175767 (n_7385, g291, n_7316);
  nand g175765 (n_7384, n_886, n_6849);
  nand g176400 (n_7383, n_6255, n_6941);
  nand g176403 (n_7382, n_6266, n_6961);
  nand g176418 (n_7381, g1367, n_7336);
  nand g176421 (n_7380, g1413, n_6974);
  nand g176428 (n_7379, n_1148, n_6918);
  nand g176431 (n_7378, n_6263, n_6905);
  nand g176432 (n_7377, n_6260, n_6962);
  nand g176436 (n_7376, g1736, n_7155);
  nand g176438 (n_7375, g1744, n_6902);
  nand g176441 (n_7374, g1752, n_6900);
  nand g176442 (n_7373, g1756, n_6917);
  nand g176455 (n_7372, g1890, n_7157);
  nand g176463 (n_7371, n_687, n_6920);
  nand g176465 (n_7370, g2016, n_7153);
  nand g176466 (n_7369, n_1207, n_6921);
  nand g176468 (n_7368, n_1375, n_6923);
  nand g176476 (n_7367, g35, n_6964);
  nand g176498 (n_7366, n_6264, n_6894);
  nand g176499 (n_7365, n_6259, n_6963);
  nand g176523 (n_7364, g890, n_6958);
  nand g176571 (n_7363, n_5520, n_6874);
  nor g176747 (n_7362, g749, n_7333);
  nand g175764 (n_7356, n_967, n_6815);
  nand g176899 (n_7355, n_7351, n_6877);
  nand g176900 (n_7354, n_7349, n_6865);
  nand g176902 (n_7353, n_7347, n_6863);
  nand g176903 (n_7352, n_7351, n_6862);
  nand g176904 (n_7350, n_7349, n_6861);
  nand g176905 (n_7348, n_7347, n_6859);
  nand g176962 (n_7346, n_8904, n_6868);
  nand g175761 (n_7345, n_6423, n_6846);
  nor g176989 (n_7344, g35, n_8296);
  nand g177007 (n_7343, n_6869, n_5019);
  nand g177009 (n_7342, n_6879, n_5510);
  nand g175760 (n_7341, n_6783, n_6866);
  nand g175759 (n_7340, n_6785, n_6845);
  not g175904 (n_7339, n_7338);
  nor g175929 (n_7337, g1367, n_7336);
  nand g177073 (n_7335, n_7331, n_6864);
  nand g177100 (n_7334, g749, n_7333);
  nand g177123 (n_7332, n_7331, n_6860);
  nand g177158 (n_7330, g35, n_6872);
  nand g175758 (n_7329, n_989, n_7016);
  nand g177382 (n_7328, n_4871, n_6858);
  nand g175928 (n_7327, g1592, n_7325);
  nand g175927 (n_7326, g1636, n_7325);
  not g175505 (n_7324, n_7125);
  nand g175926 (n_7323, g1668, n_7325);
  nor g175529 (n_7322, n_5477, n_6840);
  nand g175530 (n_7321, n_6887, n_3074);
  nand g175536 (n_7320, n_6885, n_3073);
  nand g175537 (n_7319, g4392, n_7206);
  nand g175539 (n_7318, n_6883, n_3072);
  nor g175546 (n_7317, g291, n_7316);
  nand g175554 (n_7315, n_1091, n_6798);
  nand g175559 (n_7314, n_1400, n_6819);
  nand g175562 (n_7313, n_3514, n_6795);
  nor g175574 (n_7312, n_5478, n_6841);
  nand g175582 (n_7311, n_1054, n_6832);
  nand g175594 (n_7310, n_6843, n_1997);
  nand g175602 (n_7309, n_5250, n_6855);
  nand g175604 (n_7308, n_4643, n_6802);
  nand g175605 (n_7307, n_6856, n_4798);
  nand g175606 (n_7306, n_4641, n_6797);
  nand g175607 (n_7305, g2495, n_6808);
  nand g175611 (n_7304, g2227, n_6807);
  nand g175619 (n_7303, n_6854, n_4816);
  nand g175620 (n_7302, n_4639, n_6799);
  nand g175621 (n_7301, n_6853, n_4814);
  nand g175622 (n_7300, n_4642, n_6805);
  nand g175623 (n_7299, n_4640, n_6804);
  nand g175757 (n_7298, n_6462, n_7017);
  not g175676 (n_7297, n_7117);
  not g175722 (n_7295, n_7107);
  nand g175751 (n_7293, n_1094, n_7022);
  nand g175752 (n_7292, n_8107, n_6817);
  nand g175754 (n_7291, n_497, n_6844);
  nand g175755 (n_7290, n_6598, n_7019);
  fflopd g4116_reg(.CK (clock), .D (n_6913), .Q (g4116));
  nand g175626 (n_7502, g5077, n_4656);
  fflopd g5698_reg(.CK (clock), .D (n_6806), .Q (g5698));
  fflopd g6736_reg(.CK (clock), .D (n_6800), .Q (g6736));
  fflopd g3288_reg(.CK (clock), .D (n_10156), .Q (new_g10366_));
  not g176883 (n_7656, n_7543);
  fflopd g1199_reg(.CK (clock), .D (n_6916), .Q (g1199));
  fflopd g3990_reg(.CK (clock), .D (n_10160), .Q (new_g10375_));
  fflopd g5644_reg(.CK (clock), .D (n_10150), .Q (new_g10401_));
  nand g176339 (n_7289, n_4542, n_7159);
  nand g175771 (n_7288, n_6776, n_6852);
  nand g175772 (n_7287, g2667, n_7009);
  nand g175774 (n_7286, n_7006, n_493);
  nand g175781 (n_7285, n_7611, n_7151);
  nand g175783 (n_7284, g3689, n_6980);
  nand g175793 (n_7283, g4040, n_6979);
  nand g175821 (n_7282, n_1914, n_6811);
  nand g175828 (n_7281, g5689, n_6977);
  nand g175833 (n_7280, g6381, n_6976);
  nand g175834 (n_7279, g6035, n_6975);
  nand g175837 (n_7278, n_879, n_6812);
  nand g175838 (n_7277, n_6502, n_6989);
  nand g175840 (n_7276, n_6478, n_6988);
  nand g175841 (n_7275, n_1247, n_6987);
  nand g175843 (n_7274, n_1931, n_6813);
  nand g175845 (n_7273, n_1943, n_6823);
  nand g175847 (n_7272, n_6762, n_6824);
  nand g175849 (n_7271, n_6761, n_6825);
  nand g175850 (n_7270, n_6425, n_6827);
  nand g175855 (n_7269, g5077, n_7026);
  nand g175856 (n_7268, n_1229, n_6830);
  nand g175860 (n_7267, n_6758, n_6831);
  nand g175861 (n_7266, n_6757, n_6833);
  nand g175862 (n_7265, g2399, n_6982);
  nand g175864 (n_7264, n_7263, n_6870);
  nand g175867 (n_7262, n_6880, n_2090);
  nand g175869 (n_7261, n_7260, n_6878);
  nor g175870 (n_7259, n_5465, n_6978);
  nand g175872 (n_7258, n_6889, n_2076);
  nand g175873 (n_7257, n_7038, n_2074);
  nand g175874 (n_7256, n_6882, n_2108);
  nand g175875 (n_7255, n_7037, n_2077);
  nand g175877 (n_7254, n_5787, n_6838);
  nand g175878 (n_7253, n_7036, n_2085);
  nand g175879 (n_7252, n_7034, n_2087);
  nor g175882 (n_7251, n_5463, n_6994);
  nand g175883 (n_7250, n_7032, n_2078);
  nand g175770 (n_7249, n_4180, n_7030);
  not g175886 (n_7248, n_7164);
  not g175891 (n_7247, n_7041);
  not g175903 (n_7246, n_7245);
  nor g176328 (n_7244, g2108, n_7098);
  nor g176325 (n_7243, g1772, n_7095);
  nand g176292 (n_7242, n_6966, n_2723);
  nand g175933 (n_7241, n_1257, n_6927);
  nand g176277 (n_7239, g2116, n_7237);
  nand g176276 (n_7238, g2112, n_7237);
  nand g176275 (n_7236, g2108, n_7237);
  nand g176274 (n_7235, g2089, n_7237);
  nand g176269 (n_7234, g2008, n_7237);
  nand g176268 (n_7233, g1848, n_7230);
  nand g175941 (n_7232, g1682, n_7325);
  nand g176267 (n_7231, g1844, n_7230);
  nand g176266 (n_7229, g1840, n_7230);
  nand g176265 (n_7228, g1821, n_7230);
  nand g176264 (n_7227, g1740, n_7230);
  not g176252 (n_7225, n_7173);
  not g176243 (n_7224, n_7174);
  not g176242 (n_7223, n_7175);
  not g176241 (n_7222, n_7177);
  not g176209 (n_7221, n_7192);
  not g176203 (n_7219, n_7196);
  not g176194 (n_7218, n_7198);
  not g176189 (n_7217, n_7200);
  not g176185 (n_7216, n_7085);
  nor g175959 (n_7215, n_6752, n_7096);
  not g176183 (n_7208, n_7084);
  nor g175986 (n_7487, g1906, n_7097);
  nand g175884 (n_7458, n_3986, n_7206);
  not g176258 (n_7586, n_7474);
  fflopd g542_reg(.CK (clock), .D (n_6875), .Q (g542));
  fflopd g5134_reg(.CK (clock), .D (n_6896), .Q (g5134));
  fflopd g3698_reg(.CK (clock), .D (n_6796), .Q (g3698));
  fflopd g6390_reg(.CK (clock), .D (n_6801), .Q (g6390));
  fflopd g6044_reg(.CK (clock), .D (n_6803), .Q (g6044));
  fflopd g2941_reg(.CK (clock), .D (n_6954), .Q (g2941));
  fflopd g3125_reg(.CK (clock), .D (n_6908), .Q (g3125));
  fflopd g5827_reg(.CK (clock), .D (n_6930), .Q (g5827));
  fflopd g6173_reg(.CK (clock), .D (n_6942), .Q (g6173));
  fflopd g5481_reg(.CK (clock), .D (n_6911), .Q (g5481));
  fflopd g3476_reg(.CK (clock), .D (n_6904), .Q (g3476));
  fflopd g6519_reg(.CK (clock), .D (n_6973), .Q (g6519));
  fflopd g3827_reg(.CK (clock), .D (n_6898), .Q (g3827));
  fflopd g490_reg(.CK (clock), .D (n_10366), .Q (g490));
  fflopd g1536_reg(.CK (clock), .D (n_6907), .Q (g1536));
  fflopd g1193_reg(.CK (clock), .D (n_6931), .Q (g1193));
  fflopd g3639_reg(.CK (clock), .D (n_10158), .Q (new_g10371_));
  fflopd g1418_reg(.CK (clock), .D (n_6940), .Q (g17320));
  fflopd g6682_reg(.CK (clock), .D (n_10162), .Q (new_g10413_));
  fflopd g5990_reg(.CK (clock), .D (n_10152), .Q (new_g10405_));
  fflopd g6336_reg(.CK (clock), .D (n_10154), .Q (new_g10409_));
  fflopd g4785_reg(.CK (clock), .D (n_6871), .Q (g4785));
  fflopd g5297_reg(.CK (clock), .D (n_10164), .Q (g5297));
  fflopd g5033_reg(.CK (clock), .D (n_10432), .Q (g5033));
  nand g176930 (n_7205, n_5340, n_6488);
  nand g176352 (n_7204, n_6749, n_5789);
  nand g176355 (n_7203, g4366, n_9257);
  nand g176362 (n_7202, g35, n_7039);
  nand g176363 (n_7201, g35, n_6537);
  nand g176386 (n_7200, n_1384, n_6534);
  nand g176389 (n_7199, n_6532, n_6330);
  nand g176392 (n_7198, n_6531, n_6384);
  nand g176404 (n_7197, n_244, n_6553);
  nand g176405 (n_7196, n_1160, n_6548);
  nand g176406 (n_7195, n_6546, n_6324);
  nand g176407 (n_7194, n_4328, n_7086);
  nand g176408 (n_7193, n_6545, n_6421);
  nand g176416 (n_7192, n_1195, n_6539);
  nand g176433 (n_7191, g1636, n_6909);
  nand g176439 (n_7190, n_1780, n_6517);
  nand g176440 (n_7189, g1802, n_6747);
  nand g176448 (n_7188, g1816, n_7185);
  nand g176449 (n_7187, g703, n_6515);
  nand g176450 (n_7186, g1834, n_7185);
  nand g176451 (n_7184, g35, n_6748);
  nand g176457 (n_7183, g35, n_6550);
  nand g176460 (n_7182, n_6536, n_4049);
  nand g176461 (n_7181, n_1399, n_6551);
  nand g176473 (n_7180, g2084, n_7178);
  nand g176475 (n_7179, g2102, n_7178);
  nand g176485 (n_7177, n_872, n_6529);
  nand g176486 (n_7176, n_6527, n_6417);
  nand g176488 (n_7175, n_711, n_6538);
  nand g176489 (n_7174, n_6526, n_6382);
  nand g176502 (n_7173, n_1137, n_6543);
  nand g176503 (n_7172, n_6541, n_6319);
  nand g176504 (n_7171, n_4761, n_7088);
  nand g176505 (n_7170, n_6540, n_6726);
  nand g176511 (n_7169, n_6427, n_6575);
  nand g176512 (n_7168, n_6512, n_6565);
  nand g176522 (n_7167, n_6429, n_6569);
  nand g175935 (n_7166, n_6350, n_6521);
  not g176545 (n_7165, n_7336);
  nand g175931 (n_7164, n_1050, n_6731);
  nand g176556 (n_7163, n_601, n_6479);
  nand g176608 (n_7162, n_3958, n_6477);
  nor g176746 (n_7161, n_1675, n_6492);
  not g176865 (n_7160, n_7159);
  not g176866 (n_7158, n_7157);
  not g176869 (n_7156, n_7155);
  not g176872 (n_7154, n_7153);
  not g175897 (n_7150, n_6821);
  nor g176892 (n_7149, n_6484, n_6471);
  nor g176895 (n_7148, n_6486, n_6469);
  nand g176351 (n_7147, n_6750, n_6884);
  nand g176948 (n_7146, g1996, n_7144);
  nand g176949 (n_7145, g2040, n_7144);
  nand g176950 (n_7143, g2070, n_7144);
  nand g176951 (n_7142, g2084, n_7144);
  nor g176980 (n_7138, n_4654, n_7094);
  nand g177001 (n_7137, g35, n_6500);
  nand g177011 (n_7136, g35, n_6483);
  nand g177022 (n_7135, g1728, n_7133);
  nand g177023 (n_7134, g1772, n_7133);
  nand g177024 (n_7132, g1802, n_7133);
  nand g177025 (n_7131, g1816, n_7133);
  nand g177095 (n_7130, n_1340, n_6475);
  not g177206 (n_7129, n_7333);
  not g175898 (n_7128, n_6820);
  nor g175609 (n_7127, n_6465, n_2610);
  nor g175612 (n_7126, n_6498, n_2613);
  nand g175613 (n_7125, n_6459, n_2089);
  nand g175614 (n_7124, n_6549, n_6518);
  nand g175616 (n_7123, n_6544, n_6559);
  nor g175618 (n_7122, n_6496, n_2622);
  nand g177901 (n_7121, g35, n_6466);
  nand g177903 (n_7120, n_4587, n_6857);
  nand g175750 (n_7119, n_3690, n_6767);
  nand g175756 (n_7118, g2441, n_6789);
  nand g175762 (n_7117, n_1234, n_6781);
  nand g175763 (n_7116, n_682, n_6513);
  nand g175788 (n_7115, n_6583, n_4737);
  nand g175795 (n_7114, g4040, n_6619);
  nand g175800 (n_7113, new_g10354_, n_6453);
  nand g175822 (n_7112, n_1938, n_6451);
  nand g175823 (n_7111, n_1937, n_6455);
  nand g175824 (n_7110, n_1936, n_6457);
  nand g175839 (n_7109, g2173, n_6764);
  nand g175842 (n_7108, n_1932, n_6458);
  nand g175851 (n_7107, n_1388, n_6759);
  nand g175854 (n_7106, n_1109, n_6464);
  nand g175865 (n_7105, n_6755, n_6156);
  nor g175866 (n_7104, n_6163, n_6461);
  nor g175868 (n_7103, n_6162, n_6497);
  not g175896 (n_7100, n_6822);
  not g175894 (n_7099, n_6828);
  fflopd g2856_reg(.CK (clock), .D (n_6649), .Q (g2856));
  not g176877 (n_7422, n_7098);
  not g176881 (n_7395, n_7097);
  not g176546 (n_7394, n_7096);
  not g176542 (n_7409, n_7095);
  fflopd g3949_reg(.CK (clock), .D (n_6596), .Q (g3949));
  fflopd g5228_reg(.CK (clock), .D (n_6719), .Q (g5228));
  fflopd g5244_reg(.CK (clock), .D (n_6723), .Q (g5244));
  fflopd g5236_reg(.CK (clock), .D (n_6721), .Q (g5236));
  fflopd g3255_reg(.CK (clock), .D (n_6630), .Q (g3255));
  fflopd g5551_reg(.CK (clock), .D (n_6585), .Q (g5551));
  fflopd g3598_reg(.CK (clock), .D (n_6616), .Q (g3598));
  fflopd g3897_reg(.CK (clock), .D (n_6609), .Q (g3897));
  fflopd g3917_reg(.CK (clock), .D (n_6605), .Q (g3917));
  fflopd g5268_reg(.CK (clock), .D (n_6730), .Q (g5268));
  nor g177151 (n_7418, n_5276, n_6467);
  nor g177153 (n_7414, g1936, n_7094);
  nand g177157 (n_7543, g35, n_7094);
  fflopd g6295_reg(.CK (clock), .D (n_6663), .Q (g6295));
  fflopd g5200_reg(.CK (clock), .D (n_6713), .Q (g5200));
  fflopd g3546_reg(.CK (clock), .D (n_6626), .Q (g3546));
  fflopd g3582_reg(.CK (clock), .D (n_6771), .Q (g3582));
  fflopd g3566_reg(.CK (clock), .D (n_6622), .Q (g3566));
  fflopd g3219_reg(.CK (clock), .D (n_6639), .Q (g3219));
  fflopd g5889_reg(.CK (clock), .D (n_6695), .Q (g5889));
  fflopd g6593_reg(.CK (clock), .D (n_6656), .Q (g6593));
  fflopd g6291_reg(.CK (clock), .D (n_6664), .Q (g6291));
  fflopd g5615_reg(.CK (clock), .D (n_6699), .Q (g5615));
  fflopd g5607_reg(.CK (clock), .D (n_6701), .Q (g5607));
  fflopd g6621_reg(.CK (clock), .D (n_6732), .Q (g6621));
  fflopd g5583_reg(.CK (clock), .D (n_6706), .Q (g5583));
  fflopd g5575_reg(.CK (clock), .D (n_6707), .Q (g5575));
  fflopd g5591_reg(.CK (clock), .D (n_6705), .Q (g5591));
  fflopd g6609_reg(.CK (clock), .D (n_6654), .Q (g6609));
  fflopd g6299_reg(.CK (clock), .D (n_6696), .Q (g6299));
  fflopd g3933_reg(.CK (clock), .D (n_6601), .Q (g3933));
  fflopd g3251_reg(.CK (clock), .D (n_6631), .Q (g3251));
  fflopd g4191_reg(.CK (clock), .D (n_6766), .Q (g11447));
  fflopd g5220_reg(.CK (clock), .D (n_6717), .Q (g5220));
  fflopd g5252_reg(.CK (clock), .D (n_6725), .Q (g5252));
  fflopd g6605_reg(.CK (clock), .D (n_6698), .Q (g6605));
  fflopd g6613_reg(.CK (clock), .D (n_6653), .Q (g6613));
  fflopd g6617_reg(.CK (clock), .D (n_6660), .Q (g6617));
  fflopd g6625_reg(.CK (clock), .D (n_6586), .Q (g6625));
  fflopd g6629_reg(.CK (clock), .D (n_6612), .Q (g6629));
  fflopd g6633_reg(.CK (clock), .D (n_6652), .Q (g6633));
  fflopd g6641_reg(.CK (clock), .D (n_6591), .Q (g6641));
  fflopd g6649_reg(.CK (clock), .D (n_6588), .Q (g6649));
  fflopd g3191_reg(.CK (clock), .D (n_6645), .Q (g3191));
  fflopd g3199_reg(.CK (clock), .D (n_6643), .Q (g3199));
  nand g176527 (n_7474, n_582, n_7040);
  fflopd g6287_reg(.CK (clock), .D (n_6665), .Q (g6287));
  fflopd g3215_reg(.CK (clock), .D (n_6640), .Q (g3215));
  fflopd g3223_reg(.CK (clock), .D (n_6638), .Q (g3223));
  fflopd g3227_reg(.CK (clock), .D (n_6637), .Q (g3227));
  fflopd g3231_reg(.CK (clock), .D (n_6636), .Q (g3231));
  fflopd g3239_reg(.CK (clock), .D (n_6634), .Q (g3239));
  fflopd g3243_reg(.CK (clock), .D (n_6633), .Q (g3243));
  fflopd g3247_reg(.CK (clock), .D (n_6632), .Q (g3247));
  fflopd g3259_reg(.CK (clock), .D (n_6629), .Q (g3259));
  fflopd g6741_reg(.CK (clock), .D (n_6737), .Q (new_g7097_));
  fflopd g4054_reg(.CK (clock), .D (n_6739), .Q (new_g6928_));
  nand g176345 (n_7093, n_6751, n_6886);
  nand g176336 (n_7092, n_6463, n_6567);
  nand g176334 (n_7091, n_7611, n_6573);
  nand g176333 (n_7090, n_7611, n_6571);
  nand g176331 (n_7089, n_111, n_7088);
  nand g176327 (n_7087, n_213, n_7086);
  nand g176323 (n_7085, n_6530, n_6354);
  nand g176321 (n_7084, n_6535, n_6355);
  nand g176310 (n_7083, n_982, n_6734);
  not g175907 (n_7082, g5077);
  nand g176304 (n_7081, n_488, n_6552);
  nand g176263 (n_7080, n_6352, n_6519);
  not g176256 (n_7079, n_7316);
  not g176254 (n_7078, n_6981);
  not g176251 (n_7077, n_6983);
  not g176250 (n_7076, n_6984);
  not g176247 (n_7075, n_6985);
  not g176246 (n_7074, n_6986);
  not g176240 (n_7073, n_6991);
  not g176239 (n_7072, n_6992);
  not g176227 (n_7071, n_6996);
  not g176226 (n_7070, n_6997);
  not g176220 (n_7069, n_6999);
  not g176218 (n_7068, n_7001);
  not g176219 (n_7067, n_7000);
  not g176217 (n_7066, n_7002);
  not g176215 (n_7065, n_7003);
  not g176214 (n_7064, n_7004);
  not g176213 (n_7063, n_7005);
  not g176208 (n_7062, n_7007);
  not g176207 (n_7061, n_7008);
  not g176200 (n_7060, n_7011);
  not g176201 (n_7059, n_7010);
  not g176198 (n_7058, n_7012);
  not g176197 (n_7057, n_7013);
  not g176193 (n_7056, n_7014);
  not g176192 (n_7055, n_7015);
  not g176188 (n_7054, n_7018);
  not g176187 (n_7053, n_7020);
  not g176186 (n_7052, n_7021);
  not g176179 (n_7051, n_6810);
  nand g175976 (n_7050, n_3334, n_6576);
  nand g175942 (n_7049, n_7901, n_6746);
  nor g175969 (n_7048, n_4079, n_6648);
  nand g175925 (n_7047, n_7046, n_6933);
  nand g175960 (n_7045, n_4870, n_6525);
  nand g175958 (n_7044, n_6441, n_6520);
  nand g175950 (n_7043, n_6926, n_6558);
  nand g175943 (n_7042, n_6890, n_6753);
  nand g175946 (n_7041, n_1428, n_7040);
  nor g175987 (n_7530, g19334, g990);
  nand g175989 (n_7245, g1636, n_7040);
  nand g175990 (n_7338, g1668, n_7039);
  fflopd g5957_reg(.CK (clock), .D (n_6679), .Q (g5957));
  fflopd g5953_reg(.CK (clock), .D (n_6680), .Q (g5953));
  fflopd g5949_reg(.CK (clock), .D (n_6681), .Q (g5949));
  fflopd g5945_reg(.CK (clock), .D (n_6682), .Q (g5945));
  fflopd g5941_reg(.CK (clock), .D (n_6683), .Q (g5941));
  fflopd g5933_reg(.CK (clock), .D (n_6685), .Q (g5933));
  fflopd g5929_reg(.CK (clock), .D (n_6686), .Q (g5929));
  fflopd g5925_reg(.CK (clock), .D (n_6687), .Q (g5925));
  fflopd g5917_reg(.CK (clock), .D (n_6689), .Q (g5917));
  fflopd g5913_reg(.CK (clock), .D (n_6690), .Q (g5913));
  fflopd g5909_reg(.CK (clock), .D (n_6691), .Q (g5909));
  fflopd g5893_reg(.CK (clock), .D (n_6694), .Q (g5893));
  fflopd g5897_reg(.CK (clock), .D (n_6693), .Q (g5897));
  fflopd g5543_reg(.CK (clock), .D (n_6711), .Q (g5543));
  fflopd g5611_reg(.CK (clock), .D (n_6700), .Q (g5611));
  fflopd g5603_reg(.CK (clock), .D (n_6790), .Q (g5603));
  fflopd g5599_reg(.CK (clock), .D (n_6703), .Q (g5599));
  fflopd g5595_reg(.CK (clock), .D (n_6704), .Q (g5595));
  fflopd g6239_reg(.CK (clock), .D (n_6676), .Q (g6239));
  fflopd g5587_reg(.CK (clock), .D (n_6589), .Q (g5587));
  fflopd g5579_reg(.CK (clock), .D (n_6697), .Q (g5579));
  fflopd g5571_reg(.CK (clock), .D (n_6587), .Q (g5571));
  fflopd g5567_reg(.CK (clock), .D (n_6592), .Q (g5567));
  fflopd g6589_reg(.CK (clock), .D (n_6657), .Q (g6589));
  fflopd g6601_reg(.CK (clock), .D (n_6655), .Q (g6601));
  fflopd g739_reg(.CK (clock), .D (n_6514), .Q (g739));
  fflopd g3542_reg(.CK (clock), .D (n_6627), .Q (g3542));
  fflopd g3538_reg(.CK (clock), .D (n_6628), .Q (g3538));
  fflopd g3550_reg(.CK (clock), .D (n_6625), .Q (g3550));
  fflopd g3558_reg(.CK (clock), .D (n_6624), .Q (g3558));
  fflopd g3562_reg(.CK (clock), .D (n_6623), .Q (g3562));
  fflopd g3570_reg(.CK (clock), .D (n_6621), .Q (g3570));
  fflopd g6645_reg(.CK (clock), .D (n_6651), .Q (g6645));
  fflopd g6247_reg(.CK (clock), .D (n_6674), .Q (g6247));
  fflopd g650_reg(.CK (clock), .D (n_6493), .Q (g650));
  fflopd g3574_reg(.CK (clock), .D (n_6620), .Q (g3574));
  fflopd g5041_reg(.CK (clock), .D (n_6489), .Q (g5041));
  fflopd g3578_reg(.CK (clock), .D (n_6765), .Q (g3578));
  fflopd g3586_reg(.CK (clock), .D (n_6584), .Q (g3586));
  fflopd g3235_reg(.CK (clock), .D (n_6635), .Q (g3235));
  fflopd g6259_reg(.CK (clock), .D (n_6672), .Q (g6259));
  fflopd g6263_reg(.CK (clock), .D (n_6671), .Q (g6263));
  fflopd g6267_reg(.CK (clock), .D (n_6670), .Q (g6267));
  fflopd g5921_reg(.CK (clock), .D (n_6688), .Q (g5921));
  fflopd g6275_reg(.CK (clock), .D (n_6668), .Q (g6275));
  fflopd g6279_reg(.CK (clock), .D (n_6667), .Q (g6279));
  fflopd g6581_reg(.CK (clock), .D (n_6659), .Q (g6581));
  fflopd g5901_reg(.CK (clock), .D (n_6692), .Q (g5901));
  fflopd g5961_reg(.CK (clock), .D (n_6678), .Q (g5961));
  fflopd g6585_reg(.CK (clock), .D (n_6658), .Q (g6585));
  fflopd g3211_reg(.CK (clock), .D (n_6641), .Q (g3211));
  fflopd g6271_reg(.CK (clock), .D (n_6669), .Q (g6271));
  fflopd g5937_reg(.CK (clock), .D (n_6684), .Q (g5937));
  fflopd g3195_reg(.CK (clock), .D (n_6644), .Q (g3195));
  fflopd g3207_reg(.CK (clock), .D (n_6642), .Q (g3207));
  fflopd g5555_reg(.CK (clock), .D (n_6709), .Q (g5555));
  fflopd g5563_reg(.CK (clock), .D (n_6708), .Q (g5563));
  fflopd g5547_reg(.CK (clock), .D (n_6710), .Q (g5547));
  fflopd g6255_reg(.CK (clock), .D (n_6673), .Q (g6255));
  fflopd g6235_reg(.CK (clock), .D (n_6677), .Q (g6235));
  fflopd g3590_reg(.CK (clock), .D (n_6618), .Q (g3590));
  fflopd g6243_reg(.CK (clock), .D (n_6675), .Q (g6243));
  fflopd g5264_reg(.CK (clock), .D (n_6729), .Q (g5264));
  fflopd g5260_reg(.CK (clock), .D (n_6728), .Q (g5260));
  fflopd g5256_reg(.CK (clock), .D (n_6727), .Q (g5256));
  fflopd g3187_reg(.CK (clock), .D (n_6646), .Q (g3187));
  fflopd g5248_reg(.CK (clock), .D (n_6724), .Q (g5248));
  fflopd g5240_reg(.CK (clock), .D (n_6722), .Q (g5240));
  fflopd g5232_reg(.CK (clock), .D (n_6720), .Q (g5232));
  fflopd g5224_reg(.CK (clock), .D (n_6718), .Q (g5224));
  fflopd g5216_reg(.CK (clock), .D (n_6716), .Q (g5216));
  fflopd g5208_reg(.CK (clock), .D (n_6715), .Q (g5208));
  fflopd g5204_reg(.CK (clock), .D (n_6714), .Q (g5204));
  fflopd g5196_reg(.CK (clock), .D (n_6712), .Q (g5196));
  fflopd g6283_reg(.CK (clock), .D (n_6666), .Q (g6283));
  fflopd g6303_reg(.CK (clock), .D (n_6662), .Q (g6303));
  fflopd g6307_reg(.CK (clock), .D (n_6661), .Q (g6307));
  fflopd g3961_reg(.CK (clock), .D (n_6593), .Q (g3961));
  fflopd g3957_reg(.CK (clock), .D (n_6594), .Q (g3957));
  fflopd g3953_reg(.CK (clock), .D (n_6595), .Q (g3953));
  fflopd g3945_reg(.CK (clock), .D (n_6597), .Q (g3945));
  fflopd g3941_reg(.CK (clock), .D (n_6599), .Q (g3941));
  fflopd g3937_reg(.CK (clock), .D (n_6600), .Q (g3937));
  fflopd g3929_reg(.CK (clock), .D (n_6602), .Q (g3929));
  fflopd g3925_reg(.CK (clock), .D (n_6603), .Q (g3925));
  fflopd g3921_reg(.CK (clock), .D (n_6604), .Q (g3921));
  fflopd g3913_reg(.CK (clock), .D (n_6606), .Q (g3913));
  fflopd g3909_reg(.CK (clock), .D (n_6607), .Q (g3909));
  fflopd g3901_reg(.CK (clock), .D (n_6608), .Q (g3901));
  fflopd g3893_reg(.CK (clock), .D (n_6610), .Q (g3893));
  fflopd g3889_reg(.CK (clock), .D (n_6611), .Q (g3889));
  fflopd g3610_reg(.CK (clock), .D (n_6613), .Q (g3610));
  fflopd g6637_reg(.CK (clock), .D (n_6590), .Q (g6637));
  fflopd g3606_reg(.CK (clock), .D (n_6614), .Q (g3606));
  fflopd g6653_reg(.CK (clock), .D (n_6650), .Q (g6653));
  fflopd g3602_reg(.CK (clock), .D (n_6615), .Q (g3602));
  fflopd g3594_reg(.CK (clock), .D (n_6617), .Q (g3594));
  fflopd g4801_reg(.CK (clock), .D (n_6482), .Q (g4801));
  fflopd g324_reg(.CK (clock), .D (n_10453), .Q (g324));
  fflopd g3703_reg(.CK (clock), .D (n_6555), .Q (new_g6905_));
  fflopd g5703_reg(.CK (clock), .D (n_6735), .Q (new_g7028_));
  fflopd g6049_reg(.CK (clock), .D (n_6736), .Q (new_g7051_));
  fflopd g3352_reg(.CK (clock), .D (n_6738), .Q (new_g6875_));
  fflopd g4899_reg(.CK (clock), .D (n_6490), .Q (g4899));
  fflopd g6395_reg(.CK (clock), .D (n_6556), .Q (new_g7074_));
  fflopd g1171_reg(.CK (clock), .D (n_6740), .Q (g1171));
  fflopd g5357_reg(.CK (clock), .D (n_6554), .Q (new_g7004_));
  fflopd g1116_reg(.CK (clock), .D (g19334), .Q (g13259));
  nand g176347 (n_7038, n_6439, n_7035);
  nand g176348 (n_7037, n_6888, n_6404);
  nand g176349 (n_7036, n_7035, n_6400);
  nand g176350 (n_7034, n_6366, n_7031);
  nand g176353 (n_7032, n_7031, n_6398);
  nand g176354 (n_7030, g316, n_9257);
  nand g176356 (n_7029, g35, n_6412);
  nand g176357 (n_7028, g35, n_6411);
  nand g176358 (n_7027, g35, n_6408);
  nand g176373 (n_7026, g35, n_6381);
  nand g176374 (n_7025, g35, n_6396);
  nand g176375 (n_7024, g35, n_6406);
  nand g176376 (n_7023, g35, n_6407);
  nand g176377 (n_7022, n_39, n_8107);
  nand g176378 (n_7021, n_6243, n_6431);
  nand g176379 (n_7020, g2429, n_6574);
  nand g176380 (n_7019, g2437, n_6333);
  nand g176382 (n_7018, n_6346, n_3269);
  nand g176384 (n_7017, g2445, n_6331);
  nand g176385 (n_7016, g2449, n_6336);
  nand g176390 (n_7015, n_6240, n_6328);
  nand g176391 (n_7014, n_6236, n_6432);
  nand g176398 (n_7013, n_1206, n_6383);
  nand g176399 (n_7012, g2575, n_6564);
  nand g176401 (n_7011, n_506, n_6349);
  nand g176402 (n_7010, n_522, n_6344);
  nand g176413 (n_7009, g35, n_6436);
  nand g176414 (n_7008, n_6228, n_6326);
  nand g176415 (n_7007, n_6224, n_6433);
  nand g176417 (n_7006, g35, g316);
  nand g176422 (n_7005, g1437, n_6351);
  nand g176423 (n_7004, g1467, n_6353);
  nand g176424 (n_7003, n_6223, n_6322);
  nand g176426 (n_7002, n_6220, n_6434);
  nand g176427 (n_7001, n_551, n_6337);
  nand g176429 (n_7000, g1616, n_6570);
  nand g176430 (n_6999, g1620, n_6572);
  nand g176437 (n_6998, n_6317, n_6362);
  nand g176443 (n_6997, n_6235, n_6315);
  nand g176444 (n_6996, n_6232, n_6435);
  nand g176459 (n_6995, g35, n_6388);
  nand g176467 (n_6994, n_4618, n_6371);
  nand g176474 (n_6993, n_6391, n_6360);
  nand g176477 (n_6992, n_6367, n_5786);
  nand g176478 (n_6991, g2161, n_6568);
  nand g176479 (n_6990, n_6413, n_6358);
  nand g176480 (n_6989, g2169, n_6414);
  nand g176483 (n_6988, g2177, n_6416);
  nand g176484 (n_6987, g2181, n_6335);
  nand g176496 (n_6986, n_573, n_6370);
  nand g176497 (n_6985, g2307, n_6566);
  nand g176500 (n_6984, n_692, n_6375);
  nand g176501 (n_6983, n_1180, n_6380);
  nand g176509 (n_6982, g35, n_6385);
  nand g176510 (n_6981, n_6230, n_6390);
  nand g176514 (n_6980, n_6377, n_5761);
  nand g176516 (n_6979, n_6376, n_5759);
  nand g176517 (n_6978, n_6365, n_5132);
  nand g176519 (n_6977, n_6374, n_5757);
  nand g176520 (n_6976, n_6373, n_5756);
  nand g176521 (n_6975, n_6372, n_5755);
  nand g177056 (n_6974, n_5317, n_6499);
  nand g177051 (n_6973, n_5911, n_6227);
  not g176535 (n_6966, g4366);
  not g176548 (n_6965, g19334);
  nand g176550 (n_6964, g2102, n_6928);
  nand g176555 (n_6963, n_2736, n_6270);
  nand g176559 (n_6962, n_2816, n_6275);
  nand g176564 (n_6961, n_2741, n_6272);
  nand g176575 (n_6960, n_4746, n_6910);
  nand g176599 (n_6958, g479, n_2537);
  nand g176679 (n_6954, n_1692, n_6281);
  nand g176721 (n_6950, n_6949, n_6946);
  nand g176742 (n_6947, n_2243, n_6946);
  nand g176755 (n_6944, n_5491, n_6791);
  nand g177049 (n_6943, g6173, n_6194);
  nand g177048 (n_6942, n_5895, n_6267);
  nand g177047 (n_6941, g6159, n_6273);
  not g176826 (n_6940, n_6557);
  not g176838 (n_6939, n_6524);
  not g176839 (n_6938, n_6523);
  not g176849 (n_6937, n_6511);
  not g176850 (n_6936, n_6510);
  not g176851 (n_6935, n_6509);
  nand g177045 (n_6932, g6154, n_6292);
  nand g177042 (n_6931, n_1220, n_6195);
  nand g177040 (n_6930, n_6074, n_6239);
  nand g176913 (n_6929, n_7046, n_6928);
  nand g176914 (n_6927, n_6926, n_5910);
  nor g176922 (n_6925, n_6247, n_6246);
  nor g176926 (n_6924, n_6251, n_6249);
  nand g176963 (n_6923, n_7046, n_6305);
  nand g176968 (n_6922, n_1465, n_6914);
  nand g176970 (n_6921, n_7046, n_6303);
  nand g176971 (n_6920, n_7046, n_6301);
  nand g176978 (n_6919, n_4774, n_6793);
  nand g176991 (n_6918, g479, n_9257);
  nand g177031 (n_6917, n_2054, n_6901);
  nand g176998 (n_6916, n_4570, n_6284);
  nand g177004 (n_6915, g35, n_6914);
  nand g177006 (n_6913, n_6279, n_5020);
  nand g177012 (n_6912, g35, n_6792);
  nand g177013 (n_6911, n_5905, n_6229);
  nor g176524 (n_7206, n_9257, n_6419);
  nand g176779 (n_7095, n_4423, n_6910);
  nand g176788 (n_7096, n_5371, n_6891);
  nand g176786 (n_7336, n_5373, n_6299);
  nand g176525 (n_7316, g287, n_6816);
  not g176882 (n_7325, n_6909);
  fflopd g482_reg(.CK (clock), .D (n_6320), .Q (g482));
  not g176888 (n_7237, n_7178);
  not g176887 (n_7230, n_7185);
  nand g177064 (n_6908, n_5908, n_6221);
  nand g177068 (n_6907, n_1370, n_6191);
  nand g177074 (n_6906, g3457, n_6289);
  nand g177075 (n_6905, g3462, n_6276);
  nand g177077 (n_6904, n_5903, n_6262);
  nand g177078 (n_6903, g3476, n_6189);
  nand g177081 (n_6902, n_1793, n_6901);
  nand g177084 (n_6900, n_1804, n_6901);
  nand g177086 (n_6899, g5134, n_6199);
  nand g177089 (n_6898, n_5899, n_6234);
  nand g177091 (n_6897, g1772, n_6901);
  nand g177104 (n_6896, n_5889, n_6256);
  nand g177109 (n_6895, g2040, n_6443);
  nand g177116 (n_6894, g5120, n_6269);
  nand g177121 (n_6893, g5115, n_6294);
  nor g177127 (n_6892, n_6890, n_6891);
  nand g176346 (n_6889, n_6438, n_6888);
  nand g176344 (n_6887, n_6886, n_6405);
  nand g176342 (n_6885, n_6884, n_6410);
  nand g176341 (n_6883, n_6881, n_6402);
  nand g176340 (n_6882, n_6440, n_6881);
  nand g176332 (n_6880, n_4646, n_6409);
  not g177192 (n_6879, n_6487);
  nor g176330 (n_6878, g2399, n_6448);
  nand g177236 (n_6877, g2815, n_8413);
  nand g177297 (n_6875, n_4566, n_6296);
  nor g177326 (n_6874, n_5517, n_6298);
  nand g177350 (n_6873, new_g10383_, n_6926);
  nand g177366 (n_6872, n_5277, n_6218);
  nand g177405 (n_6871, n_6216, n_5861);
  nor g176326 (n_6870, g2667, n_6447);
  not g177628 (n_6869, n_6476);
  not g177631 (n_6868, n_6473);
  nand g175916 (n_6866, g2533, n_6847);
  nand g177729 (n_6865, g2819, n_8413);
  nand g177790 (n_6864, g2771, n_8413);
  nand g177827 (n_6863, g2775, n_8413);
  nand g177859 (n_6862, g2783, n_8413);
  nand g177876 (n_6861, g2787, n_8413);
  nand g177893 (n_6860, g2803, n_8413);
  nand g177908 (n_6859, g2807, n_8413);
  not g177963 (n_6858, n_6857);
  not g175893 (n_6856, n_6460);
  nand g176316 (n_6855, n_6356, n_1952);
  not g175890 (n_6854, n_6449);
  not g175892 (n_6853, n_6579);
  nand g175911 (n_6852, g2667, n_6850);
  nand g175912 (n_6851, g2648, n_6850);
  nand g175913 (n_6849, g2567, n_6850);
  nand g175914 (n_6848, g2541, n_6847);
  nand g175915 (n_6846, g2537, n_6847);
  nand g175917 (n_6845, g2514, n_6847);
  nand g175918 (n_6844, g2433, n_6847);
  nand g175924 (n_6843, n_6437, n_481);
  nand g176308 (n_6841, n_6363, n_2869);
  nand g176307 (n_6840, n_6364, n_2978);
  nand g176299 (n_6839, n_6399, n_6454);
  nand g176298 (n_6838, n_6401, n_6456);
  nand g176297 (n_6837, n_6403, n_6450);
  nand g176291 (n_6836, g2407, n_6834);
  nand g176290 (n_6835, g2403, n_6834);
  nand g176289 (n_6833, g2399, n_6834);
  nand g175951 (n_6832, n_4452, n_6818);
  nand g176288 (n_6831, g2380, n_6834);
  nand g176287 (n_6830, g2299, n_6834);
  nand g176286 (n_6829, g2273, n_6826);
  nand g175952 (n_6828, n_3720, n_6426);
  nand g176285 (n_6827, g2269, n_6826);
  nand g176284 (n_6825, g2265, n_6826);
  nand g176283 (n_6824, g2246, n_6826);
  nand g176282 (n_6823, g4045, n_5758);
  nand g175955 (n_6822, g5348, n_4334);
  nand g175956 (n_6821, g4045, n_4335);
  nand g175957 (n_6820, g3343, n_4336);
  nand g175966 (n_6819, n_4808, n_6818);
  nor g175972 (n_6817, n_6814, n_6816);
  nand g175973 (n_6815, n_6814, n_6816);
  nand g176280 (n_6813, g3343, n_3773);
  nand g176278 (n_6812, g2165, n_6826);
  nand g176270 (n_6811, g5348, n_3767);
  nand g176262 (n_6810, g1454, n_6442);
  nand g176261 (n_6809, g2675, n_6850);
  not g176180 (n_6808, n_6504);
  not g176181 (n_6807, n_6505);
  not g176191 (n_6806, n_6786);
  not g176190 (n_6805, n_6787);
  not g176195 (n_6804, n_6784);
  not g176196 (n_6803, n_6780);
  not g176205 (n_6802, n_6778);
  not g176206 (n_6801, n_6777);
  not g176212 (n_6800, n_6773);
  not g176211 (n_6799, n_6774);
  not g176216 (n_6798, n_6772);
  not g176223 (n_6797, n_6770);
  not g176224 (n_6796, n_6769);
  not g176228 (n_6795, n_6768);
  nand g176260 (n_6794, g2671, n_6850);
  nand g177155 (n_7097, g1862, n_6793);
  nor g175988 (n_7151, g1636, n_6446);
  nand g177136 (n_7157, n_1031, n_6793);
  nand g177139 (n_7155, n_219, n_6914);
  nand g177142 (n_7153, g2070, n_6792);
  nand g177148 (n_7098, n_6016, n_6791);
  nor g177135 (n_7159, n_2894, n_6257);
  fflopd g5212_reg(.CK (clock), .D (n_6295), .Q (g5212));
  fflopd g5077_reg(.CK (clock), .D (n_6397), .Q (g5077));
  fflopd g1046_reg(.CK (clock), .D (n_6293), .Q (g1046));
  nand g177435 (n_7333, g744, n_6219);
  fflopd g5559_reg(.CK (clock), .D (n_6282), .Q (g5559));
  fflopd g5905_reg(.CK (clock), .D (n_6283), .Q (g5905));
  fflopd g3905_reg(.CK (clock), .D (n_6291), .Q (g3905));
  fflopd g3554_reg(.CK (clock), .D (n_6290), .Q (g3554));
  fflopd g3203_reg(.CK (clock), .D (n_6288), .Q (g3203));
  fflopd g6597_reg(.CK (clock), .D (n_6286), .Q (g6597));
  fflopd g6251_reg(.CK (clock), .D (n_6285), .Q (g6251));
  fflopd g5022_reg(.CK (clock), .D (n_6197), .Q (g5022));
  fflopd g4332_reg(.CK (clock), .D (n_6188), .Q (new_g12440_));
  fflopd g1312_reg(.CK (clock), .D (n_6212), .Q (g1312));
  not g177211 (n_8296, g2735);
  fflopd g969_reg(.CK (clock), .D (n_6203), .Q (g969));
  fflopd g1514_reg(.CK (clock), .D (n_6287), .Q (g1514));
  fflopd g79_reg(.CK (clock), .D (n_6280), .Q (g20899));
  fflopd g1526_reg(.CK (clock), .D (n_6193), .Q (g1526));
  fflopd g4776_reg(.CK (clock), .D (n_6196), .Q (g4776));
  fflopd g837_reg(.CK (clock), .D (n_6278), .Q (g837));
  fflopd g1500_reg(.CK (clock), .D (n_6277), .Q (g7946));
  nand g176620 (n_6790, n_1201, n_6093);
  nand g176381 (n_6789, n_1738, n_6141);
  nand g176383 (n_6788, g2495, n_6154);
  nand g176387 (n_6787, n_6152, n_4470);
  nand g176388 (n_6786, g5694, n_4472);
  nand g176393 (n_6785, g2509, n_6782);
  nand g176394 (n_6784, n_6150, n_4491);
  nand g176395 (n_6783, g2527, n_6782);
  nand g176396 (n_6781, g35, n_6169);
  nand g176397 (n_6780, g6040, n_4474);
  nand g176409 (n_6779, g2643, n_6775);
  nand g176410 (n_6778, n_6151, n_4493);
  nand g176411 (n_6777, g6386, n_4476);
  nand g176412 (n_6776, g2661, n_6775);
  nand g176419 (n_6774, n_6146, n_4489);
  nand g176420 (n_6773, g6732, n_4484);
  nand g176425 (n_6772, n_3303, n_6135);
  nand g176712 (n_6771, n_835, n_5972);
  nand g176434 (n_6770, n_6148, n_4456);
  nand g176435 (n_6769, g3694, n_4479);
  nand g176445 (n_6768, n_1069, n_6178);
  nand g176452 (n_6767, g827, n_6143);
  nand g176453 (n_6766, n_3586, n_6126);
  nand g176711 (n_6765, n_1262, n_5973);
  fflopd g1_reg(.CK (clock), .D (n_6063), .Q (g12832));
  nand g176481 (n_6764, n_1853, n_6118);
  nand g176482 (n_6763, g2227, n_6153);
  nand g176490 (n_6762, g2241, n_6760);
  nand g176491 (n_6761, g2259, n_6760);
  nand g176493 (n_6759, g35, n_6180);
  nand g176506 (n_6758, g2375, n_6756);
  nand g176508 (n_6757, g2393, n_6756);
  nor g176513 (n_6755, n_6168, n_4471);
  nor g176515 (n_6754, n_5476, n_6160);
  nor g176710 (n_6753, n_6752, n_6184);
  not g176541 (n_6751, g5348);
  not g176543 (n_6750, g3343);
  not g176544 (n_6749, g4045);
  nor g176551 (n_6748, g1848, n_6444);
  nor g176552 (n_6747, n_4524, n_6516);
  nor g176554 (n_6746, g1361, n_6522);
  nand g176572 (n_6740, n_1915, n_6069);
  nand g176576 (n_6739, n_5361, n_5942);
  nand g176577 (n_6738, n_5363, n_5984);
  nand g176578 (n_6737, n_5365, n_6005);
  nand g176579 (n_6736, n_5366, n_6023);
  nand g176580 (n_6735, n_5364, n_6098);
  nor g176582 (n_6734, n_6017, n_6186);
  nand g176584 (n_6733, n_2132, n_5915);
  nand g176585 (n_6732, n_1365, n_6171);
  nor g176586 (n_6731, g17316, n_6064);
  nand g176588 (n_6730, n_1296, n_5920);
  nand g176589 (n_6729, n_1142, n_5921);
  nand g176590 (n_6728, n_566, n_5922);
  nand g176591 (n_6727, n_1331, n_5923);
  nand g176592 (n_6726, n_6179, n_6307);
  nand g176593 (n_6725, n_516, n_5924);
  nand g176594 (n_6724, n_553, n_6025);
  nand g176595 (n_6723, n_1403, n_5925);
  nand g176596 (n_6722, n_755, n_5926);
  nand g176597 (n_6721, n_798, n_5927);
  nand g176598 (n_6720, n_733, n_5928);
  nand g176600 (n_6719, n_697, n_5929);
  nand g176601 (n_6718, n_548, n_5930);
  nand g176602 (n_6717, n_1338, n_5931);
  nand g176603 (n_6716, n_708, n_5932);
  nand g176604 (n_6715, n_642, n_6004);
  nand g176605 (n_6714, n_861, n_5933);
  nand g176606 (n_6713, n_574, n_5934);
  nand g176607 (n_6712, n_588, n_5935);
  nand g176611 (n_6711, n_1232, n_6081);
  nand g176612 (n_6710, n_1117, n_6082);
  nand g176613 (n_6709, n_783, n_6084);
  nand g176614 (n_6708, n_1127, n_6085);
  nand g176615 (n_6707, n_579, n_6088);
  nand g176616 (n_6706, n_1214, n_6089);
  nand g176617 (n_6705, n_561, n_6091);
  nand g176618 (n_6704, n_1243, n_5937);
  nand g176619 (n_6703, n_832, n_6092);
  nor g176367 (n_6702, n_5479, n_6161);
  nand g176621 (n_6701, n_784, n_6094);
  nand g176622 (n_6700, n_1278, n_6095);
  nand g176623 (n_6699, n_1150, n_6096);
  nand g176625 (n_6698, n_713, n_6109);
  nand g176626 (n_6697, n_684, n_6100);
  nand g176627 (n_6696, n_740, n_5983);
  nand g176629 (n_6695, n_1303, n_6102);
  nand g176630 (n_6694, n_1279, n_6027);
  nand g176631 (n_6693, n_498, n_6040);
  nand g176632 (n_6692, n_1002, n_6039);
  nand g176633 (n_6691, n_1244, n_6038);
  nand g176634 (n_6690, n_1249, n_6037);
  nand g176636 (n_6689, n_984, n_6036);
  nand g176637 (n_6688, n_1364, n_6035);
  nand g176638 (n_6687, n_771, n_6034);
  nand g176639 (n_6686, n_1259, n_6101);
  nand g176640 (n_6685, n_888, n_6033);
  nand g176641 (n_6684, n_1171, n_6032);
  nand g176642 (n_6683, n_928, n_6031);
  nand g176643 (n_6682, n_799, n_6030);
  nand g176644 (n_6681, n_1241, n_5962);
  nand g176645 (n_6680, n_1390, n_6029);
  nand g176646 (n_6679, n_1361, n_6028);
  nand g176647 (n_6678, n_952, n_6026);
  nand g176649 (n_6677, n_541, n_6022);
  nand g176650 (n_6676, n_1178, n_6021);
  nand g176651 (n_6675, n_674, n_6020);
  nand g176652 (n_6674, n_1110, n_6041);
  nand g176653 (n_6673, n_1359, n_6103);
  nand g176654 (n_6672, n_668, n_6042);
  nand g176655 (n_6671, n_1113, n_6043);
  nand g176656 (n_6670, n_1228, n_6044);
  nand g176657 (n_6669, n_1038, n_6045);
  nand g176658 (n_6668, n_833, n_6046);
  nand g176659 (n_6667, n_675, n_6047);
  nand g176660 (n_6666, n_1392, n_6048);
  nand g176661 (n_6665, n_1238, n_6071);
  nand g176663 (n_6664, n_1183, n_6075);
  nand g176664 (n_6663, n_754, n_6076);
  nand g176665 (n_6662, n_514, n_6077);
  nand g176666 (n_6661, n_1118, n_6078);
  nand g176667 (n_6660, n_1393, n_6170);
  nand g176668 (n_6659, n_1270, n_5941);
  nand g176669 (n_6658, n_518, n_6105);
  nand g176670 (n_6657, n_1097, n_6106);
  nand g176671 (n_6656, n_1305, n_6107);
  nand g176672 (n_6655, n_747, n_6108);
  nand g176673 (n_6654, n_870, n_6110);
  nand g176674 (n_6653, n_937, n_6111);
  nand g176675 (n_6652, n_939, n_6099);
  nand g176676 (n_6651, n_655, n_5914);
  nand g176677 (n_6650, n_780, n_6007);
  nand g176678 (n_6649, n_2052, n_6647);
  nand g176680 (n_6648, n_4912, n_6647);
  nand g176681 (n_6646, n_965, n_6003);
  nand g176682 (n_6645, n_660, n_6002);
  nand g176683 (n_6644, n_656, n_6001);
  nand g176684 (n_6643, n_818, n_6000);
  nand g176685 (n_6642, n_854, n_5999);
  nand g176686 (n_6641, n_815, n_5998);
  nand g176687 (n_6640, n_564, n_5997);
  nand g176688 (n_6639, n_1184, n_5996);
  nand g176689 (n_6638, n_1245, n_5995);
  nand g176690 (n_6637, n_997, n_5994);
  nand g176691 (n_6636, n_537, n_5993);
  nand g176692 (n_6635, n_1335, n_5992);
  nand g176693 (n_6634, n_526, n_5991);
  nand g176694 (n_6633, n_950, n_5990);
  nand g176695 (n_6632, n_1254, n_5989);
  nand g176696 (n_6631, n_874, n_5988);
  nand g176698 (n_6630, n_494, n_5987);
  nand g176699 (n_6629, n_559, n_5986);
  nand g176701 (n_6628, n_608, n_5982);
  nand g176702 (n_6627, n_1125, n_5981);
  nand g176703 (n_6626, n_529, n_5980);
  nand g176704 (n_6625, n_1285, n_5979);
  nand g176705 (n_6624, n_1286, n_5978);
  nand g176706 (n_6623, n_1233, n_5977);
  nand g176707 (n_6622, n_1326, n_5976);
  nand g176708 (n_6621, n_765, n_5975);
  nand g176709 (n_6620, n_988, n_5974);
  fflopd g4176_reg(.CK (clock), .D (n_6066), .Q (g4176));
  fflopd g2882_reg(.CK (clock), .D (n_6144), .Q (g2882));
  fflopd g4388_reg(.CK (clock), .D (n_6124), .Q (g4388));
  nor g176343 (n_6619, n_6130, n_1413);
  nand g176714 (n_6618, n_1119, n_5970);
  nand g176715 (n_6617, n_1264, n_5969);
  nand g176716 (n_6616, n_1231, n_5968);
  nand g176717 (n_6615, n_520, n_5967);
  nand g176718 (n_6614, n_917, n_5966);
  nand g176719 (n_6613, n_829, n_5965);
  nand g176722 (n_6612, n_1024, n_6173);
  nand g176723 (n_6611, n_503, n_5961);
  nand g176724 (n_6610, n_643, n_5960);
  nand g176725 (n_6609, n_777, n_5959);
  nand g176726 (n_6608, n_1386, n_5958);
  nand g176727 (n_6607, n_1145, n_5957);
  nand g176728 (n_6606, n_943, n_5956);
  nand g176729 (n_6605, n_915, n_5955);
  nand g176730 (n_6604, n_923, n_5954);
  nand g176731 (n_6603, n_944, n_5953);
  nand g176732 (n_6602, n_748, n_5952);
  nand g176733 (n_6601, n_1280, n_5951);
  nand g176734 (n_6600, n_769, n_5950);
  nand g176735 (n_6599, n_1258, n_5949);
  nand g175940 (n_6598, n_1520, n_6503);
  nand g176736 (n_6597, n_947, n_5948);
  nand g176737 (n_6596, n_766, n_5947);
  nand g176738 (n_6595, n_1013, n_5946);
  nand g176739 (n_6594, n_1168, n_5945);
  nand g176740 (n_6593, n_868, n_5944);
  nand g176744 (n_6592, n_659, n_6086);
  nand g176745 (n_6591, n_1272, n_5938);
  nand g176749 (n_6590, n_739, n_6174);
  nand g176750 (n_6589, n_670, n_6090);
  nand g176752 (n_6588, n_1389, n_5939);
  nand g176753 (n_6587, n_951, n_6087);
  nand g176756 (n_6586, n_1121, n_6172);
  nand g176757 (n_6585, n_940, n_6083);
  nand g176713 (n_6584, n_706, n_5971);
  nand g176315 (n_6583, n_6582, n_6157);
  nand g176314 (n_6581, n_6580, n_6166);
  nand g175948 (n_6579, n_6145, n_4325);
  not g176834 (n_6578, n_6348);
  not g176835 (n_6577, n_6347);
  not g176848 (n_6576, n_6389);
  not g176862 (n_6575, n_6574);
  not g176867 (n_6573, n_6572);
  not g176868 (n_6571, n_6570);
  not g176870 (n_6569, n_6568);
  not g176871 (n_6567, n_6566);
  not g176873 (n_6565, n_6564);
  nand g176313 (n_6563, n_6562, n_6158);
  nand g176312 (n_6561, n_6560, n_6155);
  nand g176311 (n_6559, n_1011, n_6176);
  wire w35, w36, w37, w38;
  nand g176891 (n_6558, w36, w38);
  nand g44 (w38, w37, n_962);
  not g43 (w37, n_5874);
  nand g42 (w36, w35, n_5874);
  not g41 (w35, n_962);
  nand g176901 (n_6557, n_1019, n_6067);
  nand g176923 (n_6556, n_5358, n_6104);
  nand g176925 (n_6555, n_5362, n_5963);
  nand g176929 (n_6554, n_5359, n_6080);
  nand g176932 (n_6553, n_2920, n_6050);
  nor g176933 (n_6552, g1772, n_6183);
  nand g176935 (n_6551, n_1994, n_6049);
  nand g176943 (n_6550, n_2619, n_6051);
  nand g176944 (n_6549, g2555, n_6547);
  nand g176945 (n_6548, g2599, n_6547);
  nand g176946 (n_6546, g2629, n_6547);
  nand g176947 (n_6545, g2643, n_6547);
  nand g176952 (n_6544, g2287, n_6542);
  nand g176953 (n_6543, g2331, n_6542);
  nand g176954 (n_6541, g2361, n_6542);
  nand g176955 (n_6540, g2375, n_6542);
  nand g176965 (n_6539, n_6011, n_6058);
  nand g176966 (n_6538, n_6019, n_6054);
  nor g176976 (n_6537, n_4653, n_6445);
  nand g176995 (n_6536, g18881, n_9257);
  nand g177017 (n_6535, g2421, n_6533);
  nand g177018 (n_6534, g2465, n_6533);
  nand g177019 (n_6532, g2495, n_6533);
  nand g177020 (n_6531, g2509, n_6533);
  nand g177026 (n_6530, g2153, n_6528);
  nand g177027 (n_6529, g2197, n_6528);
  nand g177028 (n_6527, g2227, n_6528);
  nand g177029 (n_6526, g2241, n_6528);
  nand g177043 (n_6525, g1070, n_5888);
  nand g177054 (n_6524, n_4128, n_6053);
  nand g177055 (n_6523, g1361, n_6522);
  nand g177057 (n_6521, n_5885, n_5725);
  nand g177058 (n_6520, n_5884, n_5727);
  nand g177060 (n_6519, n_5882, n_5728);
  nand g176309 (n_6518, n_1005, n_6175);
  nand g177083 (n_6517, g35, n_6516);
  nand g177092 (n_6515, n_4092, n_5897);
  nand g177097 (n_6514, n_3972, n_6068);
  nand g175930 (n_6513, n_6512, n_6394);
  nand g177105 (n_6511, g2012, n_6300);
  nand g177107 (n_6510, g2020, n_6302);
  nand g177108 (n_6509, g2024, n_6304);
  nor g176306 (n_6508, n_6167, n_2615);
  nand g176305 (n_6507, n_484, n_6164);
  nand g176303 (n_6506, n_911, n_6165);
  nand g176302 (n_6505, n_6309, n_6501);
  nand g176301 (n_6504, n_6311, n_6503);
  nand g175938 (n_6502, n_1488, n_6501);
  not g177202 (n_6500, n_6499);
  nor g176300 (n_6498, n_6114, n_5462);
  nor g176296 (n_6497, n_6128, n_5464);
  nor g176295 (n_6496, n_6129, n_4444);
  nand g177299 (n_6493, n_4828, n_5854);
  nor g177305 (n_6492, g744, n_6472);
  nand g177312 (n_6490, n_5853, n_5840);
  nand g177313 (n_6489, n_5342, n_5851);
  nor g177317 (n_6488, n_4878, n_6182);
  nand g177336 (n_6487, n_1354, n_5870);
  nor g177354 (n_6486, g2807, n_6485);
  nor g177357 (n_6484, g2775, n_6485);
  nand g177358 (n_6483, n_3308, n_5875);
  nand g177365 (n_6482, n_715, n_5865);
  nand g177379 (n_6479, n_5877, n_5550);
  nand g175937 (n_6478, n_1671, n_6501);
  fflopd g2735_reg(.CK (clock), .D (n_5859), .Q (g2735));
  not g177648 (n_6477, n_6198);
  nand g177854 (n_6476, n_851, n_5871);
  nand g177855 (n_6475, g35, n_6474);
  nand g177862 (n_6473, g744, n_6472);
  nor g177872 (n_6471, g2771, n_6468);
  nand g177878 (n_6470, n_2062, n_5867);
  nor g177883 (n_6469, g2803, n_6468);
  nand g177896 (n_6467, g146, n_6217);
  nand g178135 (n_6466, g5052, n_5879);
  nor g176294 (n_6465, n_6134, n_1409);
  nand g175923 (n_6464, n_6463, n_6392);
  nand g175939 (n_6462, n_1684, n_6503);
  nor g176293 (n_6461, n_6136, n_5466);
  nand g175949 (n_6460, n_6147, n_4327);
  nand g176281 (n_6459, g3694, n_5760);
  nand g176279 (n_6458, g6732, n_3769);
  nand g176273 (n_6457, g6386, n_6456);
  nand g176272 (n_6455, g6040, n_6454);
  nor g175964 (n_6453, g676, n_6312);
  nand g177267 (g28030, n_4764, n_5855);
  nand g176271 (n_6451, g5694, n_6450);
  nand g175944 (n_6449, n_6149, n_4323);
  fflopd g4366_reg(.CK (clock), .D (n_5940), .Q (g4366));
  not g176876 (n_7088, n_6448);
  not g176878 (n_7086, n_6447);
  not g176879 (n_7039, n_6446);
  nand g178180 (n_6857, g5052, n_5881);
  nor g177134 (n_6933, g2040, n_6185);
  nand g177156 (n_6909, g35, n_6445);
  nand g177162 (n_7185, g35, n_6444);
  nor g177146 (n_7040, g1668, n_6445);
  nand g177163 (n_7178, g35, n_6187);
  fflopd g732_reg(.CK (clock), .D (n_6181), .Q (g732));
  not g177220 (n_7094, n_6793);
  fflopd g4664_reg(.CK (clock), .D (n_6070), .Q (g4664));
  fflopd g4322_reg(.CK (clock), .D (n_6052), .Q (g4322));
  not g177218 (n_7144, n_6443);
  fflopd g4311_reg(.CK (clock), .D (n_5896), .Q (g4311));
  fflopd g5016_reg(.CK (clock), .D (n_5873), .Q (g5016));
  fflopd g812_reg(.CK (clock), .D (n_5893), .Q (g812));
  fflopd g278_reg(.CK (clock), .D (n_5936), .Q (g278));
  fflopd g827_reg(.CK (clock), .D (n_6142), .Q (g827));
  fflopd g1056_reg(.CK (clock), .D (n_5917), .Q (g19334));
  not g177223 (n_7133, n_6901);
  fflopd g4473_reg(.CK (clock), .D (n_6065), .Q (new_g6961_));
  fflopd g4392_reg(.CK (clock), .D (n_6062), .Q (g4392));
  fflopd g4975_reg(.CK (clock), .D (n_5860), .Q (g4975));
  fflopd g528_reg(.CK (clock), .D (n_5904), .Q (new_g8038_));
  fflopd g4584_reg(.CK (clock), .D (n_5862), .Q (g4584));
  nand g176924 (n_6442, n_6441, n_5624);
  not g176538 (n_6440, g6386);
  not g176539 (n_6439, g6040);
  not g176540 (n_6438, g5694);
  not g176547 (n_6437, g3694);
  nand g176553 (n_6436, g2661, n_6378);
  nand g176558 (n_6435, n_2758, n_5774);
  nand g176561 (n_6434, n_2726, n_5777);
  nand g176563 (n_6433, n_2862, n_5779);
  nand g176566 (n_6432, n_151, n_5784);
  nand g176568 (n_6431, n_2750, n_5780);
  nand g176569 (n_6430, n_6429, n_6424);
  nand g176570 (n_6428, n_6427, n_6422);
  nand g176573 (n_6426, n_6177, n_5732);
  nand g176609 (n_6425, n_2324, n_6424);
  nand g176635 (n_6423, n_2237, n_6422);
  nand g176662 (n_6421, n_5486, n_6306);
  nand g176748 (n_6419, n_144, n_6387);
  nand g177124 (n_6417, g2197, n_6415);
  nand g177122 (n_6416, n_1764, n_6415);
  nand g177117 (n_6414, n_1795, n_6415);
  nand g177115 (n_6413, g6035, n_5590);
  not g176836 (n_6412, n_6139);
  not g176837 (n_6411, n_6138);
  not g176840 (n_6410, n_6137);
  not g176841 (n_6409, n_6133);
  not g176843 (n_6408, n_6132);
  not g176844 (n_6407, n_6131);
  not g176845 (n_6406, n_6127);
  not g176846 (n_6405, n_6125);
  not g176852 (n_6404, n_6123);
  not g176853 (n_6403, n_6122);
  not g176854 (n_6402, n_6121);
  not g176855 (n_6401, n_6120);
  not g176856 (n_6400, n_6119);
  not g176857 (n_6399, n_6116);
  not g176859 (n_6398, n_6115);
  not g176860 (n_6397, n_6113);
  not g176861 (n_6396, n_6112);
  nand g177110 (n_6391, g5689, n_5566);
  nand g177106 (n_6390, g5467, n_5768);
  nand g177103 (n_6389, n_1339, n_5796);
  nand g177102 (n_6388, g4392, n_6387);
  nand g177098 (n_6386, g6500, n_5684);
  nand g176893 (n_6385, g2393, n_6368);
  nand g176896 (n_6384, n_4748, n_5823);
  nand g176897 (n_6383, n_6512, n_5831);
  nand g176898 (n_6382, n_4749, n_5729);
  nand g176906 (n_6381, n_5826, n_1026);
  nand g176907 (n_6380, n_6463, n_5839);
  nand g176908 (n_6379, n_6512, n_6378);
  nand g176910 (n_6377, n_5744, n_3627);
  nand g176911 (n_6376, n_5742, n_5154);
  nand g176912 (n_6375, n_6463, n_5837);
  nand g176915 (n_6374, n_5739, n_5152);
  nand g176916 (n_6373, n_5736, n_5150);
  nand g176917 (n_6372, n_5735, n_5148);
  nand g176918 (n_6371, n_5733, n_3272);
  nand g176919 (n_6370, n_6463, n_5835);
  nand g176920 (n_6369, n_6463, n_6368);
  nand g176921 (n_6367, n_4988, n_5762);
  not g176536 (n_6366, g6732);
  nand g176934 (n_6365, n_5740, g25114);
  nand g176939 (n_6364, n_5737, n_5130);
  nand g176940 (n_6363, n_5743, n_5128);
  nand g176957 (n_6362, n_6361, n_5567);
  nand g176958 (n_6360, n_6359, n_5565);
  nand g176959 (n_6358, n_6357, n_5591);
  nand g176960 (n_6356, n_6361, n_5741);
  nand g176967 (n_6355, n_1642, n_6342);
  nand g176969 (n_6354, n_1462, n_6339);
  nand g176974 (n_6353, n_6352, n_5628);
  nand g176979 (n_6351, n_6350, n_5596);
  nand g176981 (n_6349, n_6512, n_5833);
  nand g176982 (n_6348, n_5788, n_2974);
  nand g176983 (n_6347, n_5791, n_2975);
  nand g176986 (n_6346, g872, n_9257);
  nand g176999 (n_6345, g35, n_6308);
  nand g177002 (n_6344, n_6512, n_5829);
  nand g177003 (n_6343, g35, n_6342);
  nand g177008 (n_6341, g5481, n_5570);
  nand g177014 (n_6340, g35, n_6339);
  nand g177015 (n_6338, g35, n_6313);
  nand g177021 (n_6337, g872, n_5795);
  nand g177030 (n_6336, n_2051, n_6332);
  nand g177032 (n_6335, n_2058, n_6415);
  nand g177033 (n_6334, g5462, n_5592);
  nand g177034 (n_6333, n_2034, n_6332);
  nand g177036 (n_6331, n_1868, n_6332);
  nand g177037 (n_6330, g2465, n_6332);
  nand g177038 (n_6329, g5808, n_5816);
  nand g177039 (n_6328, g5813, n_5785);
  nand g177041 (n_6327, g5827, n_5651);
  nand g177050 (n_6326, g6505, n_5771);
  nand g177052 (n_6325, g6519, n_5669);
  nand g177053 (n_6324, g2599, n_6010);
  nand g177062 (n_6323, g3106, n_5730);
  nand g177063 (n_6322, g3111, n_5778);
  nand g177065 (n_6321, g3125, n_5745);
  nand g177067 (n_6320, n_1213, n_5820);
  nand g177069 (n_6319, g2331, n_6009);
  nand g177070 (n_6318, g3689, n_5569);
  nand g177079 (n_6317, g4040, n_5568);
  nand g177087 (n_6316, g3808, n_5627);
  nand g177088 (n_6315, g3813, n_5775);
  nand g177090 (n_6314, g3827, n_5625);
  nand g177141 (n_6566, g2361, n_6313);
  not g176875 (n_6818, n_6312);
  fflopd g316_reg(.CK (clock), .D (n_5696), .Q (g316));
  nand g177132 (n_6574, n_6311, n_6342);
  nand g177137 (n_6572, g25259, n_6310);
  nand g177138 (n_6570, n_2124, n_6310);
  nand g177140 (n_6568, n_6309, n_6339);
  nand g177150 (n_6446, g1592, n_6310);
  nand g177143 (n_6564, g2629, n_6308);
  nand g177147 (n_6448, n_5381, n_6307);
  nand g177149 (n_6447, n_5383, n_6306);
  fflopd g5348_reg(.CK (clock), .D (n_5571), .Q (g5348));
  fflopd g4045_reg(.CK (clock), .D (n_5603), .Q (g4045));
  nor g176762 (n_6816, n_4689, n_5594);
  fflopd g3343_reg(.CK (clock), .D (n_5653), .Q (g3343));
  fflopd g5062_reg(.CK (clock), .D (n_5519), .Q (g5062));
  not g176890 (n_6847, n_6782);
  not g176889 (n_6850, n_6775);
  not g176886 (n_6826, n_6760);
  not g176885 (n_6834, n_6756);
  fflopd g4005_reg(.CK (clock), .D (n_5753), .Q (g11418));
  nor g177159 (n_8107, n_9257, n_5769);
  not g177197 (n_6305, n_6304);
  not g177198 (n_6303, n_6302);
  not g177199 (n_6301, n_6300);
  not g177203 (n_6299, n_6522);
  nor g178348 (n_6298, n_5880, n_5516);
  not g178244 (n_6296, n_5907);
  nand g177254 (n_6295, n_3663, n_5527);
  nand g177255 (n_6294, g35, n_5553);
  nand g177256 (n_6293, n_4897, n_5528);
  nand g177259 (n_6292, g35, n_5547);
  nand g177260 (n_6291, n_3662, n_5530);
  nand g177261 (n_6290, n_3633, n_5531);
  nand g177262 (n_6289, g35, n_5544);
  nand g177263 (n_6288, n_3688, n_5533);
  nand g177264 (n_6287, n_2821, n_6192);
  nand g177266 (n_6286, n_3689, n_5537);
  nand g177269 (n_6285, n_3636, n_5538);
  nand g177270 (n_6284, g35, n_5561);
  nand g177271 (n_6283, n_3634, n_5539);
  nand g177273 (n_6282, n_3639, n_5540);
  nor g177291 (n_6281, n_5526, n_3354);
  nand g177294 (n_6280, n_4418, n_5535);
  nor g177303 (n_6279, n_1539, n_5557);
  nand g177309 (n_6278, n_1394, n_5529);
  nand g177316 (n_6277, n_4921, n_5534);
  nor g177320 (n_6276, g3457, n_6274);
  nor g177321 (n_6275, g3476, n_6274);
  nor g177322 (n_6273, g6154, n_6271);
  nor g177323 (n_6272, g6173, n_6271);
  nor g177324 (n_6270, g5134, n_6268);
  nor g177325 (n_6269, g5115, n_6268);
  nand g177330 (n_6267, g6173, n_6265);
  nand g177331 (n_6266, g6177, n_6265);
  nand g177332 (n_6264, g5124, n_6258);
  nand g177333 (n_6263, g3466, n_6261);
  nand g177334 (n_6262, g3476, n_6261);
  nand g177335 (n_6260, g3480, n_6261);
  nand g177337 (n_6259, g5138, n_6258);
  nand g177338 (n_6257, n_4167, n_5556);
  nand g177339 (n_6256, g5134, n_6258);
  nand g177340 (n_6255, g6163, n_6265);
  nand g177342 (n_6254, g6181, n_6265);
  nand g177347 (n_6253, g3484, n_6261);
  nand g177348 (n_6252, g5142, n_6258);
  nor g177351 (n_6251, g2819, n_6250);
  nor g177353 (n_6249, g2815, n_6248);
  nor g177355 (n_6247, g2787, n_6250);
  nor g177356 (n_6246, g2783, n_6248);
  nand g177381 (n_6245, n_5549, n_5521);
  nand g177383 (n_6244, g3133, n_6222);
  nand g177387 (n_6243, g5485, n_6241);
  nand g177388 (n_6242, g5489, n_6241);
  nand g177389 (n_6240, g5817, n_6238);
  nand g177390 (n_6239, g5827, n_6238);
  nand g177391 (n_6237, g5835, n_6238);
  nand g177392 (n_6236, g5831, n_6238);
  nand g177393 (n_6235, g3817, n_6233);
  nand g177394 (n_6234, g3827, n_6233);
  nand g177395 (n_6232, g3831, n_6233);
  nand g177396 (n_6231, g3835, n_6233);
  nand g177397 (n_6230, g5471, n_6241);
  nand g177398 (n_6229, g5481, n_6241);
  nand g177399 (n_6228, g6509, n_6226);
  nand g177400 (n_6227, g6519, n_6226);
  nand g177401 (n_6225, g6527, n_6226);
  nand g177402 (n_6224, g6523, n_6226);
  nand g177406 (n_6223, g3115, n_6222);
  nand g177407 (n_6221, g3125, n_6222);
  nand g177408 (n_6220, g3129, n_6222);
  not g177964 (n_6219, n_6472);
  not g177961 (n_6218, n_6217);
  not g177959 (n_6216, n_5863);
  not g177532 (n_6212, n_5913);
  not g177645 (n_6203, n_5891);
  nand g177907 (n_6199, g35, n_5554);
  nand g177900 (n_6198, n_3908, n_5524);
  nand g177899 (n_6197, n_3749, n_5508);
  nand g177880 (n_6196, n_4895, n_5847);
  nand g177694 (n_6195, g35, n_5506);
  nand g177704 (n_6194, g35, n_5548);
  nand g177760 (n_6193, n_3604, n_6192);
  nand g177765 (n_6191, g35, n_5523);
  nand g177778 (n_6190, g35, n_5513);
  nand g177792 (n_6189, g35, n_5545);
  nand g177861 (n_6188, n_2022, n_5522);
  not g177209 (n_6928, n_6187);
  not g177676 (n_6791, n_6186);
  not g177674 (n_6792, n_6185);
  not g177207 (n_6891, n_6184);
  nand g177483 (n_6443, g35, n_5558);
  nand g177427 (n_6499, g1542, n_5536);
  fflopd g479_reg(.CK (clock), .D (n_5512), .Q (g479));
  not g177213 (n_6946, n_6444);
  not g177678 (n_6910, n_6183);
  fflopd g6541_reg(.CK (clock), .D (n_5764), .Q (g6541));
  not g178282 (n_6926, n_6182);
  fflopd g728_reg(.CK (clock), .D (n_5542), .Q (g728));
  fflopd g645_reg(.CK (clock), .D (n_5659), .Q (g645));
  fflopd g6311_reg(.CK (clock), .D (n_5781), .Q (g6311));
  fflopd g6195_reg(.CK (clock), .D (n_5766), .Q (g6195));
  fflopd g4112_reg(.CK (clock), .D (n_5551), .Q (g4112));
  not g177679 (n_6914, n_6516);
  fflopd g6657_reg(.CK (clock), .D (n_5772), .Q (g6657));
  fflopd g4854_reg(.CK (clock), .D (n_5509), .Q (g4854));
  fflopd g718_reg(.CK (clock), .D (n_5842), .Q (g718));
  nand g177488 (n_6793, n_5660, n_5562);
  fflopd g661_reg(.CK (clock), .D (n_5507), .Q (g661));
  fflopd g4991_reg(.CK (clock), .D (n_5555), .Q (g4991));
  fflopd g681_reg(.CK (clock), .D (n_5514), .Q (g681));
  nand g177496 (n_6901, g35, n_5559);
  fflopd g655_reg(.CK (clock), .D (n_5515), .Q (g655));
  fflopd g4064_reg(.CK (clock), .D (n_5511), .Q (g4064));
  fflopd g5313_reg(.CK (clock), .D (n_5752), .Q (g12238));
  fflopd g4966_reg(.CK (clock), .D (n_5845), .Q (g4966));
  fflopd g3303_reg(.CK (clock), .D (n_5754), .Q (g11349));
  fflopd g269_reg(.CK (clock), .D (n_5782), .Q (g269));
  not g178291 (n_8413, n_6468);
  nand g176364 (n_6181, n_10369, n_5253);
  nor g176549 (n_6180, g2273, n_6014);
  nand g178474 (n_6179, n_4756, n_5285);
  nand g176574 (n_6178, n_6177, n_5731);
  nor g176581 (n_6176, n_5379, n_5666);
  nor g176583 (n_6175, n_5380, n_5663);
  not g177550 (n_6174, n_5672);
  not g177549 (n_6173, n_5673);
  not g177548 (n_6172, n_5674);
  not g177547 (n_6171, n_5675);
  not g177546 (n_6170, n_5676);
  nor g176894 (n_6169, g2541, n_6015);
  nor g176909 (n_6168, n_5433, n_4842);
  nor g176927 (n_6167, n_5413, n_1543);
  nand g176928 (n_6166, n_4171, n_5412);
  nor g176931 (n_6165, g2465, n_6013);
  nor g176936 (n_6164, g2197, n_6012);
  nor g176937 (n_6163, n_5432, n_4831);
  nor g176938 (n_6162, n_5423, n_1411);
  nor g176941 (n_6161, n_5408, n_2996);
  nor g176942 (n_6160, n_5430, n_6159);
  nand g176972 (n_6158, n_4170, n_5405);
  nand g176973 (n_6157, n_4623, n_5406);
  nor g176975 (n_6156, n_4832, n_5467);
  nand g176977 (n_6155, n_4169, n_5407);
  nor g176984 (n_6154, n_4879, n_6140);
  nor g176985 (n_6153, n_4876, n_6117);
  nand g176987 (n_6152, g5685, n_9257);
  nand g176988 (n_6151, g6377, n_9257);
  nand g176990 (n_6150, g6031, n_9257);
  nand g176992 (n_6149, g3329, n_9257);
  nand g176993 (n_6148, g3680, n_9257);
  nand g176994 (n_6147, g4031, n_9257);
  nand g176996 (n_6146, g6723, n_9257);
  nand g176997 (n_6145, g5339, n_9257);
  nand g177000 (n_6144, n_5327, n_5481);
  nand g177005 (n_6143, g35, n_5475);
  nand g177016 (n_6142, n_938, n_5482);
  nand g177035 (n_6141, g35, n_6140);
  nand g177044 (n_6139, g2571, n_5830);
  nand g177046 (n_6138, g2579, n_5832);
  nand g177059 (n_6137, g3329, g3195);
  nand g177061 (n_6136, g3329, g3211);
  nand g177066 (n_6135, n_5427, n_3310);
  nand g177071 (n_6134, g3680, g3562);
  nand g177072 (n_6133, g3680, g3546);
  nand g177076 (n_6132, g2583, n_5828);
  nand g177080 (n_6131, g2315, n_5838);
  nand g177082 (n_6130, g4031, g3897);
  nand g177085 (n_6129, g4031, g3913);
  nand g177093 (n_6128, g5339, g5220);
  nand g177094 (n_6127, g2311, n_5836);
  nand g177096 (n_6126, g35, n_5422);
  nand g177099 (n_6125, g5339, g5204);
  nand g177101 (n_6124, n_423, n_5421);
  nand g177111 (n_6123, g5685, g5551);
  nand g177112 (n_6122, g5685, g5567);
  nand g177113 (n_6121, g6377, g6243);
  nand g177114 (n_6120, g6377, g6259);
  nand g177118 (n_6119, g6031, g5897);
  nand g177119 (n_6118, g35, n_6117);
  nand g177120 (n_6116, g6031, g5913);
  nand g177125 (n_6115, g6723, g6589);
  nand g177126 (n_6114, g6723, g6605);
  nand g177130 (n_6113, g5073, n_4657);
  nand g177131 (n_6112, g2303, n_5834);
  not g177545 (n_6111, n_5677);
  not g177544 (n_6110, n_5678);
  not g177543 (n_6109, n_5679);
  not g177542 (n_6108, n_5680);
  not g177541 (n_6107, n_5681);
  not g177540 (n_6106, n_5682);
  not g177539 (n_6105, n_5683);
  not g177538 (n_6104, n_5685);
  not g177537 (n_6103, n_5686);
  not g177166 (n_6102, n_5819);
  not g177167 (n_6101, n_5818);
  not g177168 (n_6100, n_5817);
  not g177170 (n_6099, n_5815);
  not g177171 (n_6098, n_5814);
  not g177174 (n_6096, n_5812);
  not g177175 (n_6095, n_5811);
  not g177176 (n_6094, n_5810);
  not g177177 (n_6093, n_5809);
  not g177178 (n_6092, n_5808);
  not g177179 (n_6091, n_5807);
  not g177180 (n_6090, n_5806);
  not g177181 (n_6089, n_5805);
  not g177182 (n_6088, n_5804);
  not g177183 (n_6087, n_5803);
  not g177184 (n_6086, n_5802);
  not g177185 (n_6085, n_5801);
  not g177186 (n_6084, n_5800);
  not g177187 (n_6083, n_5799);
  not g177188 (n_6082, n_5798);
  not g177189 (n_6081, n_5797);
  not g177190 (n_6080, n_5793);
  not g177534 (n_6078, n_5688);
  not g177533 (n_6077, n_5689);
  not g177531 (n_6076, n_5690);
  not g177530 (n_6075, n_5691);
  nand g177226 (n_6074, g5821, n_5498);
  nand g177229 (n_6073, n_918, n_5404);
  nand g177234 (n_6072, n_2148, n_5456);
  not g177529 (n_6071, n_5692);
  nand g177258 (n_6070, n_3751, n_5331);
  nor g177272 (n_6069, n_1662, n_5314);
  nand g177292 (n_6068, n_8904, n_5315);
  nor g177293 (n_6067, g17404, n_5396);
  nand g177304 (n_6066, n_5525, n_2055);
  nand g177307 (n_6065, n_3109, n_5332);
  nand g177314 (n_6064, n_4592, n_5343);
  nand g177318 (n_6063, n_3345, n_6061);
  nand g177319 (n_6062, n_1402, n_6061);
  nor g177344 (n_6058, g1345, n_5502);
  nor g177352 (n_6054, g1002, n_6752);
  nand g177359 (n_6053, g305, n_5323);
  nand g177371 (n_6052, n_4969, n_5360);
  nand g177375 (n_6051, n_3512, n_5333);
  nor g177403 (n_6050, n_4153, n_5356);
  nor g177404 (n_6049, n_4017, n_5355);
  not g177528 (n_6048, n_5693);
  not g177527 (n_6047, n_5694);
  not g177526 (n_6046, n_5697);
  not g177525 (n_6045, n_5698);
  not g177524 (n_6044, n_5699);
  not g177523 (n_6043, n_5700);
  not g177522 (n_6042, n_5701);
  not g177521 (n_6041, n_5702);
  not g177499 (n_6040, n_5723);
  not g177500 (n_6039, n_5722);
  not g177501 (n_6038, n_5721);
  not g177502 (n_6037, n_5720);
  not g177503 (n_6036, n_5719);
  not g177504 (n_6035, n_5718);
  not g177505 (n_6034, n_5717);
  not g177506 (n_6033, n_5716);
  not g177507 (n_6032, n_5715);
  not g177508 (n_6031, n_5714);
  not g177509 (n_6030, n_5713);
  not g177510 (n_6029, n_5712);
  not g177511 (n_6028, n_5711);
  not g177512 (n_6027, n_5710);
  not g177513 (n_6026, n_5709);
  not g177514 (n_6025, n_5708);
  not g177517 (n_6023, n_5706);
  not g177518 (n_6022, n_5705);
  not g177519 (n_6021, n_5704);
  not g177520 (n_6020, n_5703);
  nand g177413 (n_6304, n_983, n_6018);
  nand g177438 (n_6184, n_6019, n_5372);
  nand g177415 (n_6300, n_1518, n_6018);
  nand g177414 (n_6302, n_6017, n_6018);
  nand g177461 (n_6187, n_6016, n_6018);
  nand g177145 (n_6312, g703, n_5425);
  nor g177144 (n_6392, g2331, n_5665);
  nor g177133 (n_6394, g2599, n_5664);
  nand g177471 (n_6444, n_1453, n_5849);
  fflopd g6386_reg(.CK (clock), .D (n_5434), .Q (g6386));
  fflopd g6040_reg(.CK (clock), .D (n_5435), .Q (g6040));
  not g177219 (n_6445, n_6310);
  fflopd g5694_reg(.CK (clock), .D (n_5484), .Q (g5694));
  fflopd g3694_reg(.CK (clock), .D (n_5428), .Q (g3694));
  nand g177165 (n_6782, g35, n_6015);
  nand g177164 (n_6775, g35, n_5661);
  nand g177161 (n_6760, g35, n_6014);
  nand g177160 (n_6756, g35, n_5662);
  nor g177154 (n_6503, n_4671, n_6013);
  nor g177152 (n_6501, n_4669, n_6012);
  fflopd g66_reg(.CK (clock), .D (n_5303), .Q (g18881));
  fflopd g6732_reg(.CK (clock), .D (n_5418), .Q (g6732));
  nand g177429 (n_6522, n_6011, n_5374);
  not g177221 (n_6533, n_6332);
  not g177216 (n_6547, n_6010);
  not g177215 (n_6542, n_6009);
  not g177222 (n_6528, n_6415);
  fflopd g209_reg(.CK (clock), .D (n_5294), .Q (g209));
  nand g177700 (n_6008, n_1253, n_5457);
  not g177552 (n_6007, n_5670);
  not g177554 (n_6005, n_5667);
  not g177556 (n_6004, n_5724);
  not g177557 (n_6003, n_5746);
  not g177558 (n_6002, n_5747);
  not g177559 (n_6001, n_5748);
  not g177560 (n_6000, n_5749);
  not g177561 (n_5999, n_5750);
  not g177562 (n_5998, n_5751);
  not g177563 (n_5997, n_5821);
  not g177564 (n_5996, n_5822);
  not g177565 (n_5995, n_5824);
  not g177566 (n_5994, n_5825);
  not g177567 (n_5993, n_5827);
  not g177568 (n_5992, n_5843);
  not g177569 (n_5991, n_5844);
  not g177570 (n_5990, n_5650);
  not g177571 (n_5989, n_5658);
  not g177572 (n_5988, n_5657);
  not g177573 (n_5987, n_5656);
  not g177574 (n_5986, n_5655);
  not g177577 (n_5984, n_5652);
  not g177579 (n_5983, n_5649);
  not g177581 (n_5982, n_5648);
  not g177582 (n_5981, n_5647);
  not g177583 (n_5980, n_5646);
  not g177584 (n_5979, n_5645);
  not g177585 (n_5978, n_5644);
  not g177586 (n_5977, n_5643);
  not g177587 (n_5976, n_5642);
  not g177588 (n_5975, n_5641);
  not g177589 (n_5974, n_5640);
  not g177590 (n_5973, n_5639);
  not g177591 (n_5972, n_5638);
  not g177592 (n_5971, n_5637);
  not g177593 (n_5970, n_5636);
  not g177594 (n_5969, n_5635);
  not g177595 (n_5968, n_5634);
  not g177596 (n_5967, n_5633);
  not g177597 (n_5966, n_5632);
  not g177598 (n_5965, n_5631);
  not g177601 (n_5963, n_5629);
  not g177606 (n_5962, n_5626);
  not g177607 (n_5961, n_5622);
  not g177608 (n_5960, n_5621);
  not g177609 (n_5959, n_5620);
  not g177610 (n_5958, n_5619);
  not g177611 (n_5957, n_5618);
  not g177612 (n_5956, n_5617);
  not g177613 (n_5955, n_5616);
  not g177614 (n_5954, n_5615);
  not g177615 (n_5953, n_5614);
  not g177616 (n_5952, n_5613);
  not g177617 (n_5951, n_5612);
  not g177618 (n_5950, n_5611);
  not g177619 (n_5949, n_5610);
  not g177620 (n_5948, n_5609);
  not g177621 (n_5947, n_5608);
  not g177622 (n_5946, n_5607);
  not g177623 (n_5945, n_5606);
  not g177624 (n_5944, n_5605);
  not g177627 (n_5942, n_5602);
  not g177629 (n_5941, n_5601);
  not g177632 (n_5940, n_5600);
  not g177633 (n_5939, n_5598);
  not g177636 (n_5938, n_5597);
  not g177637 (n_5937, n_5595);
  not g177649 (n_5936, n_5589);
  not g177650 (n_5935, n_5588);
  not g177651 (n_5934, n_5587);
  not g177652 (n_5933, n_5586);
  not g177653 (n_5932, n_5585);
  not g177654 (n_5931, n_5584);
  not g177655 (n_5930, n_5583);
  not g177656 (n_5929, n_5582);
  not g177657 (n_5928, n_5581);
  not g177658 (n_5927, n_5580);
  not g177659 (n_5926, n_5579);
  not g177660 (n_5925, n_5578);
  not g177661 (n_5924, n_5577);
  not g177662 (n_5923, n_5576);
  not g177663 (n_5922, n_5575);
  not g177664 (n_5921, n_5574);
  not g177665 (n_5920, n_5573);
  nand g178462 (n_5918, n_759, n_5326);
  wire w39, w40, w41, w42;
  nand g177681 (n_5917, w40, w42);
  nand g48 (w42, w41, g990);
  not g47 (w41, n_5916);
  nand g46 (w40, w39, n_5916);
  not g45 (w39, g990);
  nand g177689 (n_5915, g35, n_5307);
  not g177551 (n_5914, n_5671);
  nand g177720 (n_5913, g35, n_5304);
  nand g177723 (n_5912, n_2160, n_5458);
  nand g177744 (n_5911, g6513, n_5494);
  wire w43, w44, w45, w46;
  nand g177748 (n_5910, w44, w46);
  nand g52 (w46, w45, g4601);
  not g51 (w45, n_5504);
  nand g50 (w44, w43, n_5504);
  not g49 (w43, g4601);
  nand g177749 (n_5909, n_877, n_5437);
  nand g177757 (n_5908, g3119, n_5495);
  nand g178403 (n_5907, n_1049, n_5279);
  nand g177781 (n_5906, n_717, n_5460);
  nand g177785 (n_5905, g5475, n_5501);
  nand g177788 (n_5904, n_1032, n_5347);
  nand g177791 (n_5903, g3470, n_5499);
  nand g177813 (n_5902, n_2329, n_5375);
  nand g177818 (n_5901, n_797, n_5439);
  nand g177821 (n_5900, n_3703, n_5367);
  nand g177825 (n_5899, g3821, n_5496);
  nand g177848 (n_5898, n_1363, n_5461);
  nand g177850 (n_5897, n_4839, n_5440);
  nand g177860 (n_5896, n_4237, n_5345);
  nand g177863 (n_5895, g6167, n_5497);
  nand g177868 (n_5894, n_2068, n_5459);
  nand g177873 (n_5893, n_5305, n_4985);
  nand g177885 (n_5892, n_4790, n_5357);
  nand g177892 (n_5891, g35, n_5474);
  nand g177894 (n_5890, n_1029, n_5436);
  nand g177906 (n_5889, g5128, n_5500);
  nand g177920 (n_5888, n_5316, n_5560);
  nand g177926 (n_5887, n_2154, n_5489);
  nand g177929 (n_5886, n_1037, n_5455);
  nand g177931 (n_5885, n_4013, n_5883);
  nand g177933 (n_5884, n_4225, n_5883);
  nand g177934 (n_5882, n_4008, n_5883);
  nor g178879 (n_5881, n_5880, n_5878);
  nor g178638 (n_5879, n_3377, n_5878);
  nand g178609 (n_5877, g5052, n_5878);
  not g177965 (n_5875, n_5874);
  nand g178022 (n_5873, n_4723, n_5291);
  nand g178029 (n_5872, n_882, n_5284);
  nand g178061 (n_5871, n_5869, n_4625);
  nand g178062 (n_5870, n_5869, n_4534);
  nand g178074 (n_5867, g4709, n_5864);
  nand g177886 (g26877, n_5480, n_5328);
  nand g178099 (n_5865, n_4747, n_5864);
  nand g178106 (n_5863, n_964, n_5281);
  nand g178114 (n_5862, n_5293, n_4909);
  nand g178115 (n_5861, g4785, n_5864);
  nand g178116 (n_5860, n_5274, n_4916);
  nand g178496 (n_5859, n_9257, n_5848);
  nand g178349 (n_5858, g35, n_5341);
  not g178241 (n_5855, n_5505);
  not g178248 (n_5854, n_5541);
  not g178260 (n_5853, n_5841);
  not g178263 (n_5851, n_5518);
  nand g178196 (n_6474, n_3070, n_10186);
  not g177670 (n_6647, n_5563);
  fflopd g843_reg(.CK (clock), .D (n_5490), .Q (g843));
  nand g177949 (n_6185, g1996, n_6018);
  nand g177951 (n_6186, g35, n_6018);
  nand g177953 (n_6183, g35, n_5849);
  nand g178538 (n_6182, g35, n_5287);
  nor g178177 (n_6217, g168, n_5290);
  fflopd g5965_reg(.CK (clock), .D (n_5403), .Q (g5965));
  fflopd g5619_reg(.CK (clock), .D (n_5399), .Q (g5619));
  nand g178187 (n_6472, n_4672, n_5292);
  fflopd g3147_reg(.CK (clock), .D (n_5351), .Q (g3147));
  fflopd g3263_reg(.CK (clock), .D (n_5400), .Q (g3263));
  fflopd g3849_reg(.CK (clock), .D (n_5349), .Q (g3849));
  fflopd g3965_reg(.CK (clock), .D (n_5402), .Q (g3965));
  fflopd g5156_reg(.CK (clock), .D (n_5348), .Q (g5156));
  fflopd g3498_reg(.CK (clock), .D (n_5350), .Q (g3498));
  fflopd g5849_reg(.CK (clock), .D (n_5352), .Q (g5849));
  nand g178186 (n_6485, g2724, n_5848);
  fflopd g3614_reg(.CK (clock), .D (n_5401), .Q (g3614));
  fflopd g5272_reg(.CK (clock), .D (n_5398), .Q (g5272));
  fflopd g5503_reg(.CK (clock), .D (n_5353), .Q (g5503));
  nand g178547 (n_6468, n_5848, n_5503);
  nand g177954 (n_6516, g1728, n_5849);
  fflopd g411_reg(.CK (clock), .D (n_5395), .Q (g411));
  fflopd g822_reg(.CK (clock), .D (n_5419), .Q (g822));
  fflopd g1448_reg(.CK (clock), .D (n_5275), .Q (g1448));
  fflopd g1399_reg(.CK (clock), .D (n_5312), .Q (g19357));
  fflopd g3654_reg(.CK (clock), .D (n_5469), .Q (g11388));
  fflopd g6351_reg(.CK (clock), .D (n_5470), .Q (g12422));
  fflopd g6697_reg(.CK (clock), .D (n_5468), .Q (g12470));
  fflopd g5659_reg(.CK (clock), .D (n_5472), .Q (g12300));
  fflopd g6005_reg(.CK (clock), .D (n_5471), .Q (g12350));
  fflopd g703_reg(.CK (clock), .D (n_5385), .Q (g703));
  nand g178442 (n_5847, g4801, n_4884);
  nand g178475 (n_5845, n_4714, n_4915);
  nand g177774 (n_5844, n_3191, n_5070);
  nand g177773 (n_5843, n_3192, n_5147);
  nand g178424 (n_5842, n_4933, n_4717);
  nand g178453 (n_5841, n_853, n_4904);
  nand g178454 (n_5840, g35, n_4905);
  not g177193 (n_5839, n_5838);
  not g177194 (n_5837, n_5836);
  not g177195 (n_5835, n_5834);
  not g177196 (n_5833, n_5832);
  not g177200 (n_5831, n_5830);
  not g177201 (n_5829, n_5828);
  nand g177772 (n_5827, n_3193, n_4974);
  not g177205 (n_5826, g5073);
  nand g177771 (n_5825, n_3154, n_5144);
  nand g177770 (n_5824, n_3195, n_5068);
  not g177210 (n_5823, n_6013);
  nand g177769 (n_5822, n_3020, n_5121);
  nand g177768 (n_5821, n_3196, n_4964);
  nand g177767 (n_5820, g35, n_4977);
  nand g177224 (n_5819, n_3530, n_4961);
  nand g177225 (n_5818, n_3178, n_5165);
  nand g177227 (n_5817, n_3128, n_5028);
  nand g177228 (n_5816, g35, n_5113);
  nand g177230 (n_5815, n_3252, n_5041);
  nand g177231 (n_5814, n_924, n_5271);
  nand g177233 (n_5813, n_1337, n_4889);
  nand g177235 (n_5812, n_2903, n_5100);
  nand g177237 (n_5811, n_3215, n_5222);
  nand g177238 (n_5810, n_3221, n_5101);
  nand g177239 (n_5809, n_3117, n_5238);
  nand g177240 (n_5808, n_3158, n_5203);
  nand g177241 (n_5807, n_3097, n_5200);
  nand g177242 (n_5806, n_3225, n_5013);
  nand g177243 (n_5805, n_3204, n_5102);
  nand g177244 (n_5804, n_3262, n_5084);
  nand g177245 (n_5803, n_3226, n_4980);
  nand g177246 (n_5802, n_3100, n_5237);
  nand g177247 (n_5801, n_3573, n_5104);
  nand g177248 (n_5800, n_3579, n_5219);
  nand g177249 (n_5799, n_3156, n_5135);
  nand g177250 (n_5798, n_3580, n_5107);
  nand g177251 (n_5797, n_3545, n_4903);
  nand g177252 (n_5796, g14167, n_5795);
  nand g177268 (n_5794, g35, n_5176);
  nand g177274 (n_5793, n_528, n_5010);
  nand g177275 (n_5792, g4438, n_2040);
  nand g177279 (n_5791, n_6886, n_5062);
  nand g177280 (n_5790, n_5789, n_5063);
  nand g177281 (n_5788, n_6884, n_5066);
  nand g177282 (n_5787, n_6881, n_5058);
  nand g177283 (n_5786, n_6881, n_4902);
  nor g177284 (n_5785, g5808, n_5783);
  nor g177285 (n_5784, g5827, n_5783);
  nand g177286 (n_5782, n_5009, n_4065);
  nand g177287 (n_5781, n_5765, n_4198);
  nor g177289 (n_5780, g5481, n_5767);
  nor g177290 (n_5779, g6519, n_5770);
  nor g177295 (n_5778, g3106, n_5776);
  nor g177296 (n_5777, g3125, n_5776);
  nor g177300 (n_5775, g3808, n_5773);
  nor g177301 (n_5774, g3827, n_5773);
  nand g177308 (n_5772, n_5763, n_4206);
  nor g177310 (n_5771, g6500, n_5770);
  nand g177311 (n_5769, n_5289, n_5593);
  nor g177315 (n_5768, g5462, n_5767);
  nand g177327 (n_5766, n_5765, n_5248);
  nand g177328 (n_5764, n_5763, n_4950);
  nand g177367 (n_5762, n_5109, n_4159);
  nand g177369 (n_5761, n_5065, n_5760);
  nand g177370 (n_5759, n_5064, n_5758);
  nand g177376 (n_5757, n_5067, n_6450);
  nand g177377 (n_5756, n_5060, n_6456);
  nand g177378 (n_5755, n_5059, n_6454);
  nor g177384 (n_5754, g14421, n_5141);
  nor g177385 (n_5753, g14518, n_5140);
  nor g177386 (n_5752, g13039, n_5139);
  nand g177766 (n_5751, n_3150, n_4983);
  nand g177764 (n_5750, n_3558, n_5074);
  nand g177763 (n_5749, n_3559, n_5061);
  nand g177762 (n_5748, n_3369, n_5137);
  nand g177761 (n_5747, n_3560, n_5075);
  nand g177759 (n_5746, n_3561, n_4965);
  nand g177758 (n_5745, g35, n_4991);
  not g177578 (n_5744, n_5431);
  not g177580 (n_5743, n_5429);
  not g177603 (n_5742, n_5426);
  not g177605 (n_5741, n_5424);
  not g177635 (n_5740, n_5420);
  not g177639 (n_5739, n_5417);
  not g177641 (n_5737, n_5415);
  not g177642 (n_5736, n_5414);
  not g177643 (n_5735, n_5411);
  not g177647 (n_5733, n_5409);
  not g177669 (n_5732, n_5731);
  nand g177756 (n_5730, g35, n_5118);
  not g177672 (n_5729, n_6012);
  nand g177755 (n_5728, g1472, n_5726);
  nand g177753 (n_5727, g1448, n_5726);
  nand g177751 (n_5725, g1478, n_5726);
  nand g177750 (n_5724, n_3528, n_5026);
  nand g177682 (n_5723, n_3177, n_5138);
  nand g177683 (n_5722, n_3577, n_5223);
  nand g177684 (n_5721, n_3576, n_5093);
  nand g177685 (n_5720, n_3180, n_5004);
  nand g177686 (n_5719, n_3213, n_4968);
  nand g177687 (n_5718, n_3212, n_5092);
  nand g177688 (n_5717, n_3227, n_5224);
  nand g177690 (n_5716, n_3099, n_4881);
  nand g177691 (n_5715, n_3120, n_5090);
  nand g177692 (n_5714, n_3210, n_5226);
  nand g177693 (n_5713, n_3088, n_5088);
  nand g177695 (n_5712, n_3208, n_5087);
  nand g177696 (n_5711, n_3160, n_5245);
  nand g177697 (n_5710, n_3578, n_5095);
  nand g177698 (n_5709, n_2944, n_5198);
  nand g177699 (n_5708, n_3090, n_5025);
  nand g177701 (n_5707, n_2155, n_4992);
  nand g177703 (n_5706, n_695, n_5014);
  nand g177705 (n_5705, n_3544, n_5257);
  nand g177706 (n_5704, n_3540, n_5086);
  nand g177707 (n_5703, n_3205, n_5124);
  nand g177708 (n_5702, n_3575, n_5055);
  nand g177709 (n_5701, n_3214, n_5002);
  nand g177710 (n_5700, n_3203, n_4986);
  nand g177711 (n_5699, n_3201, n_5082);
  nand g177712 (n_5698, n_3200, n_5053);
  nand g177713 (n_5697, n_3199, n_5050);
  nand g177714 (n_5696, n_1290, n_5695);
  nand g177715 (n_5694, n_3220, n_5034);
  nand g177716 (n_5693, n_3113, n_5080);
  nand g177717 (n_5692, n_3236, n_5048);
  nand g177718 (n_5691, n_3171, n_5046);
  nand g177719 (n_5690, n_3239, n_4984);
  nand g177721 (n_5689, n_3115, n_5045);
  nand g177722 (n_5688, n_2939, n_5043);
  nand g177724 (n_5687, n_1116, n_4989);
  nand g177726 (n_5686, n_3574, n_5054);
  nand g177727 (n_5685, n_1196, n_4972);
  nand g177728 (n_5684, g35, n_5116);
  nand g177730 (n_5683, n_3542, n_5097);
  nand g177731 (n_5682, n_3251, n_5122);
  nand g177732 (n_5681, n_3572, n_5057);
  nand g177733 (n_5680, n_3543, n_5042);
  nand g177734 (n_5679, n_3253, n_4998);
  nand g177735 (n_5678, n_3125, n_5239);
  nand g177736 (n_5677, n_3261, n_5077);
  nand g177737 (n_5676, n_3254, n_5027);
  nand g177738 (n_5675, n_3248, n_5030);
  nand g177739 (n_5674, n_3258, n_4951);
  nand g177740 (n_5673, n_3259, n_5078);
  nand g177741 (n_5672, n_3134, n_5031);
  nand g177742 (n_5671, n_3086, n_5196);
  nand g177743 (n_5670, n_2902, n_5038);
  nand g177745 (n_5669, g35, n_5000);
  nand g177746 (n_5668, n_831, n_5241);
  nand g177747 (n_5667, n_845, n_4966);
  not g177677 (n_6307, n_5666);
  not g177675 (n_6313, n_5665);
  not g177673 (n_6308, n_5664);
  not g177671 (n_6306, n_5663);
  fflopd g3050_reg(.CK (clock), .D (n_4995), .Q (g3050));
  not g177204 (n_6368, n_5662);
  not g177208 (n_6378, n_5661);
  nand g177478 (n_6010, g35, n_5227);
  nand g177476 (n_6009, g35, n_5228);
  nor g177428 (n_6387, g4438, n_2285);
  fflopd g872_reg(.CK (clock), .D (g14167), .Q (g872));
  not g177214 (n_6424, n_6014);
  not g177212 (n_6422, n_6015);
  not g177680 (n_6339, n_6117);
  not g177217 (n_6342, n_6140);
  nand g177487 (n_6310, n_5660, n_5143);
  fflopd g239_reg(.CK (clock), .D (n_5177), .Q (g239));
  fflopd g4358_reg(.CK (clock), .D (n_5117), .Q (g4358));
  nand g177492 (n_6332, g35, n_5229);
  nand g177494 (n_6415, g35, n_5230);
  nand g178409 (n_5659, n_4927, n_4778);
  nand g177776 (n_5658, n_3189, n_4963);
  nand g177777 (n_5657, n_3188, n_5171);
  nand g177779 (n_5656, n_3187, n_5071);
  nand g177780 (n_5655, n_2973, n_5185);
  nand g177782 (n_5654, n_2151, n_4962);
  nand g177783 (n_5653, n_1000, n_5174);
  nand g177784 (n_5652, n_1252, n_4959);
  nand g177789 (n_5651, g35, n_5006);
  nand g177775 (n_5650, n_3190, n_5169);
  nand g177793 (n_5649, n_3247, n_5079);
  nand g177795 (n_5648, n_3555, n_4958);
  nand g177796 (n_5647, n_3554, n_5192);
  nand g177797 (n_5646, n_3176, n_5119);
  nand g177798 (n_5645, n_3629, n_5072);
  nand g177799 (n_5644, n_3552, n_5205);
  nand g177800 (n_5643, n_3386, n_5162);
  nand g177801 (n_5642, n_3175, n_4956);
  nand g177802 (n_5641, n_3172, n_5211);
  nand g177803 (n_5640, n_3385, n_5231);
  nand g177804 (n_5639, n_3170, n_5213);
  nand g177805 (n_5638, n_3169, n_4955);
  nand g177806 (n_5637, n_3166, n_5156);
  nand g177807 (n_5636, n_3384, n_5259);
  nand g177808 (n_5635, n_3163, n_5158);
  nand g177809 (n_5634, n_3162, n_4954);
  nand g177810 (n_5633, n_3161, n_5159);
  nand g177811 (n_5632, n_3383, n_5260);
  nand g177812 (n_5631, n_2914, n_5161);
  nand g177814 (n_5630, n_1385, n_4953);
  nand g177816 (n_5629, n_648, n_4949);
  wire w47, w48, w49, w50;
  nand g177819 (n_5628, w48, w50);
  nand g57 (w50, w49, g1472);
  not g56 (w49, n_5623);
  nand g54 (w48, w47, n_5623);
  not g53 (w47, g1472);
  nand g177824 (n_5627, g35, n_5115);
  nand g177826 (n_5626, n_3209, n_4979);
  nand g177828 (n_5625, g35, n_5235);
  wire w51, w52, w53, w54;
  nand g177829 (n_5624, w52, w54);
  nand g61 (w54, w53, g1448);
  not g60 (w53, n_5623);
  nand g59 (w52, w51, n_5623);
  not g58 (w51, g1448);
  nand g177830 (n_5622, n_3548, n_4948);
  nand g177831 (n_5621, n_3547, n_5166);
  nand g177832 (n_5620, n_3148, n_5136);
  nand g177833 (n_5619, n_3431, n_5265);
  nand g177834 (n_5618, n_3546, n_5179);
  nand g177835 (n_5617, n_3146, n_5249);
  nand g177836 (n_5616, n_3206, n_4982);
  nand g177837 (n_5615, n_3145, n_5180);
  nand g177838 (n_5614, n_3144, n_5266);
  nand g177839 (n_5613, n_3211, n_5182);
  nand g177840 (n_5612, n_3143, n_5269);
  nand g177841 (n_5611, n_3142, n_5184);
  nand g177842 (n_5610, n_3141, n_4940);
  nand g177843 (n_5609, n_3140, n_5188);
  nand g177844 (n_5608, n_3139, n_5256);
  nand g177845 (n_5607, n_3173, n_5189);
  nand g177846 (n_5606, n_3138, n_4987);
  nand g177847 (n_5605, n_2906, n_5194);
  nand g177849 (n_5604, n_2069, n_5252);
  nand g177851 (n_5603, n_934, n_5173);
  nand g177852 (n_5602, n_651, n_5246);
  nand g177856 (n_5601, n_3551, n_4967);
  nand g177864 (n_5600, g35, n_4976);
  nand g177866 (n_5599, g4438, n_2032);
  nand g177867 (n_5598, n_3270, n_5029);
  nand g177870 (n_5597, n_3126, n_5234);
  wire w55, w56, w57, w58;
  nand g177871 (n_5596, w56, w58);
  nand g65 (w58, w57, g1478);
  not g64 (w57, n_5623);
  nand g63 (w56, w55, n_5623);
  not g62 (w55, g1478);
  nand g177874 (n_5595, n_3127, n_5032);
  nand g177875 (n_5594, g283, n_5593);
  nand g177895 (n_5592, g35, n_5112);
  nand g177902 (n_5591, n_5149, n_4805);
  nand g177904 (n_5590, n_4617, n_5129);
  nand g177905 (n_5589, g35, n_5003);
  nand g177909 (n_5588, n_3536, n_5015);
  nand g177910 (n_5587, n_3529, n_5202);
  nand g177911 (n_5586, n_3216, n_5133);
  nand g177912 (n_5585, n_3527, n_5206);
  nand g177913 (n_5584, n_3102, n_5263);
  nand g177914 (n_5583, n_3096, n_5016);
  nand g177915 (n_5582, n_3095, n_5207);
  nand g177916 (n_5581, n_3149, n_5262);
  nand g177917 (n_5580, n_3093, n_5210);
  nand g177918 (n_5579, n_3092, n_5018);
  nand g177919 (n_5578, n_3091, n_5215);
  nand g177921 (n_5577, n_3224, n_5099);
  nand g177922 (n_5576, n_3089, n_4960);
  nand g177923 (n_5575, n_3119, n_5217);
  nand g177924 (n_5574, n_3108, n_5033);
  nand g177925 (n_5573, n_2905, n_5218);
  nand g177927 (n_5572, n_925, n_4923);
  nand g177928 (n_5571, n_1408, n_5167);
  nand g177930 (n_5570, g35, n_4994);
  nand g177935 (n_5569, n_4647, n_5125);
  nand g177937 (n_5568, n_4614, n_5142);
  nand g177938 (n_5567, n_5155, n_4797);
  nand g177941 (n_5566, n_4616, n_5131);
  nand g177942 (n_5565, n_5153, n_4804);
  nand g177943 (n_5564, n_5151, n_4622);
  nand g177945 (n_5563, n_5329, n_5324);
  not g177958 (n_5562, n_5369);
  not g177962 (n_5561, n_5560);
  not g177968 (n_5559, n_5849);
  not g177970 (n_5558, n_6018);
  nor g178014 (n_5557, n_5273, n_4400);
  nand g178063 (n_5556, n_1173, n_4937);
  nand g178090 (n_5555, n_640, n_4906);
  nand g178124 (n_5554, g5128, n_5552);
  nand g178125 (n_5553, n_178, n_5552);
  nand g178426 (n_5551, n_4867, n_4941);
  nand g178133 (n_5550, n_5549, n_4899);
  nand g178141 (n_5548, g6167, n_5546);
  nand g178142 (n_5547, n_159, n_5546);
  nand g178143 (n_5545, g3470, n_5543);
  nand g178144 (n_5544, n_234, n_5543);
  nand g178427 (n_5542, n_4934, n_4715);
  nand g178410 (n_5541, n_847, n_4928);
  not g178230 (n_5540, n_5309);
  not g178232 (n_5539, n_5308);
  not g178234 (n_5538, n_5306);
  not g178235 (n_5537, n_5302);
  not g178236 (n_5536, n_5301);
  not g178238 (n_5535, n_5298);
  not g178239 (n_5534, n_5376);
  not g178240 (n_5533, n_5283);
  not g178247 (n_5531, n_5485);
  not g178251 (n_5530, n_5483);
  not g178256 (n_5529, n_5295);
  not g178264 (n_5528, n_5297);
  not g178265 (n_5527, n_5473);
  not g178268 (n_5526, n_5525);
  nand g178463 (n_5524, g5037, n_4892);
  nand g178392 (n_5523, n_4379, n_4888);
  nand g178428 (n_5522, g4322, n_4944);
  nand g178465 (n_5521, n_5272, n_5520);
  nand g178466 (n_5519, n_3234, n_4894);
  nand g178464 (n_5518, n_1277, n_4898);
  nand g178676 (n_5517, n_569, n_4971);
  nand g178645 (n_5516, g5046, n_4975);
  nand g178412 (n_5515, n_4929, n_4722);
  nand g178292 (n_5514, n_4931, n_4718);
  nand g178396 (n_5513, n_5346, n_4886);
  nor g178335 (n_5512, n_9257, n_4924);
  nand g178340 (n_5511, n_9257, n_4936);
  nand g178343 (n_5510, g35, n_4901);
  nand g178350 (n_5509, n_3401, n_4900);
  nand g178351 (n_5508, g35, n_4908);
  nand g178413 (n_5507, n_4930, n_4721);
  nand g178365 (n_5506, n_4375, n_4885);
  nand g178395 (n_5505, n_4910, n_4887);
  fflopd g5752_reg(.CK (clock), .D (n_5008), .Q (g5752));
  fflopd g6098_reg(.CK (clock), .D (n_5242), .Q (g6098));
  fflopd g6444_reg(.CK (clock), .D (n_5001), .Q (g6444));
  fflopd g3752_reg(.CK (clock), .D (n_4947), .Q (g3752));
  fflopd g3401_reg(.CK (clock), .D (n_4981), .Q (g3401));
  fflopd g475_reg(.CK (clock), .D (n_4911), .Q (g475));
  fflopd g2898_reg(.CK (clock), .D (n_4913), .Q (g2898));
  nand g178194 (n_5874, g4601, n_5504);
  nand g178517 (n_6192, g35, n_4935);
  fflopd g5406_reg(.CK (clock), .D (n_4970), .Q (g5406));
  nand g178198 (n_6248, g2729, n_5503);
  fflopd g4382_reg(.CK (clock), .D (n_5108), .Q (g4382));
  not g178281 (n_7901, n_5502);
  fflopd g1389_reg(.CK (clock), .D (n_4997), .Q (g1389));
  fflopd g4669_reg(.CK (clock), .D (n_5254), .Q (g4669));
  fflopd g4408_reg(.CK (clock), .D (n_5172), .Q (g7243));
  nand g178535 (n_6271, g35, n_5546);
  nand g178526 (n_6250, g2729, g2724);
  nand g178532 (n_6274, g35, n_5543);
  nand g178536 (n_6268, g35, n_5552);
  not g178290 (n_6241, n_5501);
  not g178288 (n_6258, n_5500);
  not g178287 (n_6261, n_5499);
  fflopd g5029_reg(.CK (clock), .D (n_4891), .Q (g5029));
  not g178286 (n_6238, n_5498);
  not g178285 (n_6265, n_5497);
  not g178284 (n_6233, n_5496);
  not g178289 (n_6222, n_5495);
  not g178283 (n_6226, n_5494);
  fflopd g1472_reg(.CK (clock), .D (n_4925), .Q (g1472));
  fflopd g1478_reg(.CK (clock), .D (n_4926), .Q (g1478));
  fflopd g753_reg(.CK (clock), .D (n_4945), .Q (g753));
  fflopd g1041_reg(.CK (clock), .D (n_4907), .Q (g1041));
  fflopd g1404_reg(.CK (clock), .D (n_4996), .Q (g1404));
  fflopd g817_reg(.CK (clock), .D (n_4917), .Q (g817));
  fflopd g392_reg(.CK (clock), .D (n_4919), .Q (g392));
  nand g178066 (n_5493, n_1618, n_5492);
  nand g178443 (n_5491, n_4333, n_4796);
  nand g178441 (n_5490, n_4711, n_4706);
  nand g178064 (n_5489, g5297, n_5392);
  nand g178456 (n_5487, n_4815, n_3849);
  nand g178436 (n_5486, n_4329, n_4772);
  nand g178407 (n_5485, n_772, n_4738);
  nand g177232 (n_5484, n_1008, n_4849);
  nand g178422 (n_5483, n_633, n_4741);
  nand g177253 (n_5482, n_4854, n_4811);
  nor g177265 (n_5481, n_1792, n_5480);
  nor g177276 (n_5479, n_4800, n_2325);
  nor g177277 (n_5478, n_4858, n_2296);
  nor g177278 (n_5477, n_4699, n_2294);
  nor g177298 (n_5476, n_4818, n_1423);
  nand g177302 (n_5475, n_2854, n_4810);
  nand g178452 (n_5474, n_3712, n_4786);
  nand g178472 (n_5473, n_742, n_4744);
  nor g177360 (n_5472, g13049, n_4838);
  nor g177361 (n_5471, g13068, n_4837);
  nor g177362 (n_5470, g13085, n_4836);
  nor g177363 (n_5469, g14451, n_4835);
  nor g177364 (n_5468, g13099, n_4834);
  nor g177368 (n_5467, n_4803, n_5466);
  nor g177372 (n_5465, n_4857, n_5464);
  nor g177380 (n_5463, n_4862, n_5462);
  nand g178060 (n_5461, new_g10375_, n_5450);
  nand g178059 (n_5460, new_g10366_, n_5448);
  nand g178058 (n_5459, new_g10413_, n_5452);
  nand g178057 (n_5458, new_g10409_, n_5389);
  nand g178056 (n_5457, new_g10405_, n_5445);
  nand g178055 (n_5456, new_g10401_, n_5454);
  nand g178054 (n_5455, g5462, n_5454);
  nand g178053 (n_5453, g5011, n_5452);
  nand g178052 (n_5451, g4961, n_5450);
  nand g178051 (n_5449, g4939, n_5448);
  nand g178050 (n_5447, g4894, n_5452);
  nand g178049 (n_5446, g4831, n_5445);
  nand g178048 (n_5444, g4821, n_5454);
  nand g178047 (n_5443, g4760, n_5445);
  nand g178046 (n_5442, g4749, n_5454);
  nand g178045 (n_5441, g4035, n_5450);
  nand g178044 (n_5440, n_1076, n_10188);
  nand g178043 (n_5439, g3808, n_5450);
  nand g178042 (n_5438, g3333, n_5448);
  nand g178041 (n_5437, g3106, n_5448);
  nand g178040 (n_5436, g6500, n_5452);
  nand g177702 (n_5435, n_554, n_4848);
  nand g177725 (n_5434, n_1025, n_4847);
  nand g177752 (n_5433, g16686, g3247);
  nand g177754 (n_5432, g16686, g3255);
  nand g177786 (n_5431, g16722, g3598);
  nand g177787 (n_5430, g16722, g3606);
  nand g177794 (n_5429, g17715, g5957);
  nand g177815 (n_5428, n_521, n_4845);
  wire w59, w60, w61, w62;
  nand g177817 (n_5427, w60, w62);
  nand g69 (w62, w61, g1300);
  not g68 (w61, n_5036);
  nand g67 (w60, w59, n_5036);
  not g66 (w59, g1300);
  nand g177820 (n_5426, g16748, g3949);
  nand g177822 (n_5425, n_4417, n_4840);
  nand g177823 (n_5424, g16748, g3957);
  nand g177853 (n_5423, g17639, g5264);
  nand g177857 (n_5422, n_593, n_4844);
  nand g177865 (n_5421, g4401, n_4264);
  nand g177869 (n_5420, g17639, g5256);
  nand g177877 (n_5419, n_1267, n_4855);
  nand g177879 (n_5418, n_1332, n_4846);
  nand g177881 (n_5417, g17678, g5603);
  nand g177882 (n_5416, n_3714, n_4763);
  nand g177884 (n_5415, g17678, g5611);
  nand g177887 (n_5414, g17743, g6295);
  nand g177888 (n_5413, g17743, g6303);
  nor g177889 (n_5412, n_4850, n_4447);
  nand g177890 (n_5411, g17715, g5949);
  nand g177891 (n_5410, n_3724, n_4856);
  nand g177897 (n_5409, g17764, g6641);
  nand g177898 (n_5408, g17764, g6649);
  nor g177932 (n_5407, n_4843, n_4443);
  nor g177936 (n_5406, n_4841, n_3873);
  nor g177939 (n_5405, n_4833, n_4446);
  nand g178039 (n_5404, g5808, n_5445);
  nand g178036 (n_5403, n_4745, n_4196);
  nand g178035 (n_5402, n_4742, n_4197);
  nand g178034 (n_5401, n_4740, n_4200);
  nand g178033 (n_5400, n_4736, n_4203);
  nand g178032 (n_5399, n_4729, n_4211);
  nand g178031 (n_5398, n_4739, n_4202);
  not g177960 (n_5397, n_5111);
  nand g178007 (n_5396, n_107, n_4725);
  nand g178008 (n_5395, n_3841, n_4758);
  nand g178010 (n_5394, g3684, n_5386);
  nand g178012 (n_5393, g21245, n_5392);
  nand g178018 (n_5391, g4704, n_5392);
  nand g178019 (n_5390, g4771, n_5389);
  nand g178020 (n_5388, g4826, n_5389);
  nand g178021 (n_5387, g4950, n_5386);
  nand g178028 (n_5385, n_4377, n_4866);
  fflopd g4888_reg(.CK (clock), .D (n_4709), .Q (g4888));
  nand g177948 (n_5664, g2555, n_5384);
  nand g177946 (n_5663, g35, n_5384);
  nand g177944 (n_5731, g703, n_4830);
  nand g177453 (n_5661, n_5383, n_5384);
  nand g177952 (n_5666, g35, n_5382);
  nand g177430 (n_5662, n_5381, n_5382);
  nand g177417 (n_5828, n_1006, n_5384);
  nand g177416 (n_5830, n_1511, n_5384);
  nand g177412 (n_5832, n_5380, n_5384);
  nand g177411 (n_5834, n_1493, n_5382);
  nand g177410 (n_5836, n_5379, n_5382);
  nand g177409 (n_5838, n_565, n_5382);
  nand g177950 (n_5665, g2287, n_5382);
  nand g177947 (n_6012, g35, n_5378);
  fflopd g5685_reg(.CK (clock), .D (g17678), .Q (g5685));
  fflopd g6377_reg(.CK (clock), .D (g17743), .Q (g6377));
  fflopd g6031_reg(.CK (clock), .D (g17715), .Q (g6031));
  fflopd g6723_reg(.CK (clock), .D (g17764), .Q (g6723));
  fflopd g5073_reg(.CK (clock), .D (n_4827), .Q (g5073));
  nand g177480 (n_6140, g2421, n_5377);
  nand g177473 (n_6014, n_1461, n_5378);
  nand g177469 (n_6015, n_1606, n_5377);
  fflopd g4031_reg(.CK (clock), .D (g16748), .Q (g4031));
  nand g177462 (n_6013, g35, n_5377);
  fflopd g5339_reg(.CK (clock), .D (g17639), .Q (g5339));
  fflopd g3680_reg(.CK (clock), .D (g16722), .Q (g3680));
  fflopd g3329_reg(.CK (clock), .D (g16686), .Q (g3329));
  nand g177955 (n_6117, g2153, n_5378);
  fflopd g3119_reg(.CK (clock), .D (n_4694), .Q (g3119));
  nand g178390 (n_5376, n_1135, n_4733);
  nand g178070 (n_5375, new_g10371_, n_5386);
  nand g178071 (n_5374, n_1825, n_5492);
  nand g178073 (n_5373, n_11, n_5492);
  nand g178080 (n_5372, n_3237, n_7889);
  nand g178081 (n_5371, n_6890, n_7889);
  nand g178082 (n_5370, n_7535, n_7889);
  nand g178089 (n_5369, n_5368, n_4773);
  nand g178415 (n_5367, n_1563, n_4775);
  nand g178091 (n_5366, new_g7051_, n_5445);
  nand g178092 (n_5365, new_g7097_, n_5452);
  nand g178093 (n_5364, new_g7028_, n_5454);
  nand g178094 (n_5363, new_g6875_, n_5448);
  nand g178095 (n_5362, new_g6905_, n_5386);
  nand g178097 (n_5361, new_g6928_, n_5450);
  nand g178098 (n_5360, g4322, n_4869);
  nand g178100 (n_5359, new_g7004_, n_5392);
  nand g178101 (n_5358, new_g7074_, n_5389);
  nand g178105 (n_5357, n_1562, n_4768);
  nor g178108 (n_5356, n_2606, n_4719);
  nor g178113 (n_5355, n_2611, n_4713);
  nand g178118 (n_5354, n_1430, n_4821);
  nand g178127 (n_5353, n_4788, n_4354);
  nand g178128 (n_5352, n_4789, n_4355);
  nand g178129 (n_5351, n_4767, n_4356);
  nand g178130 (n_5350, n_4752, n_4357);
  nand g178131 (n_5349, n_4751, n_4359);
  nand g178132 (n_5348, n_4750, n_4361);
  nand g178401 (n_5347, n_5346, n_4732);
  nand g178151 (n_5345, n_3691, n_4783);
  nand g178067 (n_5344, n_87, n_5492);
  nand g178476 (n_5343, n_2716, n_4781);
  nand g178896 (n_5342, g35, n_4766);
  nor g178883 (n_5341, n_5340, n_5286);
  not g178228 (n_5338, n_5022);
  not g178253 (n_5333, n_5268);
  not g178254 (n_5332, n_5236);
  not g178255 (n_5331, n_5247);
  not g178269 (n_5328, n_5327);
  nand g178881 (n_5326, n_2649, n_4760);
  not g178272 (n_5323, n_5695);
  nand g178327 (n_5317, n_3903, n_5300);
  nand g178330 (n_5316, n_3969, n_5313);
  wire w63, w64, w65, w66;
  nand g178331 (n_5315, w64, w66);
  nand g73 (w66, w65, g739);
  not g72 (w65, n_4882);
  nand g71 (w64, w63, n_4882);
  not g70 (w63, g739);
  nor g178332 (n_5314, n_9257, n_5313);
  wire w67, w68, w69, w70;
  nand g178333 (n_5312, w68, w70);
  nand g77 (w70, w69, g1333);
  not g76 (w69, n_4920);
  nand g75 (w68, w67, n_4920);
  not g74 (w67, g1333);
  nand g178843 (n_5311, g20763, n_5310);
  nand g178357 (n_5309, n_921, n_4728);
  nand g178361 (n_5308, n_598, n_4743);
  nand g178363 (n_5307, n_2544, n_5313);
  nand g178368 (n_5306, n_639, n_4731);
  nand g178370 (n_5305, g812, n_4712);
  nand g178371 (n_5304, n_3131, n_4785);
  nand g178374 (n_5303, n_1200, n_4819);
  nand g178375 (n_5302, n_615, n_4730);
  nand g178380 (n_5301, n_3506, n_5300);
  nand g178382 (n_5299, n_4817, n_3707);
  nand g178386 (n_5298, n_4734, n_4624);
  nand g178468 (n_5297, n_753, n_4724);
  nand g178400 (n_5296, n_4436, n_4770);
  nand g178440 (n_5295, n_4707, n_4769);
  nand g178478 (n_5294, n_1342, n_4727);
  not g178787 (n_5293, n_4946);
  not g178779 (n_5292, n_4883);
  not g178775 (n_5291, n_4893);
  nand g178673 (n_5290, n_1934, n_5289);
  nand g178667 (n_5287, new_g10383_, n_5286);
  nand g178660 (n_5285, g2375, n_4762);
  nand g178654 (n_5284, n_2719, n_5280);
  nand g178391 (n_5283, n_857, n_4735);
  nand g178621 (n_5281, n_486, n_5280);
  nand g178586 (n_5279, g542, n_8904);
  nand g178585 (n_5278, g554, n_8904);
  nand g178581 (n_5277, n_5276, n_5289);
  nand g178575 (n_5275, n_4583, n_4757);
  not g178551 (n_5274, n_4918);
  nand g178542 (n_5498, g35, n_4793);
  nand g178543 (n_5499, g35, n_4873);
  nand g178544 (n_5500, g35, n_4874);
  nand g178545 (n_5495, g35, n_4791);
  nand g178546 (n_5501, g35, n_4792);
  nand g178539 (n_5494, g35, n_4795);
  fflopd g433_reg(.CK (clock), .D (n_4823), .Q (g433));
  nand g178537 (n_5502, g35, n_5492);
  not g178270 (n_6061, n_4943);
  nand g178521 (n_5525, g35, g4072);
  nand g178541 (n_5497, g35, n_4875);
  nand g178540 (n_5496, g35, n_4794);
  fflopd g4698_reg(.CK (clock), .D (n_4710), .Q (g4698));
  nand g178178 (n_5560, n_4073, n_5313);
  fflopd g460_reg(.CK (clock), .D (n_4779), .Q (g460));
  not g178795 (n_5869, n_5273);
  nor g178964 (n_5864, n_9257, n_5280);
  fflopd g832_reg(.CK (clock), .D (n_4807), .Q (g832));
  fflopd g1216_reg(.CK (clock), .D (n_4700), .Q (g1216));
  nor g178191 (n_5883, n_5035, n_5623);
  fflopd g699_reg(.CK (clock), .D (n_4865), .Q (g699));
  not g179043 (n_5878, n_5272);
  nand g178533 (n_6752, g35, n_7889);
  not g178560 (n_5848, g2729);
  fflopd g6167_reg(.CK (clock), .D (n_4753), .Q (g6167));
  fflopd g6513_reg(.CK (clock), .D (n_4701), .Q (g6513));
  fflopd g1559_reg(.CK (clock), .D (n_10375), .Q (g1559));
  fflopd g3821_reg(.CK (clock), .D (n_4704), .Q (g3821));
  fflopd g5128_reg(.CK (clock), .D (n_4754), .Q (g5128));
  nand g178210 (n_5849, n_3988, n_4780);
  fflopd g3470_reg(.CK (clock), .D (n_4703), .Q (g3470));
  fflopd g5475_reg(.CK (clock), .D (n_4755), .Q (g5475));
  fflopd g182_reg(.CK (clock), .D (n_4726), .Q (g182));
  fflopd g4349_reg(.CK (clock), .D (n_4765), .Q (g4349));
  nand g178219 (n_6018, n_4000, n_4784);
  fflopd g4793_reg(.CK (clock), .D (n_4705), .Q (g4793));
  nand g178483 (n_5271, n_459, n_5270);
  nand g178461 (n_5269, n_5186, n_5255);
  nand g178431 (n_5268, n_512, n_5267);
  nand g178315 (n_5266, n_5181, n_5264);
  nand g178314 (n_5265, n_5178, n_5264);
  nand g178459 (n_5263, new_g7704_, n_5261);
  nand g178313 (n_5262, n_5208, n_5261);
  nand g178312 (n_5260, n_5160, n_5258);
  nand g178311 (n_5259, n_5157, n_5258);
  nand g178490 (n_5257, n_5085, n_5123);
  nand g178457 (n_5256, n_5193, n_5255);
  nand g178439 (n_5254, n_3752, n_4590);
  nand g177010 (n_5253, g35, n_4658);
  nand g178455 (n_5252, n_5250, n_5251);
  nand g178423 (n_5249, new_g7121_, n_5264);
  nor g178489 (n_5248, n_4613, n_4173);
  nand g178438 (n_5247, n_714, n_4645);
  nand g178437 (n_5246, n_908, n_5251);
  nand g178420 (n_5245, n_5197, n_5225);
  nand g178405 (n_5242, n_3350, n_4621);
  nand g178421 (n_5241, n_5126, n_5240);
  nand g178435 (n_5239, n_5076, n_5233);
  nand g178481 (n_5238, n_5220, n_5134);
  nand g178471 (n_5237, new_g7738_, n_5221);
  nand g178433 (n_5236, n_4619, n_2144);
  nand g178419 (n_5235, g3821, n_5114);
  nand g178432 (n_5234, n_5195, n_5233);
  nand g178310 (n_5231, n_5212, n_5258);
  not g177966 (n_5230, n_5378);
  not g177967 (n_5229, n_5377);
  not g177969 (n_5228, n_5382);
  not g177971 (n_5227, n_5384);
  nand g177973 (n_5226, n_5089, n_5225);
  nand g177974 (n_5224, n_5163, n_5225);
  nand g177975 (n_5223, n_5094, n_5225);
  nand g177976 (n_5222, n_5220, n_5221);
  nand g177977 (n_5219, n_5105, n_5221);
  nand g177978 (n_5218, n_5216, n_5209);
  nand g177979 (n_5217, n_5216, n_5214);
  nand g177980 (n_5215, n_5098, n_5214);
  nand g177981 (n_5213, n_5212, n_5204);
  nand g177982 (n_5211, n_5212, n_5191);
  nand g177983 (n_5210, n_5208, n_5209);
  nand g177984 (n_5207, n_5208, n_5214);
  nand g177985 (n_5206, n_5201, n_5209);
  nand g177986 (n_5205, n_5190, n_5204);
  nand g177987 (n_5203, n_5199, n_5103);
  nand g177988 (n_5202, n_5201, n_5214);
  nand g177989 (n_5200, n_5199, n_5106);
  nand g177990 (n_5198, n_5197, n_5164);
  nand g177991 (n_5196, n_5195, n_5096);
  nand g177992 (n_5194, n_5193, n_5187);
  nand g177993 (n_5192, n_5190, n_5191);
  nand g177994 (n_5189, n_5193, n_5183);
  nand g177995 (n_5188, n_5186, n_5187);
  nand g177996 (n_5185, n_5170, n_5168);
  nand g177997 (n_5184, n_5186, n_5183);
  nand g177998 (n_5182, n_5181, n_5187);
  nand g177999 (n_5180, n_5181, n_5183);
  nand g178000 (n_5179, n_5178, n_5187);
  nand g178001 (n_5177, n_4663, n_4067);
  nor g178004 (n_5176, n_4138, n_5175);
  nand g178009 (n_5174, n_2079, n_4676);
  nand g178013 (n_5173, n_2103, n_4688);
  nand g178016 (n_5172, n_2748, n_4605);
  nand g178017 (n_5171, n_5170, n_5146);
  nand g178023 (n_5169, n_5145, n_5168);
  nand g178024 (n_5167, n_2081, n_4660);
  nand g178025 (n_5166, n_5178, n_5183);
  nand g178026 (n_5165, n_5163, n_5164);
  nand g178408 (n_5162, new_g10323_, n_5258);
  nand g178027 (n_5161, n_5160, n_5204);
  nand g178030 (n_5159, n_5160, n_5191);
  nand g178037 (n_5158, n_5157, n_5204);
  nand g178038 (n_5156, n_5157, n_5191);
  nand g178072 (n_5155, n_4606, n_5154);
  nand g178075 (n_5153, n_4611, n_5152);
  nand g178076 (n_5151, n_4599, n_5150);
  nand g178077 (n_5149, n_4603, n_5148);
  nand g178078 (n_5147, n_5145, n_5146);
  nand g178079 (n_5144, n_5120, n_5168);
  nor g178088 (n_5143, g1135, g27831);
  nand g178096 (n_5142, n_4608, n_5250);
  nand g178102 (n_5141, n_3858, n_4632);
  nand g178103 (n_5140, n_3795, n_4630);
  nand g178104 (n_5139, n_3352, n_4628);
  nand g178107 (n_5138, new_g7766_, n_4978);
  nand g178109 (n_5137, new_g10295_, n_4973);
  nand g178110 (n_5136, new_g7121_, n_5255);
  nand g178112 (n_5135, new_g7738_, n_5134);
  nand g178117 (n_5133, new_g7704_, n_5017);
  nand g178120 (n_5132, n_4604, n_4922);
  nand g178121 (n_5131, n_4601, n_5130);
  nand g178122 (n_5129, n_4602, n_5128);
  nand g178123 (n_5127, n_4609, n_5126);
  nand g178126 (n_5125, n_4610, n_4952);
  nand g178134 (n_5124, new_g7791_, n_5123);
  nand g178137 (n_5122, new_g7812_, n_5233);
  nand g178138 (n_5121, n_5120, n_5146);
  nand g178139 (n_5119, new_g10323_, n_4957);
  nand g178140 (n_5118, n_67, n_4990);
  nand g178429 (n_5117, n_1921, n_4588);
  nand g178145 (n_5116, n_164, n_4999);
  nand g178146 (n_5115, n_172, n_5114);
  nand g178147 (n_5113, n_141, n_5005);
  nand g178148 (n_5112, n_127, n_4993);
  nand g178149 (n_5111, n_2872, n_5110);
  nand g178150 (n_5109, g6381, n_4600);
  nand g178152 (n_5108, n_4109, n_10192);
  nand g178153 (n_5107, n_5105, n_5106);
  nand g178154 (n_5104, n_5105, n_5103);
  nand g178155 (n_5102, n_5083, n_5103);
  nand g178156 (n_5101, n_5220, n_5106);
  nand g178157 (n_5100, n_5220, n_5103);
  nand g178158 (n_5099, n_5098, n_5209);
  nand g178159 (n_5097, n_5056, n_5096);
  nand g178160 (n_5095, n_5094, n_5091);
  nand g178161 (n_5093, n_5094, n_5164);
  nand g178162 (n_5092, n_5163, n_5091);
  nand g178163 (n_5090, n_5089, n_5091);
  nand g178164 (n_5088, n_5089, n_5164);
  nand g178165 (n_5087, n_5197, n_5091);
  nand g178166 (n_5086, n_5085, n_5081);
  nand g178167 (n_5084, n_5083, n_5106);
  nand g178168 (n_5082, n_5051, n_5081);
  nand g178169 (n_5080, n_5047, n_5081);
  nand g178170 (n_5079, n_5044, n_5081);
  nand g178171 (n_5078, n_5039, n_5096);
  nand g178172 (n_5077, n_5076, n_5096);
  nand g178173 (n_5075, n_5073, n_5146);
  nand g178174 (n_5074, n_5073, n_5168);
  nand g178309 (n_5072, n_5190, n_5258);
  nand g178308 (n_5071, n_5170, n_5069);
  nand g178307 (n_5070, n_5145, n_5069);
  nand g178306 (n_5068, n_5120, n_5069);
  not g178233 (n_5067, n_4806);
  not g178237 (n_5066, n_4802);
  not g178242 (n_5065, n_4851);
  not g178249 (n_5064, n_4829);
  not g178250 (n_5063, n_4853);
  not g178252 (n_5062, n_4863);
  nand g178305 (n_5061, n_5073, n_5069);
  not g178257 (n_5060, n_4799);
  not g178258 (n_5059, n_4864);
  not g178259 (n_5058, n_4860);
  nand g178293 (n_5057, n_5056, n_5040);
  nand g178294 (n_5055, n_5085, n_5052);
  nand g178295 (n_5054, n_5085, n_5049);
  nand g178296 (n_5053, n_5051, n_5052);
  nand g178297 (n_5050, n_5051, n_5049);
  nand g178298 (n_5048, n_5047, n_5052);
  nand g178299 (n_5046, n_5047, n_5049);
  nand g178300 (n_5045, n_5044, n_5052);
  nand g178301 (n_5043, n_5044, n_5049);
  nand g178302 (n_5042, n_5056, n_5037);
  nand g178303 (n_5041, n_5039, n_5040);
  nand g178304 (n_5038, n_5195, n_5037);
  fflopd g4933_reg(.CK (clock), .D (n_4684), .Q (g4933));
  fflopd g4955_reg(.CK (clock), .D (n_4687), .Q (g4955));
  fflopd g6537_reg(.CK (clock), .D (n_4549), .Q (g6537));
  fflopd g3143_reg(.CK (clock), .D (n_4552), .Q (g3143));
  nand g178179 (n_5593, n_4395, n_10190);
  fflopd g6191_reg(.CK (clock), .D (n_4562), .Q (g6191));
  fflopd g4754_reg(.CK (clock), .D (n_4679), .Q (g4754));
  fflopd g4765_reg(.CK (clock), .D (n_4680), .Q (g4765));
  nor g178190 (n_5726, n_5035, n_5036);
  fflopd g4438_reg(.CK (clock), .D (n_4598), .Q (g4438));
  fflopd g887_reg(.CK (clock), .D (g14147), .Q (g14167));
  fflopd g1300_reg(.CK (clock), .D (n_4548), .Q (g1300));
  nand g178492 (n_5034, n_5047, n_5123);
  nand g178318 (n_5033, n_5216, n_5261);
  nand g178319 (n_5032, n_5199, n_5221);
  nand g178320 (n_5031, n_5039, n_5037);
  nand g178321 (n_5030, n_5076, n_5037);
  nand g178322 (n_5029, n_5195, n_5040);
  nand g178323 (n_5028, n_5083, n_5221);
  nand g178324 (n_5027, n_5076, n_5040);
  nand g178325 (n_5026, n_5201, n_5261);
  nand g178326 (n_5025, n_5098, n_5261);
  nand g178329 (n_5022, n_2819, n_5251);
  wire w71, w72, w73, w74;
  nand g178334 (n_5021, w72, w74);
  nand g81 (w74, w73, n_13);
  not g80 (w73, n_5276);
  nand g79 (w72, w71, n_5276);
  not g78 (w71, n_13);
  nand g178341 (n_5020, g35, n_4607);
  nand g178342 (n_5019, g35, n_4626);
  nand g178345 (n_5018, n_5098, n_5017);
  nand g178346 (n_5016, n_5208, n_5017);
  nand g178347 (n_5015, n_5201, n_5017);
  nand g178488 (n_5014, n_478, n_5023);
  nand g178352 (n_5013, n_5199, n_5134);
  nand g178354 (n_5010, n_902, n_5243);
  nand g178356 (n_5009, g14147, n_5795);
  nand g178358 (n_5008, n_3346, n_4620);
  nand g178360 (n_5006, g5821, n_5005);
  nand g178362 (n_5004, new_g7766_, n_5225);
  nand g178364 (n_5003, n_4181, n_4638);
  nand g178369 (n_5002, new_g7791_, n_5052);
  nand g178372 (n_5001, n_3235, n_4649);
  nand g178373 (n_5000, g6513, n_4999);
  nand g178376 (n_4998, new_g7812_, n_5040);
  nand g178377 (n_4997, n_4188, n_4666);
  nand g178378 (n_4996, n_4420, n_4674);
  nand g178381 (n_4995, n_3348, n_4650);
  nand g178384 (n_4994, g5475, n_4993);
  nand g178387 (n_4992, n_5128, n_5023);
  nand g178388 (n_4991, g3119, n_4990);
  nand g178494 (n_4989, n_4988, n_5110);
  nand g178317 (n_4987, n_5193, n_5264);
  nand g178491 (n_4986, n_5051, n_5123);
  nand g178389 (n_4985, g843, n_4665);
  nand g178493 (n_4984, n_5044, n_5123);
  nand g178393 (n_4983, new_g10295_, n_5069);
  nand g178469 (n_4982, n_5181, n_5255);
  nand g178397 (n_4981, n_3349, n_4651);
  nand g178402 (n_4980, n_5083, n_5134);
  nand g178487 (n_4979, n_5197, n_4978);
  nand g178394 (n_4977, n_5346, n_4612);
  nand g178430 (n_4976, n_2620, n_5267);
  not g179266 (n_4975, n_4872);
  nand g178501 (n_4974, n_5145, n_4973);
  nand g178495 (n_4972, n_822, n_5110);
  nand g179077 (n_4971, n_225, n_4877);
  nand g178477 (n_4970, n_3233, n_4661);
  not g179020 (n_4969, n_4698);
  nand g178484 (n_4968, n_5163, n_4978);
  nand g178497 (n_4967, n_5056, n_5233);
  nand g178498 (n_4966, n_904, n_5240);
  nand g178499 (n_4965, n_5073, n_4973);
  nand g178500 (n_4964, n_5120, n_4973);
  nand g178502 (n_4963, n_5170, n_4973);
  nand g178503 (n_4962, n_4168, n_5011);
  nand g178485 (n_4961, n_5094, n_4978);
  nand g178504 (n_4960, n_5216, n_5017);
  nand g178505 (n_4959, n_901, n_5011);
  nand g178506 (n_4958, n_5190, n_4957);
  nand g178507 (n_4956, n_5212, n_4957);
  nand g178508 (n_4955, n_5157, n_4957);
  nand g178509 (n_4954, n_5160, n_4957);
  nand g178510 (n_4953, n_4952, n_8166);
  nand g178511 (n_4951, n_5039, n_5233);
  nor g178512 (n_4950, n_4596, n_4175);
  nand g178513 (n_4949, n_482, n_8166);
  nand g178515 (n_4948, n_5178, n_5255);
  nand g178411 (n_4947, n_3181, n_4652);
  nand g178939 (n_4946, n_663, n_4582);
  nand g178933 (n_4945, n_4496, n_4561);
  nand g178931 (n_4944, g35, n_4683);
  nand g178524 (n_4943, n_4129, n_10192);
  nand g178926 (n_4941, new_g6946_, n_4302);
  nand g178316 (n_4940, n_5186, n_5264);
  not g178552 (n_4937, n_4820);
  not g178553 (n_4936, g4072);
  not g178554 (n_4935, n_5300);
  nand g178566 (n_4934, g728, n_4932);
  nand g178567 (n_4933, g718, n_4932);
  nand g178568 (n_4931, g681, n_4932);
  nand g178569 (n_4930, g661, n_4932);
  nand g178570 (n_4929, g655, n_4932);
  nand g178571 (n_4928, g650, n_4932);
  nand g178572 (n_4927, g645, n_4932);
  nand g178573 (n_4926, n_4312, n_4573);
  nand g178574 (n_4925, n_4311, n_4572);
  nand g178587 (n_4924, n_4541, n_2478);
  nand g178480 (n_4923, n_4922, n_5243);
  nand g178605 (n_4921, n_10400, n_4920);
  nand g178606 (n_4919, n_4309, n_4543);
  nand g178607 (n_4918, n_732, n_4544);
  nand g178612 (n_4917, n_3697, n_4577);
  nand g178614 (n_4916, g4975, n_4914);
  nand g178617 (n_4915, g4966, n_4914);
  nand g178619 (n_4913, n_2177, n_4912);
  nand g178623 (n_4911, n_3735, n_4574);
  nand g178624 (n_4910, n_3881, n_4685);
  nand g178631 (n_4909, g4584, n_4578);
  nor g178646 (n_4908, g9497, n_4530);
  nand g178647 (n_4907, n_4569, n_4337);
  nand g178648 (n_4906, n_4127, n_4914);
  nand g178658 (n_4905, n_2506, n_4565);
  nand g178672 (n_4904, g4899, n_4914);
  nand g178479 (n_4903, n_5105, n_5134);
  nand g178446 (n_4902, n_4644, n_3282);
  not g178784 (n_4901, n_4716);
  not g178788 (n_4900, n_4708);
  not g178796 (n_4899, n_5520);
  nand g178819 (n_4898, n_4594, n_4567);
  nand g178858 (n_4897, g35, n_4571);
  nand g178868 (n_4895, g35, n_4576);
  nand g178870 (n_4894, g35, n_4563);
  nand g178877 (n_4893, n_2709, n_4585);
  nand g178878 (n_4892, n_4579, n_4759);
  nand g178880 (n_4891, n_3656, n_4586);
  nand g178892 (n_4890, g355, n_4693);
  nand g178482 (n_4889, n_5130, n_5270);
  nand g178900 (n_4888, g1536, n_4553);
  nand g178901 (n_4887, n_2815, n_4554);
  nand g178902 (n_4886, g490, n_4696);
  nand g178904 (n_4885, g1193, n_4547);
  nand g178908 (n_4884, g35, n_4581);
  nand g178910 (n_4883, g739, n_4882);
  nand g178486 (n_4881, n_5089, n_4978);
  fflopd g5499_reg(.CK (clock), .D (n_4545), .Q (g5499));
  nand g178525 (n_5324, g35, n_4635);
  nand g178523 (n_5327, g35, n_4636);
  nand g178522 (n_5765, new_g7791_, n_5049);
  nand g178519 (n_5329, g35, n_4633);
  nand g178518 (n_5763, new_g7812_, n_5037);
  nand g178962 (n_5273, g35, new_g6946_);
  nor g178966 (n_5916, n_9257, n_4880);
  not g179277 (n_6427, n_4879);
  nor g178722 (n_5504, n_5340, n_4878);
  fflopd g4944_reg(.CK (clock), .D (n_4686), .Q (g4944));
  fflopd g3845_reg(.CK (clock), .D (n_4559), .Q (g3845));
  fflopd g3494_reg(.CK (clock), .D (n_4558), .Q (g3494));
  fflopd g5845_reg(.CK (clock), .D (n_4546), .Q (g5845));
  fflopd g4743_reg(.CK (clock), .D (n_4681), .Q (g4743));
  fflopd g5152_reg(.CK (clock), .D (n_4550), .Q (g5152));
  nand g179222 (n_5272, g5046, n_4877);
  fflopd g2886_reg(.CK (clock), .D (n_4667), .Q (g2886));
  not g179285 (n_6429, n_4876);
  fflopd g1233_reg(.CK (clock), .D (n_4655), .Q (g10500));
  fflopd g2729_reg(.CK (clock), .D (n_4584), .Q (g2729));
  nand g178531 (n_5783, g35, n_5005);
  nand g178534 (n_5773, g35, n_5114);
  nand g178530 (n_5767, g35, n_4993);
  not g178797 (n_5546, n_4875);
  fflopd g504_reg(.CK (clock), .D (n_4555), .Q (g504));
  not g178798 (n_5552, n_4874);
  not g178799 (n_5543, n_4873);
  nand g178527 (n_5695, g35, n_5175);
  nand g178528 (n_5776, g35, n_4990);
  nand g178529 (n_5770, g35, n_4999);
  fflopd g1384_reg(.CK (clock), .D (n_4551), .Q (g1384));
  fflopd g1351_reg(.CK (clock), .D (n_4589), .Q (g1351));
  fflopd g262_reg(.CK (clock), .D (n_4637), .Q (g262));
  not g179291 (n_6463, n_4868);
  fflopd g1008_reg(.CK (clock), .D (n_4677), .Q (g1008));
  fflopd g4983_reg(.CK (clock), .D (n_4682), .Q (g4983));
  nand g179443 (n_4872, n_4593, n_4871);
  nor g178641 (n_4870, n_1498, n_4341);
  nor g178637 (n_4869, n_4477, n_4782);
  nand g179483 (n_4868, g35, n_4481);
  nand g178634 (n_4867, g4112, n_4303);
  nor g178633 (n_4866, n_859, n_4500);
  nand g178632 (n_4865, n_4305, n_4288);
  nand g178448 (n_4864, g14673, g5933);
  nand g178425 (n_4863, g14597, g5248);
  nand g178458 (n_4862, g14749, g6625);
  nand g178473 (n_4861, g35, n_4450);
  nand g178450 (n_4860, g14705, g6287);
  nand g178451 (n_4858, g14673, g5941);
  nand g178434 (n_4857, g14597, g5240);
  nand g178449 (n_4856, n_1446, n_4453);
  nand g178418 (n_4855, n_4854, n_4449);
  nand g178417 (n_4853, g13906, g3941);
  nor g178630 (n_4852, n_4501, n_4503);
  nand g178398 (n_4851, g13881, g3582);
  nor g177972 (n_4850, n_4399, n_3789);
  nand g178002 (n_4849, n_2075, n_4410);
  nand g178003 (n_4848, n_2073, n_4519);
  nand g178005 (n_4847, n_2107, n_4412);
  nand g178006 (n_4846, n_2086, n_4394);
  nand g178011 (n_4845, n_2088, n_4408);
  nand g178015 (n_4844, n_33, n_4430);
  nor g178068 (n_4843, n_4419, n_4842);
  nor g178069 (n_4841, n_4413, n_899);
  nand g178416 (n_4840, g35, n_4839);
  nand g178083 (n_4838, n_3786, n_4428);
  nand g178084 (n_4837, n_3791, n_4439);
  nand g178085 (n_4836, n_3784, n_4440);
  nand g178086 (n_4835, n_3355, n_4441);
  nand g178087 (n_4834, n_3788, n_4442);
  nor g178111 (n_4833, n_4402, n_445);
  nor g178119 (n_4832, n_4416, n_4831);
  nor g178136 (n_4830, g691, n_4839);
  nand g178414 (n_4829, g13906, g3933);
  nand g178628 (n_4828, g681, n_4777);
  nand g178467 (n_4827, n_4486, n_3155);
  nor g178627 (n_4826, n_4269, n_4504);
  nor g178626 (n_4825, n_4507, n_4508);
  nor g178625 (n_4824, n_4271, n_4510);
  nand g178622 (n_4823, n_4044, n_4308);
  nor g178620 (n_4822, n_1529, n_4346);
  nand g178613 (n_4821, n_3339, n_4383);
  nand g178610 (n_4820, n_3738, n_4360);
  nand g178608 (n_4819, g4340, n_4314);
  nand g178399 (n_4818, g13881, g3590);
  nand g178603 (n_4817, g3263, n_4368);
  nand g178602 (n_4816, g3338, n_4300);
  nand g178599 (n_4815, g6657, n_4369);
  nand g178597 (n_4814, g25219, n_4298);
  nand g178595 (n_4813, g3965, n_4370);
  nand g178594 (n_4812, g5619, n_4371);
  wire w75, w76, w77, w78;
  nand g178336 (n_4811, w76, w78);
  nand g85 (w78, w77, n_170);
  not g84 (w77, n_4809);
  nand g83 (w76, w75, n_4809);
  not g82 (w75, n_170);
  wire w79, w80, w81, w82;
  nand g178338 (n_4810, w80, w82);
  nand g89 (w82, w81, n_1043);
  not g88 (w81, n_4809);
  nand g87 (w80, w79, n_4809);
  not g86 (w79, n_1043);
  wire w83, w84, w85, w86;
  nand g178339 (n_4808, w84, w86);
  nand g93 (w86, w85, n_239);
  not g92 (w85, n_4373);
  nand g91 (w84, w83, n_4373);
  not g90 (w83, n_239);
  nand g178355 (n_4807, n_527, n_4499);
  nand g178366 (n_4806, g14635, g5587);
  nor g178367 (n_4805, n_3872, n_4437);
  nor g178379 (n_4804, n_3871, n_4448);
  nand g178383 (n_4803, g13865, g3231);
  nand g178385 (n_4802, g13865, g3239);
  nand g178593 (n_4801, g5965, n_4372);
  nand g178470 (n_4800, g14749, g6633);
  nand g178447 (n_4799, g14705, g6279);
  nand g178589 (n_4798, g4040, n_4299);
  nor g178514 (n_4797, n_3870, n_4445);
  nand g178588 (n_4796, g2084, n_4295);
  not g178555 (n_4795, n_4999);
  not g178556 (n_4794, n_5114);
  not g178557 (n_4793, n_5005);
  not g178558 (n_4792, n_4993);
  not g178559 (n_4791, n_4990);
  nand g178584 (n_4790, g6311, n_4690);
  nand g178563 (n_4789, n_4787, n_2440);
  nand g178564 (n_4788, n_4787, n_2381);
  nand g178576 (n_4786, n_6019, n_4506);
  nand g178577 (n_4785, n_6011, n_4497);
  nand g178578 (n_4784, g1087, n_4292);
  nor g178579 (n_4783, n_3510, n_4782);
  nor g178516 (n_5480, n_9257, n_4432);
  nand g179466 (n_4879, g35, n_4670);
  fflopd g2848_reg(.CK (clock), .D (n_10194), .Q (g2848));
  nand g179475 (n_4876, g35, n_4668);
  fflopd g4401_reg(.CK (clock), .D (n_4429), .Q (g4401));
  fflopd g4859_reg(.CK (clock), .D (n_4505), .Q (g4859));
  fflopd g1211_reg(.CK (clock), .D (n_4385), .Q (g1211));
  fflopd g255_reg(.CK (clock), .D (n_4348), .Q (g255));
  fflopd g3325_reg(.CK (clock), .D (g13865), .Q (g16686));
  fflopd g3676_reg(.CK (clock), .D (g13881), .Q (g16722));
  fflopd g4027_reg(.CK (clock), .D (g13906), .Q (g16748));
  fflopd g5335_reg(.CK (clock), .D (g14597), .Q (g17639));
  not g178561 (n_5623, n_5036);
  nand g178203 (n_5377, n_4425, n_4433);
  nand g178202 (n_5378, n_4427, n_4434);
  fflopd g6027_reg(.CK (clock), .D (g14673), .Q (g17715));
  fflopd g5681_reg(.CK (clock), .D (g14635), .Q (g17678));
  fflopd g6373_reg(.CK (clock), .D (g14705), .Q (g17743));
  fflopd g6719_reg(.CK (clock), .D (g14749), .Q (g17764));
  fflopd g1395_reg(.CK (clock), .D (n_4431), .Q (g1395));
  fflopd g513_reg(.CK (clock), .D (n_4512), .Q (g513));
  fflopd g232_reg(.CK (clock), .D (n_4350), .Q (g232));
  fflopd g518_reg(.CK (clock), .D (n_4511), .Q (g518));
  nand g178220 (n_5384, n_4010, n_4513);
  nand g178217 (n_5382, n_4480, n_4403);
  nand g178895 (n_4781, g35, n_4366);
  nand g178661 (n_4780, g17316, n_4321);
  nand g178663 (n_4779, n_3306, n_4306);
  nand g178665 (n_4778, g446, n_4777);
  nand g178669 (n_4775, n_3066, n_4382);
  nor g178670 (n_4774, n_1728, n_4296);
  nand g178671 (n_4773, g17400, n_4344);
  nand g178674 (n_4772, g2643, n_4294);
  nand g178675 (n_4771, n_1553, n_4352);
  nand g178678 (n_4770, n_1566, n_4353);
  nand g178682 (n_4769, g847, n_4378);
  nand g178685 (n_4768, n_3371, n_4384);
  nand g178687 (n_4767, n_4787, n_2433);
  nand g179342 (n_4766, n_4458, n_4871);
  nand g179333 (n_4765, n_4250, n_4485);
  nand g179332 (n_4764, n_3968, n_4459);
  nand g178444 (n_4763, n_1444, n_4454);
  nor g179309 (n_4762, n_5381, n_4761);
  not g179270 (n_4760, n_4759);
  not g178777 (n_4758, n_4675);
  not g179246 (n_4757, n_4591);
  nand g179155 (n_4756, n_74, n_4761);
  nand g179141 (n_4755, n_3591, n_4460);
  nand g179139 (n_4754, n_3449, n_4461);
  nand g179126 (n_4753, n_3455, n_4466);
  nand g178805 (n_4752, n_4787, n_2452);
  nand g178806 (n_4751, n_4787, n_2432);
  nand g178807 (n_4750, n_4787, n_2373);
  wire w87, w88, w89, w90;
  nand g178808 (n_4749, w88, w90);
  nand g97 (w90, w89, n_1736);
  not g96 (w89, n_4218);
  nand g95 (w88, w87, n_4218);
  not g94 (w87, n_1736);
  wire w91, w92, w93, w94;
  nand g178809 (n_4748, w92, w94);
  nand g101 (w94, w93, n_1735);
  not g100 (w93, n_4217);
  nand g99 (w92, w91, n_4217);
  not g98 (w91, n_1735);
  wire w95, w96, w97, w98;
  nand g178814 (n_4747, w96, w98);
  nand g105 (w98, w97, g4801);
  not g104 (w97, n_4580);
  nand g103 (w96, w95, n_4580);
  not g102 (w95, g4801);
  wire w99, w100, w101, w102;
  nand g178816 (n_4746, w100, w102);
  nand g109 (w102, w101, n_1758);
  not g108 (w101, n_4245);
  nand g107 (w100, w99, n_4245);
  not g106 (w99, n_1758);
  nand g178817 (n_4745, n_3007, n_4787);
  nand g178818 (n_4744, n_2342, n_4787);
  nand g178822 (n_4743, n_2343, n_4787);
  nand g178823 (n_4742, n_3011, n_4787);
  nand g178824 (n_4741, n_2353, n_4787);
  nand g178826 (n_4740, n_3013, n_4787);
  nand g178827 (n_4739, g26801, n_4787);
  nand g178828 (n_4738, n_2372, n_4787);
  nand g178829 (n_4737, n_1567, n_4345);
  nand g178832 (n_4736, n_3009, n_4787);
  nand g178833 (n_4735, n_2344, n_4787);
  nand g178854 (n_4734, g35, n_4381);
  nand g178855 (n_4733, g35, n_4364);
  nand g178857 (n_4732, n_4100, n_4313);
  nand g178861 (n_4731, n_2340, n_4787);
  nand g178862 (n_4730, n_2341, n_4787);
  nand g178866 (n_4729, n_3005, n_4787);
  nand g178867 (n_4728, n_2708, n_4787);
  nand g178869 (n_4727, g35, n_4498);
  nand g178872 (n_4726, n_3582, n_4310);
  nand g178893 (n_4725, n_2715, n_4415);
  nand g178659 (n_4724, n_4143, n_4331);
  nand g178905 (n_4723, g5022, n_4316);
  nand g178913 (n_4722, g650, n_4720);
  nand g178915 (n_4721, g718, n_4720);
  nand g178920 (n_4719, n_2646, n_4386);
  nand g178921 (n_4718, g645, n_4720);
  nand g178924 (n_4717, g655, n_4720);
  nand g178929 (n_4716, g4122, n_4533);
  nand g178930 (n_4715, g661, n_4720);
  nand g178934 (n_4714, g4991, n_4517);
  nand g178938 (n_4713, n_2644, n_4495);
  nand g178940 (n_4712, n_2061, n_4711);
  nand g178942 (n_4710, n_4262, n_4340);
  nand g178945 (n_4709, n_4270, n_4339);
  nand g178946 (n_4708, n_869, n_4293);
  nand g178949 (n_4707, g837, n_4290);
  nand g178951 (n_4706, g837, n_4315);
  nand g178952 (n_4705, n_4186, n_4351);
  nand g179116 (n_4704, n_3464, n_4462);
  nand g179112 (n_4703, n_3436, n_4463);
  nand g179096 (n_4701, n_3439, n_4465);
  nand g179093 (n_4700, n_3626, n_4467);
  nand g178445 (n_4699, g14635, g5595);
  nand g179084 (n_4698, n_844, n_4478);
  nand g179046 (n_4694, n_3444, n_4464);
  not g179041 (n_5286, n_4878);
  fflopd g4072_reg(.CK (clock), .D (n_4304), .Q (g4072));
  not g179282 (n_5310, n_4693);
  nand g178991 (n_4873, n_4692, n_8312);
  nand g178989 (n_4874, n_4691, g28753);
  nand g178977 (n_4875, n_4690, n_8355);
  fflopd g1489_reg(.CK (clock), .D (n_4307), .Q (g1489));
  not g179034 (n_5280, n_4568);
  nand g178965 (n_5520, g35, n_4297);
  fflopd g4414_reg(.CK (clock), .D (n_4397), .Q (g7257));
  nand g178715 (n_5300, n_1851, n_4380);
  not g179287 (n_5289, n_4689);
  nand g178744 (n_5313, n_1880, n_4376);
  nor g178971 (n_5392, n_9257, g28753);
  nor g178973 (n_5389, n_9257, n_8355);
  fflopd g417_reg(.CK (clock), .D (n_4421), .Q (g417));
  nor g178967 (n_5386, n_9257, n_8312);
  not g178800 (n_5445, n_4557);
  not g178802 (n_5450, n_4538);
  fflopd g5821_reg(.CK (clock), .D (n_4349), .Q (g5821));
  not g178803 (n_5452, n_4536);
  not g178804 (n_5454, n_4532);
  fflopd g1554_reg(.CK (clock), .D (n_4514), .Q (g1554));
  not g178801 (n_5448, n_4540);
  nor g178770 (n_5492, g1312, n_4342);
  nor g178769 (n_7889, g969, n_4338);
  not g179295 (n_8904, n_4673);
  nand g178925 (n_4688, n_1616, n_4629);
  nand g179388 (n_4687, n_3911, n_4228);
  nand g179390 (n_4686, n_3962, n_4229);
  nand g179393 (n_4685, n_3487, n_10378);
  nand g179399 (n_4684, n_3957, n_4232);
  nand g179412 (n_4683, n_4222, n_4422);
  nand g179423 (n_4682, n_3909, n_4221);
  nand g179371 (n_4681, n_3915, n_4231);
  nand g179436 (n_4680, n_3913, n_4227);
  nand g179437 (n_4679, n_3914, n_4230);
  nand g178919 (n_4678, n_1443, n_4131);
  nand g178914 (n_4677, n_4137, n_4144);
  nand g178903 (n_4676, n_1454, n_4631);
  nand g178894 (n_4675, n_542, n_4134);
  nand g178891 (n_4674, g1404, n_4172);
  nand g179487 (n_4673, g35, n_4672);
  not g179499 (n_4671, n_4670);
  not g179501 (n_4669, n_4668);
  nand g178889 (n_4667, n_2652, n_4130);
  nand g178888 (n_4666, g1384, n_4187);
  nand g178886 (n_4665, g35, n_4185);
  nand g178885 (n_4664, n_2409, n_4139);
  nand g178876 (n_4663, g14125, n_5795);
  nor g178643 (g32185, n_3118, n_10380);
  nand g178874 (n_4661, g35, n_4152);
  nand g178873 (n_4660, n_1456, n_4627);
  not g177630 (n_4658, n_4451);
  nand g178871 (n_4657, g35, n_4656);
  nand g178863 (n_4655, n_2147, n_4115);
  wire w103, w104, w105, w106;
  nand g178337 (n_4654, w104, w106);
  nand g113 (w106, w105, n_1759);
  not g112 (w105, n_4072);
  nand g111 (w104, w103, n_4072);
  not g110 (w103, n_1759);
  wire w107, w108, w109, w110;
  nand g178344 (n_4653, w108, w110);
  nand g117 (w110, w109, n_1757);
  not g116 (w109, n_4071);
  nand g115 (w108, w107, n_4071);
  not g114 (w107, n_1757);
  nand g178860 (n_4652, g35, n_4156);
  nand g178856 (n_4651, g35, n_4158);
  nand g178852 (n_4650, g35, n_4161);
  nand g178851 (n_4649, g35, n_4162);
  nand g178565 (n_4647, n_4646, n_4118);
  nand g178580 (n_4645, n_3834, n_4151);
  nand g178582 (n_4644, g6381, n_4111);
  nand g178583 (n_4643, g6381, n_4103);
  nand g178590 (n_4642, g5689, n_4119);
  nand g178591 (n_4641, g3689, n_4120);
  nand g178592 (n_4640, g6035, n_4121);
  nand g178598 (n_4639, g6727, n_4102);
  nand g178601 (n_4638, g278, n_4184);
  nand g178615 (n_4637, n_4135, n_4055);
  nand g178629 (n_4636, n_21, n_4157);
  nand g178640 (n_4635, n_62, n_4155);
  nand g178644 (n_4633, n_189, n_4148);
  nor g178655 (n_4632, n_4631, n_4176);
  nor g178656 (n_4630, n_4629, n_4177);
  nor g178657 (n_4628, n_4627, n_4178);
  nor g178662 (n_4626, n_66, n_4625);
  nand g178664 (n_4624, g20899, n_4104);
  nand g178679 (n_4623, n_4114, n_5760);
  nand g178686 (n_4622, n_4110, n_6456);
  nand g178850 (n_4621, g35, n_4146);
  nand g178849 (n_4620, g35, n_4163);
  nand g178845 (n_4619, g4369, n_9257);
  nand g178839 (n_4618, n_7031, n_4116);
  nand g178838 (n_4617, n_7035, n_4112);
  nand g178837 (n_4616, n_6888, n_4117);
  nand g178836 (n_4615, n_6886, n_4108);
  nand g178835 (n_4614, n_5789, n_4113);
  nor g178830 (n_4613, g6195, n_4595);
  wire w111, w112, w113, w114;
  nand g178813 (n_4612, w112, w114);
  nand g121 (w114, w113, g482);
  not g120 (w113, n_4238);
  nand g119 (w112, w111, n_4238);
  not g118 (w111, g482);
  not g178776 (n_4611, n_4502);
  not g178778 (n_4610, n_4414);
  not g178780 (n_4609, n_4406);
  not g178781 (n_4608, n_4405);
  not g178783 (n_4607, n_4401);
  not g178782 (n_4606, n_4404);
  not g178785 (n_4605, n_4398);
  not g178786 (n_4604, n_4396);
  not g178789 (n_4603, n_4392);
  not g178790 (n_4602, n_4391);
  not g178791 (n_4601, n_4390);
  not g178792 (n_4600, n_4389);
  not g178793 (n_4599, n_4388);
  not g178794 (n_4598, n_4597);
  nor g178812 (n_4596, g6541, n_4595);
  fflopd g429_reg(.CK (clock), .D (n_4282), .Q (g429));
  nand g179454 (n_4759, n_2881, n_4594);
  nor g179458 (n_4882, n_3920, n_4224);
  nand g179471 (n_4693, g35, n_4240);
  nand g179477 (n_4689, g691, n_4258);
  not g179512 (n_4877, n_4593);
  fflopd g452_reg(.CK (clock), .D (n_4276), .Q (g452));
  fflopd g424_reg(.CK (clock), .D (n_4261), .Q (g424));
  fflopd g884_reg(.CK (clock), .D (g14125), .Q (g14147));
  fflopd g437_reg(.CK (clock), .D (n_4280), .Q (g437));
  nor g178774 (n_5036, g1319, n_2201);
  nand g178707 (n_5267, n_3415, n_4265);
  fflopd g962_reg(.CK (clock), .D (n_4252), .Q (g962));
  fflopd g1306_reg(.CK (clock), .D (n_4236), .Q (g1306));
  nor g178720 (g27831, n_4592, n_4142);
  fflopd g4646_reg(.CK (clock), .D (n_4154), .Q (g4646));
  fflopd g499_reg(.CK (clock), .D (n_4274), .Q (g499));
  nor g178734 (n_4990, n_4526, n_4539);
  fflopd g174_reg(.CK (clock), .D (n_4272), .Q (g174));
  fflopd g168_reg(.CK (clock), .D (n_4273), .Q (g168));
  fflopd g4633_reg(.CK (clock), .D (n_4166), .Q (g4633));
  nor g179478 (n_4914, n_9257, n_4564);
  nor g178727 (n_4999, n_4528, n_4535);
  nor g178729 (n_5114, n_4523, n_4537);
  nor g178730 (n_5005, n_4522, n_4556);
  nor g178731 (n_4993, n_4525, n_4531);
  fflopd g405_reg(.CK (clock), .D (n_4191), .Q (g405));
  fflopd g847_reg(.CK (clock), .D (n_4266), .Q (g847));
  nand g179367 (n_4591, n_1197, n_4220);
  nand g178941 (n_4590, g4664, n_4263);
  nand g178944 (n_4589, n_3733, n_4145);
  nand g178932 (n_4588, g4349, n_4279);
  nand g179339 (n_4587, n_5549, n_4594);
  nand g179338 (n_4586, n_2828, n_4594);
  nand g179337 (n_4585, n_994, n_4594);
  nand g179331 (n_4584, n_9257, n_5503);
  nand g179325 (n_4583, g35, n_4226);
  nand g179318 (n_4582, n_1445, n_4521);
  nand g179317 (n_4581, n_1299, n_4580);
  nand g179310 (n_4579, n_2771, n_4594);
  not g179284 (n_4578, n_4782);
  not g179265 (n_4577, n_4494);
  not g179254 (n_4576, n_4509);
  not g179253 (n_4575, n_4515);
  not g179252 (n_4574, n_4516);
  not g179249 (n_4573, n_4518);
  not g179248 (n_4572, n_4520);
  not g179244 (n_4571, n_4387);
  not g179241 (n_4570, n_4367);
  not g179240 (n_4569, n_4365);
  nand g179178 (n_4568, g4776, n_4580);
  nor g179157 (n_4567, n_4457, n_4216);
  nand g179149 (n_4566, n_1592, n_4672);
  nand g179146 (n_4565, n_2721, n_4564);
  nor g179140 (n_4563, g9553, n_4248);
  nand g179137 (n_4562, n_532, n_4208);
  nand g179119 (n_4561, g753, n_4560);
  nand g179117 (n_4559, n_1294, n_4199);
  nand g179114 (n_4558, n_751, n_4201);
  nand g178995 (n_4557, g35, n_4556);
  nand g179110 (n_4555, n_3184, n_4214);
  nor g179108 (n_4554, n_3230, n_4527);
  nand g179106 (n_4553, g1413, n_4242);
  nand g179105 (n_4552, n_502, n_4204);
  nand g179100 (n_4551, n_4205, n_4035);
  nand g179098 (n_4550, n_496, n_4209);
  nand g179097 (n_4549, n_1343, n_4207);
  nand g179094 (n_4548, n_3951, n_4215);
  nand g179092 (n_4547, g1070, n_4244);
  nand g179091 (n_4546, n_1181, n_4210);
  nand g179085 (n_4545, n_933, n_4212);
  nand g179051 (n_4544, n_913, n_4564);
  nand g179049 (n_4543, n_4542, n_4249);
  not g179044 (n_4541, n_5276);
  nand g179010 (n_4540, g35, n_4539);
  nand g179011 (n_4538, g35, n_4537);
  nand g179012 (n_4536, g35, n_4535);
  not g179028 (n_4534, n_4533);
  nand g179014 (n_4532, g35, n_4531);
  not g179024 (n_4530, n_4317);
  nand g178959 (n_8351, g6500, n_4528);
  nand g179164 (n_4880, n_1996, n_4247);
  nand g179166 (n_4696, g482, n_4239);
  nor g179163 (n_4912, n_3880, n_4527);
  nand g178960 (n_8359, g3106, n_4526);
  nand g178961 (n_8382, g5462, n_4525);
  not g179278 (n_6949, n_4524);
  not g179283 (n_4920, n_4490);
  nand g178957 (n_8357, g3808, n_4523);
  nand g178958 (n_8384, g5808, n_4522);
  fflopd g401_reg(.CK (clock), .D (n_4190), .Q (g401));
  nand g178963 (n_5175, n_2429, n_4147);
  fflopd g2975_reg(.CK (clock), .D (n_4132), .Q (g2975));
  nand g179192 (n_4878, g4584, n_4521);
  fflopd g441_reg(.CK (clock), .D (n_4278), .Q (g441));
  fflopd g4145_reg(.CK (clock), .D (n_4213), .Q (new_g6946_));
  nor g178982 (n_5243, n_9257, n_4285);
  nor g178981 (n_5270, n_9257, n_4531);
  nor g178980 (n_5204, n_1418, n_4595);
  nor g178979 (n_5023, n_9257, n_4556);
  nor g178978 (n_5191, n_1706, n_4595);
  nor g178976 (n_5110, n_9257, n_4287);
  nor g178975 (n_5240, n_9257, n_4535);
  nor g178986 (n_5011, n_9257, n_4539);
  nor g178994 (n_5164, n_1417, n_4595);
  nor g178974 (n_5146, n_1724, n_4595);
  nor g178993 (n_5103, n_1420, n_4595);
  nor g178992 (n_5187, n_1422, n_4595);
  nor g178990 (n_5214, n_1720, n_4595);
  nor g178972 (n_5168, n_1421, n_4595);
  nor g178985 (n_5081, n_1710, n_4595);
  nor g178970 (n_5091, n_1722, n_4595);
  nor g178969 (n_5096, n_1715, n_4595);
  nor g178968 (n_5106, n_1721, n_4595);
  nor g178988 (n_5183, n_1707, n_4595);
  nor g178987 (n_5209, n_1425, n_4595);
  nor g178984 (n_8166, n_9257, n_4286);
  nor g178983 (n_5251, n_9257, n_4537);
  nor g179015 (n_5049, n_1548, n_4595);
  nor g179013 (n_5052, n_2811, n_4595);
  nor g179009 (n_5069, n_2796, n_4595);
  nor g179008 (n_4978, n_1194, n_4595);
  nor g179007 (n_5221, n_2957, n_4595);
  nor g179006 (n_5123, n_607, n_4595);
  nor g179005 (n_5017, n_591, n_4595);
  nor g179004 (n_5258, n_969, n_4595);
  nor g179003 (n_4973, n_1705, n_4595);
  nor g179002 (n_5261, n_2733, n_4595);
  nor g179001 (n_4957, n_618, n_4595);
  nor g179000 (n_5134, n_838, n_4595);
  nor g178999 (n_5037, n_1419, n_4595);
  nor g178998 (n_5264, n_2766, n_4595);
  nor g178997 (n_5255, n_600, n_4595);
  nor g178996 (n_5233, n_594, n_4595);
  nor g179017 (n_5040, n_2738, n_4595);
  nor g179016 (n_5225, n_2761, n_4595);
  not g179292 (n_6512, n_4487);
  not g179289 (n_7046, n_4488);
  not g179294 (n_4932, n_4720);
  nand g179376 (n_4520, n_701, n_3995);
  nand g178887 (n_4519, n_1406, n_4438);
  nand g179377 (n_4518, n_1198, n_3993);
  nand g179380 (n_4517, g35, n_3967);
  nand g179384 (n_4516, n_587, n_4045);
  nand g179385 (n_4515, n_1190, n_3905);
  nand g179386 (n_4514, n_3477, n_3940);
  nand g178884 (n_4513, g1430, n_3885);
  nand g179391 (n_4512, n_3524, n_3937);
  nand g179394 (n_4511, n_3516, n_3936);
  nand g179396 (n_4510, n_4005, n_4004);
  nand g179398 (n_4509, g4776, n_4194);
  nand g179400 (n_4508, n_3974, n_3705);
  nand g179402 (n_4507, n_3704, n_3901);
  nand g179403 (n_4506, n_3129, n_4006);
  nand g179405 (n_4505, n_3400, n_3912);
  nand g179406 (n_4504, n_4003, n_4002);
  nand g179410 (n_4503, n_3899, n_3702);
  nand g178882 (n_4502, g17813, g5579);
  nand g179413 (n_4501, n_3701, n_3900);
  nand g179417 (n_4500, n_4046, n_3742);
  nand g178875 (n_4499, n_4854, n_3879);
  nand g179420 (n_4498, n_3719, n_4050);
  nand g179428 (n_4497, n_3103, n_3997);
  nand g179432 (n_4496, g732, n_4195);
  nand g179441 (n_4495, n_2253, n_4031);
  nand g179442 (n_4494, n_842, n_3966);
  nand g178865 (n_4493, n_4492, n_4475);
  nand g178859 (n_4491, n_6357, n_4473);
  nand g179472 (n_4490, g35, n_4363);
  nand g178853 (n_4489, n_6580, n_4483);
  nand g179480 (n_4488, g35, n_4001);
  nand g179484 (n_4487, g35, n_4011);
  nand g178848 (n_4486, g5069, n_9257);
  not g179490 (n_4485, n_4233);
  nand g178847 (n_4484, g6727, n_4483);
  nand g178846 (n_4482, g4423, n_9257);
  nand g179620 (n_4481, g1585, n_4480);
  nand g178844 (n_4479, g3689, n_4455);
  nand g179655 (n_4478, n_3509, n_4477);
  nand g178842 (n_4476, g6381, n_4475);
  nand g178841 (n_4474, g6035, n_4473);
  nand g178840 (n_4472, g5689, n_4469);
  nor g178834 (n_4471, n_4030, n_1547);
  nand g178831 (n_4470, n_6359, n_4469);
  not g179750 (n_4467, n_4235);
  not g179760 (n_4466, n_4253);
  not g179762 (n_4465, n_4254);
  not g179768 (n_4464, n_4255);
  not g179772 (n_4463, n_4256);
  not g179775 (n_4462, n_4257);
  not g179788 (n_4461, n_4259);
  not g179790 (n_4460, n_4260);
  not g179796 (n_4459, n_4527);
  nand g179848 (n_4458, n_4457, n_4426);
  nand g178825 (n_4456, n_6582, n_4455);
  nand g178821 (n_4454, n_3340, n_3883);
  nand g178820 (n_4453, n_3341, n_3882);
  wire w115, w116, w117, w118;
  nand g178815 (n_4452, w116, w118);
  nand g125 (w118, w117, g671);
  not g124 (w117, n_4140);
  nand g123 (w116, w115, n_4140);
  not g122 (w115, g671);
  nand g177858 (n_4451, n_4283, n_3921);
  wire w119, w120, w121, w122;
  nand g178811 (n_4450, w120, w122);
  nand g129 (w122, w121, g8358);
  not g128 (w121, n_3759);
  nand g127 (w120, w119, n_3759);
  not g126 (w119, g8358);
  wire w123, w124, w125, w126;
  nand g178810 (n_4449, w124, w126);
  nand g133 (w126, w125, g822);
  not g132 (w125, n_4101);
  nand g131 (w124, w123, n_4101);
  not g130 (w123, g822);
  nor g178684 (n_4448, n_4089, n_3616);
  nor g178683 (n_4447, n_3894, n_5462);
  nor g178681 (n_4446, n_4094, n_5464);
  nor g178680 (n_4445, n_4093, n_4444);
  nor g178677 (n_4443, n_3924, n_5466);
  nor g178653 (n_4442, n_4393, n_3833);
  nor g178652 (n_4441, n_4407, n_3830);
  nor g178651 (n_4440, n_4411, n_3799);
  nor g178650 (n_4439, n_4438, n_3804);
  nor g178562 (n_4437, n_4097, n_3614);
  nand g178596 (n_4436, g3614, n_4692);
  nand g178600 (n_4435, g5272, n_4691);
  nand g178604 (n_4434, g17320, n_3878);
  nand g178611 (n_4433, g17423, n_3875);
  nor g178616 (n_4432, g2625, n_3869);
  nand g178618 (n_4431, n_10216, n_3896);
  nand g178636 (n_4430, n_592, n_3868);
  nand g178639 (n_4429, n_6, n_3874);
  nor g178649 (n_4428, n_4409, n_3798);
  nand g179679 (n_4668, n_4424, n_4427);
  nand g179704 (n_4593, g5041, n_4426);
  fflopd g2999_reg(.CK (clock), .D (n_3887), .Q (g2999));
  nand g179672 (n_4670, n_4424, n_4425);
  nand g179467 (n_4524, g35, n_4423);
  fflopd g4287_reg(.CK (clock), .D (n_4088), .Q (g9019));
  nand g179707 (n_4761, new_g6832_, n_4480);
  fflopd g385_reg(.CK (clock), .D (n_4041), .Q (g385));
  nand g178708 (n_4839, g681, n_3866);
  fflopd g4462_reg(.CK (clock), .D (n_3888), .Q (g4462));
  fflopd g2917_reg(.CK (clock), .D (n_4033), .Q (g2917));
  fflopd g667_reg(.CK (clock), .D (n_3929), .Q (g667));
  nand g179473 (n_4782, g35, n_4422);
  fflopd g6715_reg(.CK (clock), .D (g17871), .Q (g14749));
  fflopd g6369_reg(.CK (clock), .D (g17845), .Q (g14705));
  fflopd g4023_reg(.CK (clock), .D (g16955), .Q (g13906));
  fflopd g3321_reg(.CK (clock), .D (g16874), .Q (g13865));
  fflopd g3672_reg(.CK (clock), .D (g16924), .Q (g13881));
  fflopd g5813_reg(.CK (clock), .D (n_3960), .Q (g5813));
  fflopd g6159_reg(.CK (clock), .D (n_3955), .Q (g6159));
  fflopd g3462_reg(.CK (clock), .D (n_3934), .Q (g3462));
  fflopd g3111_reg(.CK (clock), .D (n_3943), .Q (g3111));
  fflopd g4836_reg(.CK (clock), .D (n_4019), .Q (g4836));
  fflopd g4659_reg(.CK (clock), .D (n_3867), .Q (g4659));
  fflopd g6533_reg(.CK (clock), .D (n_3907), .Q (g6533));
  fflopd g3490_reg(.CK (clock), .D (n_3933), .Q (g3490));
  fflopd g5841_reg(.CK (clock), .D (n_3946), .Q (g5841));
  fflopd g3139_reg(.CK (clock), .D (n_3942), .Q (g3139));
  fflopd g5148_reg(.CK (clock), .D (n_3950), .Q (g5148));
  fflopd g3841_reg(.CK (clock), .D (n_3927), .Q (g3841));
  fflopd g370_reg(.CK (clock), .D (n_3895), .Q (g370));
  fflopd g6187_reg(.CK (clock), .D (n_3953), .Q (g6187));
  fflopd g6023_reg(.CK (clock), .D (g17819), .Q (g14673));
  fflopd g6505_reg(.CK (clock), .D (n_3931), .Q (g6505));
  fflopd g5677_reg(.CK (clock), .D (g17813), .Q (g14635));
  fflopd g5331_reg(.CK (clock), .D (g17787), .Q (g14597));
  fflopd g3179_reg(.CK (clock), .D (n_4032), .Q (g3179));
  fflopd g4340_reg(.CK (clock), .D (n_4087), .Q (g4340));
  fflopd g6227_reg(.CK (clock), .D (n_4039), .Q (g6227));
  fflopd g3530_reg(.CK (clock), .D (n_4022), .Q (g3530));
  fflopd g5535_reg(.CK (clock), .D (n_4040), .Q (g5535));
  fflopd g5881_reg(.CK (clock), .D (n_4034), .Q (g5881));
  nand g179486 (n_4720, g35, n_4059);
  nand g179368 (n_4421, n_4043, n_3842);
  nand g178890 (n_4420, g1395, n_3897);
  nand g178897 (n_4419, g16874, g3223);
  nand g178898 (n_4418, g728, n_4417);
  nand g178899 (n_4416, g16874, g3215);
  nand g179365 (n_4415, g35, n_3945);
  nand g178906 (n_4414, g16924, g3566);
  nand g178907 (n_4413, g16924, g3574);
  nand g178909 (n_4412, n_609, n_4411);
  nand g178911 (n_4410, n_726, n_4409);
  nand g178912 (n_4408, n_828, n_4407);
  nand g178916 (n_4406, g17871, g6609);
  nand g178917 (n_4405, g16955, g3917);
  nand g178918 (n_4404, g16955, g3925);
  nand g178922 (n_4403, g17404, n_3889);
  nand g178923 (n_4402, g17787, g5232);
  nand g178927 (n_4401, g4116, n_4400);
  nand g178928 (n_4399, g17871, g6617);
  nand g178935 (n_4398, n_664, n_4106);
  nand g178936 (n_4397, n_2033, n_3877);
  nand g178937 (n_4396, g17787, g5224);
  nand g178943 (n_4395, g278, n_4183);
  nand g178947 (n_4394, n_619, n_4393);
  nand g178948 (n_4392, g17819, g5925);
  nand g178950 (n_4391, g17819, g5917);
  nand g178953 (n_4390, g17813, g5571);
  nand g178954 (n_4389, g17845, g6263);
  nand g178955 (n_4388, g17845, g6271);
  nand g179356 (n_4387, g1046, n_4330);
  nand g179353 (n_4386, n_2208, n_4007);
  nand g179352 (n_4385, n_3473, n_3956);
  not g179018 (n_4384, n_4165);
  not g179019 (n_4383, n_4164);
  not g179021 (n_4382, n_4160);
  not g179023 (n_4381, n_4141);
  not g179025 (n_4380, n_4379);
  not g179030 (n_4378, n_4377);
  not g179031 (n_4376, n_4375);
  not g179035 (n_4372, n_4522);
  not g179036 (n_4371, n_4525);
  not g179037 (n_4370, n_4523);
  not g179038 (n_4369, n_4528);
  not g179039 (n_4368, n_4526);
  nand g179346 (n_4367, n_707, n_3971);
  nand g179345 (n_4366, g1211, n_4246);
  nand g179344 (n_4365, n_530, n_4012);
  nor g179050 (n_4364, n_10400, n_4363);
  nand g179053 (n_4361, n_4358, n_3687);
  nand g179054 (n_4360, n_2376, n_4060);
  nand g179058 (n_4359, n_4358, n_3680);
  nand g179059 (n_4357, n_4358, n_3681);
  nand g179061 (n_4356, n_4358, n_3683);
  nand g179064 (n_4355, n_4358, n_3686);
  nand g179066 (n_4354, n_4358, n_3682);
  nand g179079 (n_4353, n_3772, n_4064);
  nand g179080 (n_4352, n_3774, n_4062);
  nand g179081 (n_4351, g4793, n_4083);
  nand g179087 (n_4350, n_3754, n_4053);
  nand g179089 (n_4349, n_3459, n_4054);
  nand g179090 (n_4348, n_3264, n_4066);
  nor g179101 (n_4346, g1413, n_4241);
  nand g179111 (n_4345, n_3287, n_4061);
  nand g179118 (n_4344, n_4343, n_4320);
  nand g179120 (n_4342, n_3123, n_4069);
  nor g179122 (n_4341, g1070, n_4243);
  nand g179124 (n_4340, g4698, n_4075);
  nand g179130 (n_4339, g4888, n_4077);
  nand g179135 (n_4338, n_3105, n_4070);
  nand g179138 (n_4337, g1041, n_4082);
  nand g179143 (n_4336, n_1298, n_4322);
  nand g179144 (n_4335, n_1368, n_4326);
  nand g179145 (n_4334, n_805, n_4324);
  nand g179147 (n_4333, n_165, n_4332);
  nor g179148 (n_4331, g1046, n_4330);
  nand g179150 (n_4329, n_221, n_4328);
  nand g179151 (n_4327, n_1617, n_4326);
  nand g179152 (n_4325, n_1457, n_4324);
  nand g179154 (n_4323, n_1455, n_4322);
  nand g179156 (n_4321, n_4319, n_4320);
  nand g179161 (n_4317, n_1040, n_4015);
  nand g179335 (n_4316, g35, n_3996);
  nand g179334 (n_4315, g35, n_4020);
  nor g179330 (n_4314, n_2423, n_3902);
  nand g179328 (n_4313, g35, n_4051);
  nand g179327 (n_4312, g35, n_4014);
  nand g179326 (n_4311, g35, n_4009);
  not g179238 (n_4310, n_4136);
  not g179245 (n_4309, n_4189);
  not g179247 (n_4308, n_4281);
  not g179250 (n_4307, n_4277);
  not g179251 (n_4306, n_4275);
  not g179258 (n_4305, n_4268);
  not g179260 (n_4304, n_4267);
  not g179269 (n_4303, n_4302);
  nand g179312 (n_4301, g351, n_9257);
  not g179272 (n_4300, n_4631);
  not g179279 (n_4299, n_4629);
  not g179281 (n_4298, n_4627);
  nor g179311 (n_4297, g5046, n_4871);
  not g179290 (n_4296, n_7798);
  nor g179308 (n_4295, n_6016, n_4332);
  nor g179307 (n_4294, n_5383, n_4328);
  nand g179297 (n_4293, n_2969, n_4036);
  nand g179300 (n_4292, n_4291, n_4320);
  nand g179304 (n_4290, n_3570, n_4048);
  nand g179165 (n_4711, g837, n_3918);
  nand g178956 (n_4597, g35, g4423);
  not g179042 (n_4690, n_4289);
  not g179271 (n_4777, n_4288);
  nand g179169 (n_4533, g4064, n_4057);
  fflopd g1576_reg(.CK (clock), .D (n_4099), .Q (g10527));
  fflopd g5467_reg(.CK (clock), .D (n_3906), .Q (g5467));
  nand g179224 (n_5276, g518, n_4063);
  not g179288 (n_8355, n_4287);
  fflopd g5495_reg(.CK (clock), .D (n_3964), .Q (g5495));
  not g179045 (n_8312, n_4286);
  fflopd g5120_reg(.CK (clock), .D (n_3922), .Q (g5120));
  fflopd g3813_reg(.CK (clock), .D (n_3928), .Q (g3813));
  fflopd g3881_reg(.CK (clock), .D (n_4028), .Q (g3881));
  fflopd g5188_reg(.CK (clock), .D (n_4024), .Q (g5188));
  fflopd g6573_reg(.CK (clock), .D (n_4037), .Q (g6573));
  not g179293 (g28753, n_4285);
  not g179296 (n_4787, n_4595);
  nand g179372 (n_4282, n_3566, n_3844);
  nand g179373 (n_4281, n_955, n_3846);
  nand g179374 (n_4280, n_3565, n_3847);
  nand g179375 (n_4279, g35, n_3748);
  nand g179378 (n_4278, n_3564, n_3803);
  nand g179379 (n_4277, g35, n_3727);
  nand g179381 (n_4276, n_3563, n_3764);
  nand g179383 (n_4275, n_945, n_3763);
  nand g179389 (n_4274, n_3315, n_3725);
  nand g179392 (n_4273, n_3430, n_3762);
  nand g179395 (n_4272, n_3581, n_3780);
  nand g179397 (n_4271, n_3723, n_3794);
  nand g179404 (n_4270, g4894, n_4076);
  nand g179409 (n_4269, n_3721, n_3793);
  nand g179414 (n_4268, n_1336, n_3743);
  nand g179421 (n_4267, g35, n_3814);
  nand g179429 (n_4266, n_3556, n_3836);
  nand g179431 (n_4265, g4608, n_3734);
  nand g179434 (n_4264, g35, n_3832);
  nand g179435 (n_4263, g35, n_3835);
  nand g179440 (n_4262, g4704, n_4074);
  nand g179369 (n_4261, n_3567, n_3843);
  nand g179990 (n_4260, n_1004, n_3659);
  nand g179983 (n_4259, n_942, n_3664);
  nand g179973 (n_4258, n_4223, n_3641);
  nand g179934 (n_4257, n_866, n_3660);
  nand g179917 (n_4256, n_792, n_3640);
  nand g179895 (n_4255, n_1319, n_3637);
  nand g179873 (n_4254, n_1246, n_3635);
  nand g179863 (n_4253, n_779, n_3638);
  nand g179838 (n_4252, n_3402, n_3685);
  nand g179830 (n_4250, g35, n_3655);
  not g179489 (n_4249, n_4042);
  not g179497 (n_4248, n_3998);
  not g179500 (n_4247, n_4246);
  not g179502 (n_4245, n_3989);
  not g179505 (n_4244, n_4243);
  not g179507 (n_4242, n_4241);
  not g179511 (n_4240, g351);
  not g179514 (n_4239, n_4238);
  nand g179828 (n_4237, g35, n_3692);
  nand g179823 (n_4236, n_3398, n_3684);
  nand g179813 (n_4235, n_770, n_3675);
  nand g179548 (n_4233, n_960, n_3674);
  nand g179594 (n_4232, g4933, n_3652);
  nand g179597 (n_4231, g4743, n_3650);
  nand g179602 (n_4230, g4754, n_3648);
  nand g179603 (n_4229, g4944, n_3644);
  nand g179604 (n_4228, g4955, n_3654);
  nand g179605 (n_4227, g4765, n_3646);
  nor g179617 (n_4226, n_4225, n_4219);
  nand g179630 (n_4224, n_3673, n_4223);
  nand g179636 (n_4222, n_1805, n_3865);
  nand g179660 (n_4221, g4983, n_3642);
  nand g179664 (n_4220, n_4225, n_4219);
  nor g179681 (n_4218, new_g6832_, n_3863);
  nor g179682 (n_4217, new_g6832_, n_3864);
  nand g179808 (n_4216, n_3862, n_3678);
  not g179784 (n_4215, n_3910);
  not g179748 (n_4214, n_4084);
  not g179751 (n_4213, n_3973);
  not g179752 (n_4212, n_3963);
  not g179753 (n_4211, n_3961);
  not g179756 (n_4210, n_3959);
  not g179759 (n_4209, n_3954);
  not g179761 (n_4208, n_3952);
  not g179763 (n_4207, n_3949);
  not g179765 (n_4206, n_3948);
  not g179766 (n_4205, n_3947);
  not g179769 (n_4204, n_3941);
  not g179770 (n_4203, n_3939);
  not g179771 (n_4202, n_3938);
  not g179773 (n_4201, n_3932);
  not g179774 (n_4200, n_3930);
  not g179776 (n_4199, n_3926);
  not g179778 (n_4198, n_3925);
  not g179779 (n_4197, n_3923);
  not g179781 (n_4196, n_3919);
  nand g179479 (n_4287, g4688, n_3761);
  nand g179453 (n_4302, g35, n_3801);
  nand g179459 (n_4288, g35, n_4058);
  not g179798 (n_4560, n_4195);
  nand g179485 (n_4285, g4646, n_3817);
  not g179516 (n_4521, n_4422);
  not g179517 (n_4580, n_4194);
  not g179515 (n_4564, n_3991);
  not g179801 (n_8302, n_9193);
  not g179518 (n_5503, g2724);
  fflopd g4273_reg(.CK (clock), .D (n_3855), .Q (g4273));
  nand g180020 (n_4527, n_4193, n_3658);
  nand g179697 (n_4672, g11678, n_3679);
  nand g179474 (n_4556, g4681, n_3808);
  nand g179470 (n_4627, g35, n_3984);
  nand g179468 (n_4629, g35, n_3982);
  nand g179461 (n_4531, g4674, n_3812);
  nand g179460 (n_4631, g35, n_3983);
  fflopd g1442_reg(.CK (clock), .D (n_3728), .Q (g1442));
  fflopd g5170_reg(.CK (clock), .D (n_3665), .Q (g5170));
  fflopd g6555_reg(.CK (clock), .D (n_3670), .Q (g6555));
  fflopd g6209_reg(.CK (clock), .D (n_3671), .Q (g6209));
  not g179800 (n_4594, n_5880);
  nand g179482 (n_7798, n_575, n_4192);
  nand g179481 (n_7611, n_1216, n_4192);
  nand g179488 (n_4595, g35, n_4174);
  nand g179364 (n_4191, n_3569, n_3840);
  nand g179363 (n_4190, n_3571, n_3839);
  nand g179362 (n_4189, n_649, n_3837);
  nand g179359 (n_4188, g1389, n_3826);
  nand g179358 (n_4187, g35, n_3729);
  nand g179355 (n_4186, g35, n_3776);
  nand g179354 (n_4185, g837, n_3827);
  not g179027 (n_4184, n_4183);
  nand g179350 (n_4180, g35, g311);
  nand g179047 (n_4179, n_2274, n_3698);
  nor g179052 (n_4178, n_3000, n_3778);
  fflopd g1319_reg(.CK (clock), .D (n_3696), .Q (g1319));
  nor g179057 (n_4177, n_3004, n_3781);
  nor g179060 (n_4176, n_3002, n_3783);
  nor g179062 (n_4175, n_4174, n_3597);
  nor g179063 (n_4173, n_4174, n_3469);
  nand g179068 (n_4172, n_2002, n_3851);
  nand g179070 (n_4171, n_3694, n_5126);
  nand g179073 (n_4170, n_3746, n_4922);
  nand g179074 (n_4169, n_3695, n_4168);
  nand g179075 (n_4167, g417, n_4133);
  nand g179076 (n_4166, n_3535, n_3838);
  nand g179082 (n_4165, n_3766, n_2536);
  nand g179083 (n_4164, n_3768, n_2539);
  nor g179088 (n_4163, g9680, n_3806);
  nor g179095 (n_4162, g9817, n_3816);
  nor g179102 (n_4161, g8277, n_3824);
  nand g179103 (n_4160, n_3771, n_3065);
  nand g179104 (n_4159, n_4492, n_3745);
  nor g179109 (n_4158, g8342, n_3820);
  nor g179113 (n_4157, g2047, n_3807);
  nor g179115 (n_4156, g8398, n_3815);
  nor g179121 (n_4155, g1978, n_3828);
  nor g179123 (n_4154, n_4153, n_4150);
  nor g179125 (n_4152, g9615, n_3805);
  nor g179127 (n_4151, g4664, n_4150);
  nor g179129 (n_4148, g2537, n_3818);
  nand g179131 (n_4147, g311, n_205);
  nor g179132 (n_4146, g9741, n_3829);
  nand g179133 (n_4145, n_1893, n_3741);
  nand g179136 (n_4144, n_4143, n_3747);
  nor g179142 (n_4142, n_1560, n_3975);
  nand g179159 (n_4141, g661, n_4140);
  nand g179160 (n_4139, g311, n_4138);
  nand g179349 (n_4137, g969, n_4081);
  nand g179341 (n_4136, n_661, n_3782);
  nand g179336 (n_4135, g14096, n_5795);
  nand g179329 (n_4134, n_4047, n_4133);
  nand g179322 (n_4132, n_1588, n_3750);
  nand g179321 (n_4131, n_3770, n_3526);
  nand g179320 (n_4130, g35, n_10212);
  nand g179315 (n_4129, g35, n_3756);
  nand g179313 (n_4128, g311, n_9257);
  wire w127, w128, w129, w130;
  nand g179305 (n_4127, w128, w130);
  nand g137 (w130, w129, g4991);
  not g136 (w129, n_3990);
  nand g135 (w128, w127, n_3990);
  not g134 (w127, g4991);
  nand g179303 (n_4126, n_2272, n_3708);
  nand g179302 (n_4125, n_2259, n_3722);
  nand g179301 (n_4124, n_2266, n_3716);
  nand g179299 (n_4123, n_2261, n_3730);
  nand g179298 (n_4122, n_2277, n_3706);
  not g179286 (n_4121, n_4438);
  not g179280 (n_4120, n_4407);
  not g179276 (n_4119, n_4409);
  not g179237 (n_4118, n_3890);
  not g179239 (n_4117, n_3891);
  not g179242 (n_4116, n_3892);
  not g179243 (n_4115, n_3893);
  not g179255 (n_4114, n_4098);
  not g179256 (n_4113, n_4096);
  not g179259 (n_4112, n_4095);
  not g179261 (n_4111, n_4091);
  not g179262 (n_4110, n_4090);
  not g179263 (n_4109, n_4086);
  not g179264 (n_4108, n_4085);
  not g179268 (n_4105, n_4078);
  not g179273 (n_4104, n_4417);
  not g179274 (n_4103, n_4411);
  not g179275 (n_4102, n_4393);
  nand g179225 (n_4286, g4871, n_3819);
  nand g179200 (n_4289, g6381, n_3785);
  nand g179195 (n_4809, g822, n_4101);
  nand g179455 (g31521, n_1956, n_3813);
  not g179040 (n_4656, g5069);
  nand g179162 (n_4379, g7946, n_3853);
  nor g179168 (n_4625, g4064, n_4056);
  nand g179171 (n_4377, g703, n_3700);
  fflopd g4369_reg(.CK (clock), .D (n_3717), .Q (g4369));
  nand g179174 (n_4375, g7916, n_3852);
  nand g179175 (n_4373, g671, n_4140);
  nand g179191 (n_4537, g4878, n_3831);
  nand g179179 (n_4522, g6035, n_3792);
  nand g179180 (n_4539, g4864, n_3823);
  nand g179182 (n_4525, g5689, n_3787);
  nand g179177 (n_4535, g4836, n_3809);
  nand g179183 (n_4523, g4040, n_3796);
  nand g179184 (n_4528, g6727, n_3790);
  nand g179185 (n_4526, g3338, n_3859);
  fflopd g881_reg(.CK (clock), .D (g14096), .Q (g14125));
  fflopd g86_reg(.CK (clock), .D (n_3857), .Q (g20557));
  fflopd g1495_reg(.CK (clock), .D (n_3726), .Q (g1495));
  fflopd g5517_reg(.CK (clock), .D (n_3672), .Q (g5517));
  fflopd g3161_reg(.CK (clock), .D (n_3669), .Q (g3161));
  fflopd g3512_reg(.CK (clock), .D (n_3668), .Q (g3512));
  fflopd g5863_reg(.CK (clock), .D (n_3666), .Q (g5863));
  fflopd g3863_reg(.CK (clock), .D (n_3667), .Q (g3863));
  nand g179571 (n_4100, n_1747, n_3985);
  nand g179387 (n_4099, n_3587, n_2460);
  nand g179401 (n_4098, g3550, g14451);
  nand g179407 (n_4097, g5901, g13068);
  nand g179408 (n_4096, g3889, g14518);
  nand g179415 (n_4095, g5889, g13068);
  nand g179416 (n_4094, g5208, g13039);
  nand g179418 (n_4093, g3901, g14518);
  nand g179419 (n_4092, new_g10354_, n_3978);
  nand g179422 (n_4091, g6235, g13085);
  nand g179424 (n_4090, g6247, g13085);
  nand g179425 (n_4089, g5555, g13049);
  nand g179427 (n_4088, n_3585, n_2018);
  nand g179430 (n_4087, n_1036, n_3583);
  nand g179433 (n_4086, n_931, n_3539);
  nand g179438 (n_4085, g5196, g13039);
  nand g179810 (n_4084, n_3344, n_3553);
  not g179797 (n_4083, n_4150);
  not g179794 (n_4082, n_4081);
  nand g179449 (n_4078, g35, g10306);
  not g179792 (n_4077, n_4076);
  not g179791 (n_4075, n_4074);
  not g179789 (n_4073, n_3709);
  nand g179456 (n_4072, n_3429, n_5660);
  nand g179457 (n_4071, n_3525, n_5660);
  not g179787 (n_4070, n_3710);
  not g179785 (n_4069, n_3711);
  not g179783 (n_4068, n_3713);
  not g179782 (n_4067, n_3715);
  not g179764 (n_4066, n_3731);
  not g179758 (n_4065, n_3797);
  not g179491 (n_4064, n_3821);
  not g179493 (n_4063, n_3802);
  not g179495 (n_4062, n_3800);
  not g179496 (n_4061, n_3777);
  not g179498 (n_4060, n_3765);
  not g179503 (n_4059, n_4058);
  not g179504 (n_4057, n_4056);
  not g179757 (n_4055, n_3848);
  not g179755 (n_4054, n_3760);
  not g179754 (n_4053, n_3757);
  not g179747 (n_4051, n_3744);
  nand g179522 (n_4050, n_3758, n_3407);
  nand g179534 (n_4049, g4643, n_3424);
  nand g179536 (n_4048, n_1897, n_4047);
  nand g179537 (n_4046, n_2843, n_4047);
  nand g179538 (n_4045, g246, n_4047);
  nand g179539 (n_4044, g269, n_4047);
  nand g179540 (n_4043, g446, n_4047);
  nand g179541 (n_4042, g854, n_4047);
  nand g179545 (n_4041, n_1906, n_3419);
  nand g179549 (n_4040, n_3084, n_3397);
  nand g179551 (n_4039, n_3062, n_3395);
  nand g179555 (n_4037, n_3033, n_3394);
  nor g179557 (n_4036, g4854, n_4018);
  nand g179558 (n_4035, g1384, n_3428);
  nand g179561 (n_4034, n_3060, n_3396);
  nand g179562 (n_4033, n_2824, n_3603);
  nand g179567 (n_4032, n_3056, n_3391);
  nand g179570 (n_4031, n_2310, n_3494);
  nand g179370 (n_4030, g3187, g14421);
  nand g179577 (n_4028, n_3049, n_3382);
  nand g179585 (n_4024, n_3085, n_3421);
  nand g179587 (n_4022, n_2775, n_3608);
  nand g179590 (n_4020, n_3916, n_3917);
  nor g179591 (n_4019, n_4017, n_4018);
  nand g179598 (n_4015, g9553, n_3521);
  nor g179609 (n_4014, n_4013, n_3992);
  nand g179612 (n_4012, n_1632, n_3987);
  nand g179614 (n_4011, g1585, n_4010);
  nor g179616 (n_4009, n_4008, n_3994);
  nand g179621 (n_4007, n_2187, n_3492);
  nand g179623 (n_4006, g1008, n_3489);
  nand g179627 (n_4005, g2638, n_7349);
  nand g179628 (n_4004, g2504, n_7351);
  nand g179631 (n_4003, g2079, n_7349);
  nand g179632 (n_4002, g1945, n_7351);
  nand g179644 (n_4001, g23683, n_4000);
  nand g179647 (n_3999, n_2263, n_3467);
  nand g179648 (n_3998, n_1916, n_3490);
  nand g179649 (n_3997, g1351, n_3610);
  nand g179661 (n_3996, n_1891, n_3861);
  nand g179665 (n_3995, n_4008, n_3994);
  nand g179666 (n_3993, n_4013, n_3992);
  nand g179711 (n_3991, g4966, n_3990);
  nand g179684 (n_3989, new_g6821_, n_3988);
  nand g179680 (n_4330, n_966, n_3987);
  nor g179686 (n_4363, n_1770, n_3944);
  nand g179690 (n_4243, g1199, n_3970);
  nand g179692 (n_4241, g1542, n_3904);
  nand g179445 (n_4106, n_3986, n_3876);
  nand g179706 (n_4238, n_1746, n_3985);
  nor g179446 (n_4469, n_9257, n_3981);
  nor g179447 (n_4473, n_9257, n_3976);
  nand g179678 (n_4423, g23683, n_3988);
  nor g179448 (n_4475, n_9257, n_3979);
  nand g179730 (n_4194, g4793, n_3508);
  nor g179450 (n_4483, n_9257, n_3980);
  nand g179677 (n_4246, n_2826, n_3987);
  nor g179451 (n_4455, n_9257, n_3977);
  not g179513 (n_4324, n_3984);
  not g179509 (n_4322, n_3983);
  not g179508 (n_4326, n_3982);
  nand g179452 (n_4400, g4064, n_3622);
  nand g179465 (n_4409, g35, n_3981);
  nand g179464 (n_4393, g35, n_3980);
  nand g179463 (n_4411, g35, n_3979);
  nand g179462 (n_4417, g35, n_3978);
  nand g179469 (n_4407, g35, n_3977);
  nand g179476 (n_4438, g35, n_3976);
  fflopd g351_reg(.CK (clock), .D (n_3393), .Q (g351));
  fflopd g2724_reg(.CK (clock), .D (n_3589), .Q (g2724));
  nand g179714 (n_4422, new_g12440_, n_3511);
  not g179799 (n_4320, n_3975);
  nand g179710 (n_4332, new_g6821_, n_4000);
  nand g179709 (n_4328, new_g6832_, n_4010);
  not g179521 (n_4358, n_4174);
  nand g179997 (n_3974, n_35, n_7349);
  nand g179816 (n_3973, g4104, n_9257);
  nand g179819 (n_3972, g736, n_9257);
  nand g179822 (n_3971, n_3969, n_3970);
  nor g179826 (n_3968, n_2813, n_3392);
  nand g179827 (n_3967, n_1260, n_3990);
  nand g179831 (n_3966, n_3497, n_3422);
  nand g179841 (n_3964, n_3462, n_3228);
  nand g179842 (n_3963, n_3006, n_3461);
  nand g179845 (n_3962, g4950, n_3643);
  nand g179847 (n_3961, n_1112, n_3480);
  nand g179850 (n_3960, n_3460, n_3223);
  nand g179852 (n_3959, n_3008, n_3448);
  nand g179855 (n_3958, g35, n_3860);
  nand g179858 (n_3957, g4939, n_3651);
  nand g179859 (n_3956, g1216, n_3389);
  nand g179861 (n_3955, n_3457, n_3168);
  nand g179862 (n_3954, n_3015, n_3474);
  nand g179864 (n_3953, n_3454, n_3207);
  nand g179865 (n_3952, n_2850, n_3453);
  nand g179866 (n_3951, g1300, n_3405);
  nand g179867 (n_3950, n_3447, n_3250);
  nand g179875 (n_3949, n_2998, n_3601);
  nand g179880 (n_3948, n_790, n_3481);
  nand g179881 (n_3947, n_1070, n_3486);
  nand g179885 (n_3946, n_3458, n_3249);
  nand g179888 (n_3945, g1554, n_3944);
  nand g179893 (n_3943, n_3446, n_3358);
  nand g179897 (n_3942, n_3443, n_3359);
  nand g179898 (n_3941, n_3010, n_3442);
  nand g179907 (n_3940, g1559, n_3390);
  nand g179908 (n_3939, n_970, n_3440);
  nand g179910 (n_3938, n_1291, n_3596);
  nand g179912 (n_3937, g504, n_3935);
  nand g179913 (n_3936, g513, n_3935);
  nand g179916 (n_3934, n_3438, n_3179);
  nand g179918 (n_3933, n_3441, n_3165);
  nand g179919 (n_3932, n_3014, n_3435);
  nand g179926 (n_3931, n_3450, n_3111);
  nand g179929 (n_3930, n_545, n_3432);
  nand g179931 (n_3929, n_3157, n_3515);
  nand g179933 (n_3928, n_3479, n_3153);
  nand g179935 (n_3927, n_3466, n_3152);
  nand g179936 (n_3926, n_3012, n_3468);
  nand g179938 (n_3925, n_710, n_3451);
  nand g179366 (n_3924, g3199, g14421);
  nand g179945 (n_3923, n_883, n_3471);
  nand g179950 (n_3922, n_3463, n_3136);
  nand g179953 (n_3921, g732, n_3920);
  nand g179955 (n_3919, n_1033, n_3594);
  nor g179963 (n_3918, n_3916, n_3917);
  nand g179966 (n_3915, g4749, n_3649);
  nand g179967 (n_3914, g4760, n_3647);
  nand g179968 (n_3913, g4771, n_3645);
  nand g179972 (n_3912, g4854, n_3399);
  nand g179974 (n_3911, g4961, n_3653);
  nand g179975 (n_3910, n_764, n_3482);
  nand g179976 (n_3909, g35, n_3465);
  nand g179981 (n_3908, g5033, n_3406);
  nand g179984 (n_3907, n_3599, n_3114);
  nand g179989 (n_3906, n_3592, n_3219);
  nand g179995 (n_3905, n_3903, n_3904);
  nand g179811 (n_3902, n_2867, n_3507);
  nand g179999 (n_3901, n_194, n_7351);
  nand g180003 (n_3900, n_83, n_7351);
  nand g180005 (n_3899, n_142, n_7349);
  nand g180010 (n_3898, n_2724, n_3513);
  nand g179361 (n_3897, g35, n_3625);
  nand g179360 (n_3896, g35, n_3850);
  nand g179357 (n_3895, n_584, n_3584);
  nand g179351 (n_3894, g6593, g13099);
  nand g179348 (n_3893, n_3588, n_1928);
  nand g179347 (n_3892, g6581, g13099);
  nand g179343 (n_3891, g5543, g13049);
  nand g179340 (n_3890, g3538, g14451);
  nand g179324 (n_3889, n_2157, n_3884);
  not g180378 (n_3888, n_3693);
  nor g179323 (n_3887, n_9257, n_3623);
  nand g179319 (n_3885, n_1561, n_3884);
  nor g179316 (n_3883, n_2295, n_3617);
  nor g179314 (n_3882, n_2297, n_3615);
  not g179795 (n_3881, n_3880);
  wire w131, w132, w133, w134;
  nand g179306 (n_3879, w132, w134);
  nand g141 (w134, w133, n_3739);
  not g140 (w133, n_3740);
  nand g139 (w132, w131, n_3740);
  not g138 (w131, n_3739);
  nand g179048 (n_3878, n_1950, n_3884);
  nand g179056 (n_3877, g4392, n_3876);
  nand g179065 (n_3875, n_2856, n_3884);
  nand g179067 (n_3874, n_3986, n_3618);
  nor g179069 (n_3873, n_3557, n_6159);
  nor g179071 (n_3872, n_3533, n_1410);
  nor g179072 (n_3871, n_3531, n_1540);
  nor g179078 (n_3870, n_3550, n_1545);
  nand g179086 (n_3869, n_163, n_3624);
  nand g179134 (n_3868, n_60, n_3621);
  nand g179153 (n_3867, n_3534, n_2953);
  not g179257 (n_3866, n_3856);
  fflopd g5069_reg(.CK (clock), .D (n_3537), .Q (g5069));
  fflopd g4423_reg(.CK (clock), .D (g10306), .Q (g4423));
  nand g180022 (n_4195, g35, n_3920);
  not g180049 (n_4477, n_3865);
  not g180050 (n_4425, n_3864);
  not g180054 (n_4427, n_3863);
  not g180055 (n_4426, n_3862);
  nand g179170 (n_4181, g269, n_3427);
  nor g179167 (n_4183, g269, n_3613);
  wire w135, w136, w137, w138;
  nand g178520 (n_4283, w136, w138);
  nand g147 (w138, w137, n_2304);
  not g145 (w137, n_3370);
  nand g144 (w136, w135, n_3370);
  not g143 (w135, n_2304);
  nor g179206 (n_4692, n_6582, n_3628);
  fflopd g1532_reg(.CK (clock), .D (n_3605), .Q (g1532));
  nor g179221 (n_4691, n_6562, n_3612);
  fflopd g1189_reg(.CK (clock), .D (n_3602), .Q (g1189));
  nand g180025 (n_5880, g35, n_3861);
  not g180053 (n_4480, n_3661);
  fflopd g862_reg(.CK (clock), .D (n_3488), .Q (g862));
  fflopd g1521_reg(.CK (clock), .D (n_3478), .Q (g1521));
  fflopd g4643_reg(.CK (clock), .D (n_3418), .Q (g4643));
  fflopd g1178_reg(.CK (clock), .D (n_3483), .Q (g1178));
  fflopd g5673_reg(.CK (clock), .D (g13049), .Q (g17813));
  fflopd g5327_reg(.CK (clock), .D (g13039), .Q (g17787));
  fflopd g6365_reg(.CK (clock), .D (g13085), .Q (g17845));
  fflopd g6711_reg(.CK (clock), .D (g13099), .Q (g17871));
  fflopd g3668_reg(.CK (clock), .D (g14451), .Q (g16924));
  fflopd g4019_reg(.CK (clock), .D (g14518), .Q (g16955));
  nand g180024 (n_4871, n_4457, n_3860);
  fflopd g3317_reg(.CK (clock), .D (g14421), .Q (g16874));
  fflopd g6019_reg(.CK (clock), .D (g13068), .Q (g17819));
  nand g180026 (n_9193, g35, new_g10233_);
  nor g179625 (n_3859, n_3858, n_4842);
  nand g179382 (n_3857, n_1977, n_3363);
  nand g179411 (n_3856, g699, n_3367);
  nand g179426 (n_3855, n_2029, n_3362);
  nand g179439 (n_3854, g35, n_3365);
  not g179492 (n_3853, n_3620);
  not g179494 (n_3852, n_3619);
  not g179506 (n_3851, n_3850);
  nand g179871 (n_3849, n_7031, n_3274);
  nand g179853 (n_3848, n_689, n_3266);
  nand g179523 (n_3847, g437, n_3845);
  nand g179524 (n_3846, g433, n_3845);
  nand g179525 (n_3844, g429, n_3845);
  nand g179526 (n_3843, g424, n_3845);
  nand g179527 (n_3842, g417, n_3845);
  nand g179528 (n_3841, g411, n_3845);
  nand g179529 (n_3840, g405, n_3845);
  nand g179530 (n_3839, g401, n_3845);
  nand g179531 (n_3838, n_2866, n_3241);
  nand g179532 (n_3837, g392, n_3845);
  nand g179533 (n_3836, g847, n_3845);
  nand g179535 (n_3835, n_3834, n_3775);
  nor g179542 (n_3833, n_3499, n_3278);
  nand g179543 (n_3832, g4392, n_3755);
  nand g179544 (n_3831, n_2311, n_3822);
  nor g179546 (n_3830, n_3504, n_3285);
  nor g179550 (n_3829, g6098, n_3331);
  nand g179553 (n_3828, n_227, n_3319);
  nor g179554 (n_3827, g812, n_3502);
  nand g179559 (n_3826, n_2312, n_3732);
  nor g179564 (n_3824, g3050, n_3328);
  nand g179565 (n_3823, n_2172, n_3822);
  nand g179566 (n_3821, n_3342, n_3067);
  nor g179568 (n_3820, g3401, n_3326);
  nand g179569 (n_3819, n_3493, n_3822);
  nand g179573 (n_3818, n_229, n_3318);
  nand g179574 (n_3817, n_2346, n_3811);
  nor g179575 (n_3816, g6444, n_3330);
  nor g179576 (n_3815, g3752, n_3325);
  nand g179580 (n_3814, g4098, n_3323);
  nand g179582 (n_3813, n_2870, n_3324);
  nand g179588 (n_3812, n_2315, n_3811);
  nand g179593 (n_3809, n_2348, n_3822);
  nand g179595 (n_3808, n_3491, n_3811);
  nand g179599 (n_3807, n_173, n_3317);
  nor g179600 (n_3806, g5752, n_3332);
  nor g179601 (n_3805, g5406, n_3316);
  nor g179606 (n_3804, n_3500, n_3293);
  nand g179608 (n_3803, g441, n_3845);
  nand g179611 (n_3802, g203, n_1347);
  nand g179618 (n_3801, n_1955, n_3737);
  nand g179619 (n_3800, n_3338, n_3068);
  nor g179622 (n_3799, n_3498, n_3292);
  nor g179624 (n_3798, n_3503, n_3294);
  nand g179860 (n_3797, n_605, n_3335);
  nor g179626 (n_3796, n_3795, n_896);
  nand g179629 (n_3794, g2370, n_7347);
  nand g179633 (n_3793, g1811, n_7347);
  nor g179635 (n_3792, n_3791, n_448);
  nor g179637 (n_3790, n_3788, n_3789);
  nor g179638 (n_3787, n_3786, n_892);
  nor g179639 (n_3785, n_3784, n_900);
  nor g179640 (n_3783, g16718, n_3300);
  nand g179641 (n_3782, g182, n_3779);
  nor g179642 (n_3781, g16775, n_3299);
  nand g179643 (n_3780, g174, n_3779);
  nor g179645 (n_3778, g17674, n_3297);
  nand g179646 (n_3777, n_2530, n_3286);
  nor g179650 (n_3776, g4793, n_3775);
  nand g179651 (n_3774, n_3246, n_3773);
  nand g179652 (n_3772, n_3064, n_5760);
  nand g179653 (n_3771, n_3245, n_5758);
  nand g179654 (n_3770, n_3244, n_3769);
  nand g179656 (n_3768, n_3242, n_3767);
  nand g179658 (n_3766, n_3063, n_6456);
  nand g179663 (n_3765, n_2695, n_3337);
  nand g179667 (n_3764, g452, n_3779);
  nand g179668 (n_3763, g460, n_3779);
  nand g179669 (n_3762, g168, n_3779);
  nand g179670 (n_3761, n_2188, n_3811);
  nand g179851 (n_3760, n_768, n_3232);
  nor g179687 (n_3759, n_3718, n_3758);
  nand g179849 (n_3757, n_490, n_3268);
  nor g179846 (n_3756, n_3986, n_3755);
  nand g179839 (n_3754, g14217, n_5795);
  nand g179835 (n_3753, g35, n_3238);
  nand g179833 (n_3752, g35, n_3243);
  nand g179832 (n_3751, g35, n_3240);
  nor g179825 (n_3750, n_2331, n_3356);
  nand g179818 (n_3749, g5112, n_9257);
  wire w139, w140, w141, w142;
  nand g179809 (n_3748, w140, w142);
  nand g152 (w142, w141, g4358);
  not g151 (w141, n_3379);
  nand g149 (w140, w139, n_3379);
  not g148 (w139, g4358);
  nand g179806 (n_3747, n_6019, n_3106);
  not g179777 (n_3746, n_3549);
  not g179780 (n_3745, n_3541);
  nand g179802 (n_3744, new_g8038_, n_3505);
  nand g179803 (n_3743, g699, n_3845);
  nand g179804 (n_3742, g703, n_3845);
  nand g179805 (n_3741, n_6011, n_3124);
  nor g179695 (n_4101, n_3739, n_3740);
  fflopd g2844_reg(.CK (clock), .D (n_3295), .Q (g2844));
  nand g179705 (n_3984, g12238, n_3279);
  nor g179685 (n_4058, n_2980, n_3159);
  nand g179696 (n_3983, g11349, n_3288);
  not g179510 (n_4133, n_3738);
  nand g179694 (n_3982, g11418, n_3281);
  nand g179689 (n_4056, g4057, n_3737);
  nand g179688 (n_9273, n_3736, n_3321);
  not g179519 (n_4140, n_3978);
  fflopd g878_reg(.CK (clock), .D (g14217), .Q (g14096));
  nand g179746 (n_4174, g4180, n_3368);
  fflopd g311_reg(.CK (clock), .D (n_3217), .Q (g311));
  nand g179914 (n_3735, g475, n_3845);
  nand g179874 (n_3734, n_595, n_3309);
  nand g179877 (n_3733, g1312, n_3732);
  nand g179879 (n_3731, n_796, n_3229);
  nand g179882 (n_3730, n_3275, n_2532);
  nand g179884 (n_3729, g1351, n_3307);
  nand g179889 (n_3728, n_2930, n_3304);
  nand g179899 (n_3727, n_2507, n_3360);
  nand g179900 (n_3726, n_2927, n_3301);
  nand g179909 (n_3725, g499, n_3186);
  nand g179911 (n_3724, n_7035, n_3271);
  nand g179921 (n_3723, g2236, n_7331);
  nand g179927 (n_3722, n_3276, n_2527);
  nand g179930 (n_3721, g1677, n_7331);
  nand g179939 (n_3720, g691, n_3194);
  nand g179947 (n_3719, g209, n_3718);
  nand g179956 (n_3717, n_323, n_3182);
  nand g179958 (n_3716, n_3277, n_2528);
  nand g179959 (n_3715, n_1126, n_3267);
  nand g179965 (n_3714, n_6888, n_3280);
  nand g179969 (n_3713, n_3736, n_3121);
  nand g179971 (n_3712, g969, n_3630);
  nand g179977 (n_3711, n_2639, n_3098);
  nand g179979 (n_3710, n_2641, n_3107);
  nand g179988 (n_3709, g1199, n_3501);
  nand g179991 (n_3708, n_3273, n_2526);
  nand g179992 (n_3707, n_6884, n_3291);
  nand g179993 (n_3706, n_3289, n_2531);
  nand g179998 (n_3705, n_220, n_7347);
  nand g180000 (n_3704, n_156, n_7331);
  nand g180001 (n_3703, n_5789, n_3284);
  nand g180002 (n_3702, n_166, n_7347);
  nand g180004 (n_3701, n_15, n_7331);
  nor g180007 (n_3700, g837, n_3372);
  nand g180008 (n_3699, n_6886, n_3351);
  nand g180009 (n_3698, n_3336, n_2529);
  nand g180011 (n_3697, n_3081, n_3845);
  nand g179872 (n_3696, n_2035, n_3260);
  not g179767 (n_3695, n_3568);
  not g179786 (n_3694, n_3532);
  nand g180611 (n_3693, new_g6961_, n_3071);
  nor g180604 (n_3692, n_3691, n_3631);
  nand g180429 (n_3690, n_1044, n_4854);
  nand g180428 (n_3689, g35, n_3044);
  nand g180422 (n_3688, g35, n_3055);
  not g180028 (n_3687, n_3609);
  not g180029 (n_3686, n_3611);
  not g180030 (n_3685, n_3485);
  not g180031 (n_3684, n_3484);
  not g180032 (n_3683, n_3475);
  not g180034 (n_3682, n_3452);
  not g180037 (n_3681, n_3434);
  not g180038 (n_3680, n_3433);
  not g180043 (n_3679, g736);
  not g180051 (n_3678, n_3860);
  not g180059 (n_3677, new_g10233_);
  nand g180080 (n_3675, n_1350, n_3032);
  nand g180103 (n_3674, n_1920, n_3022);
  nand g180138 (n_3673, g12184, n_3076);
  nand g180228 (n_3672, n_1709, n_3083);
  nand g180229 (n_3671, n_1727, n_3058);
  nand g180230 (n_3670, n_1726, n_3053);
  nand g180231 (n_3669, n_1708, n_3057);
  nand g180232 (n_3668, n_1711, n_3052);
  nand g180233 (n_3667, n_1716, n_3050);
  nand g180234 (n_3666, n_1723, n_3046);
  nand g180235 (n_3665, n_1713, n_3038);
  nand g180420 (n_3664, g35, n_3040);
  nand g180419 (n_3663, g35, n_3035);
  nand g180418 (n_3662, g35, n_3048);
  nand g180310 (n_3661, n_4225, n_3632);
  nand g180417 (n_3660, g35, n_3021);
  nand g180416 (n_3659, g35, n_3043);
  not g180361 (n_3658, n_3404);
  not g180373 (n_3656, n_3381);
  not g180374 (n_3655, n_3380);
  not g180384 (n_3654, n_3653);
  not g180385 (n_3652, n_3651);
  not g180386 (n_3650, n_3649);
  not g180389 (n_3648, n_3647);
  not g180390 (n_3646, n_3645);
  not g180391 (n_3644, n_3643);
  not g180395 (n_3642, n_4018);
  not g180397 (n_3641, n_3920);
  nand g180405 (n_3640, g35, n_3023);
  nand g180406 (n_3639, g35, n_3054);
  nand g180408 (n_3638, g35, n_3041);
  nand g180409 (n_3637, g35, n_3037);
  nand g180410 (n_3636, g35, n_3026);
  nand g180411 (n_3635, g35, n_3034);
  nand g180412 (n_3634, g35, n_3045);
  nand g180415 (n_3633, g35, n_3051);
  nand g180314 (n_3862, g5033, n_3079);
  nand g180311 (n_3863, n_4013, n_3632);
  nand g180307 (n_3864, n_4008, n_3632);
  nand g180306 (n_3865, g4311, n_3631);
  nor g180283 (n_4219, n_3378, n_3069);
  nand g180023 (n_3975, g979, n_3101);
  nand g180013 (n_4074, g35, n_3519);
  nand g180019 (n_3880, n_2200, n_3231);
  nand g180018 (n_4081, g35, n_3630);
  nand g180014 (n_4076, g35, n_3517);
  nand g180016 (n_4192, g35, n_3343);
  nand g180017 (n_4079, n_3408, n_3410);
  nand g180021 (n_4150, g35, n_3775);
  fflopd g4621_reg(.CK (clock), .D (n_3314), .Q (g4621));
  fflopd g1564_reg(.CK (clock), .D (n_3312), .Q (g1564));
  fflopd g4628_reg(.CK (clock), .D (n_3366), .Q (g4628));
  fflopd g4849_reg(.CK (clock), .D (n_3313), .Q (g4849));
  fflopd g4269_reg(.CK (clock), .D (n_3322), .Q (g4269));
  fflopd g5097_reg(.CK (clock), .D (n_3327), .Q (g5097));
  fflopd g1221_reg(.CK (clock), .D (n_3311), .Q (g1221));
  nand g179924 (n_3629, g3550, n_2989);
  nand g179634 (n_3628, g16656, n_3627);
  nand g180146 (n_3626, g1216, n_3472);
  nand g179547 (n_3625, n_3496, n_2841);
  nor g179556 (n_3624, g2491, n_2995);
  nor g179563 (n_3623, g2932, g2999);
  nor g179581 (n_3622, g4057, n_3198);
  nor g179583 (n_3621, g8788, n_2993);
  nand g179610 (n_3620, n_2547, n_2934);
  nand g179613 (n_3619, n_2545, n_2827);
  nor g179615 (n_3618, n_1694, n_3538);
  nor g179657 (n_3617, n_2893, n_3616);
  nor g179659 (n_3615, n_2891, n_3614);
  nand g179662 (n_3613, g246, n_2887);
  nand g179671 (n_3612, g17577, g25114);
  nand g180144 (n_3611, g5849, n_3593);
  nor g180142 (n_3610, n_3122, n_2818);
  nand g180140 (n_3609, g5156, n_3595);
  nor g180137 (n_3608, n_568, n_2865);
  nand g180132 (n_3606, g1559, n_3476);
  nand g180131 (n_3605, n_1961, n_2836);
  nor g180130 (n_3604, n_2607, n_2789);
  nor g180128 (n_3603, n_1822, n_3425);
  nand g180124 (n_3602, n_1960, n_2834);
  nand g180121 (n_3601, g6537, n_3598);
  nand g180120 (n_3599, g6533, n_3598);
  nand g180119 (n_3597, g6541, n_3598);
  nand g180118 (n_3596, g5272, n_3595);
  nand g180117 (n_3594, g5965, n_3593);
  nand g180116 (n_3592, g5467, n_3590);
  nand g180115 (n_3591, g5475, n_3590);
  not g180027 (n_3589, n_3347);
  nand g179814 (n_3588, new_g6821_, n_9257);
  nand g179815 (n_3587, new_g6832_, n_9257);
  nand g179817 (n_3586, g2946, n_9257);
  nand g179820 (n_3585, new_g8703_, n_9257);
  nand g179824 (n_3584, g35, n_2932);
  nand g179829 (n_3583, g35, n_2919);
  nand g179837 (n_3582, g35, n_2981);
  nand g179840 (n_3581, g182, n_3562);
  nand g179843 (n_3580, g5547, n_2917);
  nand g179844 (n_3579, g5555, n_2951);
  nand g179854 (n_3578, g5893, n_2938);
  nand g179856 (n_3577, g5901, n_2901);
  nand g179857 (n_3576, g5909, n_2896);
  nand g179868 (n_3575, g6247, n_2940);
  nand g179869 (n_3574, g6255, n_2943);
  nand g179870 (n_3573, g5563, n_2949);
  nand g179876 (n_3572, g6593, n_2935);
  nand g179886 (n_3571, g429, n_3570);
  nand g179887 (n_3569, g392, n_3570);
  nand g179890 (n_3568, g3203, g16624);
  nand g179891 (n_3567, g411, n_3570);
  nand g179892 (n_3566, g433, n_3570);
  nand g179894 (n_3565, g441, n_3570);
  nand g179896 (n_3564, g475, n_3570);
  nand g179901 (n_3563, g460, n_3562);
  nand g179902 (n_3561, g3187, n_2926);
  nand g179903 (n_3560, g3191, n_2925);
  nand g179904 (n_3559, g3199, n_2923);
  nand g179906 (n_3558, g3207, n_2922);
  nand g179915 (n_3557, g3554, g16656);
  nand g179920 (n_3556, g854, n_3570);
  nand g179922 (n_3555, g3538, n_2990);
  nand g179923 (n_3554, g3542, n_2912);
  nand g180102 (n_3553, g504, n_3523);
  nand g179925 (n_3552, g3558, n_2915);
  nand g179928 (n_3551, g6581, n_2987);
  nand g179932 (n_3550, g3905, g16693);
  nand g179937 (n_3549, g5212, g17577);
  nand g179940 (n_3548, g3889, n_2986);
  nand g179941 (n_3547, g3893, n_2911);
  nand g179942 (n_3546, g3909, n_2909);
  nand g179943 (n_3545, g5543, n_2992);
  nand g179944 (n_3544, g6235, n_2985);
  nand g179946 (n_3543, g6601, n_2948);
  nand g179949 (n_3542, g6585, n_2945);
  nand g179951 (n_3541, g6251, g17685);
  nand g179954 (n_3540, g6239, n_2941);
  nand g179957 (n_3539, n_2749, n_3538);
  nand g179960 (n_3537, n_630, n_2889);
  nand g179961 (n_3536, g5196, n_2984);
  nand g179962 (n_3535, g4628, n_2839);
  nand g179964 (n_3534, g4653, n_2899);
  nand g179970 (n_3533, g5905, g17646);
  nand g179978 (n_3532, g6597, g17722);
  nand g179980 (n_3531, g5559, g17604);
  nand g179982 (n_3530, g5889, n_2991);
  nand g179985 (n_3529, g5200, n_2890);
  nand g179986 (n_3528, g5208, n_2946);
  nand g179987 (n_3527, g5216, n_2955);
  nor g179994 (n_3526, n_2326, n_2997);
  nor g179996 (n_3525, g1135, new_g6821_);
  nand g180101 (n_3524, g513, n_3523);
  not g180039 (n_3521, g5112);
  nand g180100 (n_3516, g518, n_3523);
  nand g180098 (n_3515, g667, n_3523);
  nand g180097 (n_3514, g686, n_3523);
  nand g180092 (n_3513, n_3512, n_2830);
  nor g180086 (n_3511, n_3509, n_3510);
  not g180058 (n_3508, n_3775);
  nor g180081 (n_3507, n_2000, n_3423);
  fflopd g4104_reg(.CK (clock), .D (n_2963), .Q (g4104));
  not g180056 (n_3904, n_3506);
  not g180052 (n_3985, n_3505);
  nand g179673 (n_3977, g16627, n_3504);
  nand g179674 (n_3981, g17580, n_3503);
  not g180044 (n_3917, n_3502);
  nor g180015 (n_3876, n_9257, n_3538);
  not g180057 (n_3970, n_3501);
  nand g179675 (n_3976, g17607, n_3500);
  nand g179676 (n_3980, g17688, n_3499);
  nand g179683 (n_3979, g17649, n_3498);
  nand g179700 (n_3738, n_1911, n_3016);
  nor g179691 (n_3850, g1322, n_2936);
  nand g179742 (n_3978, n_3497, n_2983);
  not g180065 (n_3987, n_3630);
  not g180048 (n_3988, n_3255);
  not g180047 (n_4000, n_3257);
  nor g179719 (n_3884, n_3496, n_2982);
  fflopd g6000_reg(.CK (clock), .D (g17646), .Q (g13068));
  fflopd g6346_reg(.CK (clock), .D (g17685), .Q (g13085));
  fflopd g6692_reg(.CK (clock), .D (g17722), .Q (g13099));
  fflopd g5654_reg(.CK (clock), .D (g17604), .Q (g13049));
  fflopd g5308_reg(.CK (clock), .D (g17577), .Q (g13039));
  fflopd g3649_reg(.CK (clock), .D (g16656), .Q (g14451));
  fflopd g3298_reg(.CK (clock), .D (g16624), .Q (g14421));
  fflopd g4000_reg(.CK (clock), .D (g16693), .Q (g14518));
  fflopd g3873_reg(.CK (clock), .D (n_2783), .Q (g3873));
  nor g180149 (n_3494, n_3493, n_2746);
  nor g180152 (n_3492, n_3491, n_2794);
  nand g180153 (n_3490, g9497, n_2874);
  nor g180154 (n_3489, n_3104, n_2822);
  nand g180159 (n_3488, n_1985, n_2880);
  nand g180160 (n_3487, n_10218, n_3403);
  nand g180169 (n_3486, n_2313, n_3375);
  nand g180177 (n_3485, n_1330, n_2853);
  nand g180178 (n_3484, n_1242, n_2857);
  nand g180180 (n_3483, n_2181, n_2882);
  nand g180181 (n_3482, n_2567, n_2852);
  nand g180184 (n_3481, g6657, n_3598);
  nand g180185 (n_3480, g5619, n_3590);
  nand g180186 (n_3479, g3813, n_3470);
  nand g180189 (n_3478, n_2185, n_2832);
  nand g180190 (n_3477, g1554, n_3476);
  nand g180191 (n_3475, g3147, n_3445);
  nand g180192 (n_3474, g5152, n_3595);
  nand g180193 (n_3473, g1211, n_3472);
  nand g180215 (n_3471, g3965, n_3470);
  nand g180220 (n_3469, g6195, n_3456);
  nand g180226 (n_3468, g3845, n_3470);
  nand g180236 (n_3467, n_2525, n_2848);
  nand g180237 (n_3466, g3841, n_3470);
  nor g180239 (n_3465, g4983, n_3374);
  nand g180240 (n_3464, g3821, n_3470);
  nand g180241 (n_3463, g5120, n_3595);
  nand g180242 (n_3462, g5495, n_3590);
  nand g180243 (n_3461, g5499, n_3590);
  nand g180247 (n_3460, g5813, n_3593);
  nand g180248 (n_3459, g5821, n_3593);
  nand g180249 (n_3458, g5841, n_3593);
  nand g180251 (n_3457, g6159, n_3456);
  nand g180252 (n_3455, g6167, n_3456);
  nand g180253 (n_3454, g6187, n_3456);
  nand g180254 (n_3453, g6191, n_3456);
  nand g180255 (n_3452, g5503, n_3590);
  nand g180256 (n_3451, g6311, n_3456);
  nand g180257 (n_3450, g6505, n_3598);
  nand g180258 (n_3449, g5128, n_3595);
  nand g180261 (n_3448, g5845, n_3593);
  nand g180263 (n_3447, g5148, n_3595);
  nand g180264 (n_3446, g3111, n_3445);
  nand g180265 (n_3444, g3119, n_3445);
  nand g180266 (n_3443, g3139, n_3445);
  nand g180268 (n_3442, g3143, n_3445);
  nand g180269 (n_3441, g3490, n_3437);
  nand g180270 (n_3440, g3263, n_3445);
  nand g180271 (n_3439, g6513, n_3598);
  nand g180272 (n_3438, g3462, n_3437);
  nand g180273 (n_3436, g3470, n_3437);
  nand g180274 (n_3435, g3494, n_3437);
  nand g180275 (n_3434, g3498, n_3437);
  nand g180276 (n_3433, g3849, n_3470);
  nand g180277 (n_3432, g3614, n_3437);
  nand g179878 (n_3431, g3901, n_2838);
  nand g179883 (n_3430, g174, n_3562);
  nor g179948 (n_3429, g1129, new_g6821_);
  not g180393 (n_3428, n_3732);
  nor g180012 (n_3427, g246, n_2979);
  nand g180135 (g28041, n_3425, n_2825);
  nor g180670 (n_3424, g4340, n_3423);
  nor g180668 (n_3422, g817, n_3017);
  nand g180654 (n_3421, g35, n_2735);
  not g180363 (n_3419, n_3353);
  nand g180147 (n_3418, n_941, n_2868);
  not g180375 (n_3415, n_3133);
  not g180392 (n_3407, n_3718);
  nand g180648 (n_3406, g35, n_2755);
  nand g180610 (n_3405, n_2929, n_2774);
  nand g180413 (n_3404, n_3387, n_3403);
  nand g180423 (n_3402, g35, n_2829);
  nand g180424 (n_3401, g35, n_2883);
  nand g180425 (n_3400, g35, n_2801);
  nand g180426 (n_3399, g35, n_2970);
  nand g180427 (n_3398, g35, n_2833);
  nand g180433 (n_3397, g35, n_2958);
  nand g180448 (n_3396, g35, n_2762);
  nand g180462 (n_3395, g35, n_2812);
  nand g180480 (n_3394, g35, n_2740);
  nand g180491 (n_3393, n_1633, n_2966);
  nand g180507 (n_3392, n_2203, n_10222);
  nand g180511 (n_3391, g35, n_2797);
  nand g180523 (n_3390, g35, n_10220);
  nand g180539 (n_3389, g35, n_3031);
  nand g180550 (n_3386, g3562, n_2972);
  nand g180555 (n_3385, g3574, n_2859);
  nand g180561 (n_3384, g3590, n_2860);
  nand g180566 (n_3383, g3606, n_2858);
  nand g180578 (n_3382, g35, n_2767);
  nand g180601 (n_3381, n_2400, n_2730);
  nand g180605 (n_3380, g4349, n_3379);
  fflopd g546_reg(.CK (clock), .D (n_2861), .Q (g546));
  nor g180281 (n_3992, n_3378, n_2851);
  not g180394 (n_3861, n_3377);
  nand g180671 (n_3653, g35, n_2820);
  nand g180672 (n_3651, g35, n_3024);
  nand g180673 (n_3649, g35, n_3027);
  nand g180675 (n_3935, g35, n_2976);
  nand g180679 (n_3647, g35, n_3077);
  nand g180680 (n_3645, g35, n_2873);
  nand g180681 (n_3643, g35, n_3376);
  fflopd g736_reg(.CK (clock), .D (g11678), .Q (g736));
  nand g180287 (n_3944, n_2933, n_3375);
  nor g180282 (n_3994, n_3378, n_2847);
  nor g180308 (n_3860, g5033, n_2968);
  fflopd g4537_reg(.CK (clock), .D (n_2994), .Q (g10306));
  nand g180685 (n_4018, g35, n_3374);
  nor g180317 (n_4010, g1300, n_3018);
  nor g180319 (n_3990, n_998, n_3374);
  fflopd g4653_reg(.CK (clock), .D (n_2921), .Q (g4653));
  fflopd g4581_reg(.CK (clock), .D (n_2745), .Q (new_g10233_));
  nand g180687 (n_3920, n_2879, n_3305);
  fflopd g3522_reg(.CK (clock), .D (n_2778), .Q (g3522));
  fflopd g5873_reg(.CK (clock), .D (n_2809), .Q (g5873));
  fflopd g6219_reg(.CK (clock), .D (n_2808), .Q (g6219));
  fflopd g5180_reg(.CK (clock), .D (n_2956), .Q (g5180));
  fflopd g6565_reg(.CK (clock), .D (n_2725), .Q (g6565));
  fflopd g5527_reg(.CK (clock), .D (n_2960), .Q (g5527));
  fflopd g3171_reg(.CK (clock), .D (n_2791), .Q (g3171));
  nor g180343 (n_7351, new_g7717_, n_3373);
  fflopd g5092_reg(.CK (clock), .D (n_2729), .Q (g5092));
  nor g180688 (n_7349, n_3373, n_3197);
  not g180398 (n_4047, n_3372);
  nand g180238 (n_3371, n_2513, n_4988);
  wire w143, w144, w145, w146;
  nand g179444 (n_3370, w144, w146);
  nand g158 (w146, w145, g269);
  not g156 (w145, n_2303);
  nand g155 (w144, w143, n_2303);
  not g154 (w143, g269);
  nand g180514 (n_3369, g3195, n_2483);
  not g180041 (n_3368, new_g8703_);
  nor g179607 (n_3367, g650, n_2702);
  nand g179807 (n_3366, n_930, n_2707);
  wire w147, w148, w149, w150;
  nand g179821 (n_3365, w148, w150);
  nand g163 (w150, w149, g4527);
  not g162 (w149, n_3364);
  nand g161 (w148, w147, n_3364);
  not g159 (w147, g4527);
  nand g179905 (n_3363, g5097, n_2697);
  nand g179952 (n_3362, g4269, n_2696);
  nand g180509 (n_3360, g1489, n_2568);
  nand g180508 (n_3359, g3133, n_3357);
  nand g180506 (n_3358, g3147, n_3357);
  nand g180502 (n_3356, n_273, n_2654);
  not g180064 (n_3355, g16656);
  nand g180500 (n_3354, n_250, n_2653);
  nand g180498 (n_3353, n_1976, n_2496);
  not g180069 (n_3352, g17577);
  nor g180070 (n_3351, n_3296, n_2275);
  nand g180072 (n_3350, g6148, n_9257);
  nand g180073 (n_3349, g3451, n_9257);
  nand g180074 (n_3348, g3100, n_9257);
  nand g180075 (n_3347, new_g7753_, n_9257);
  nand g180076 (n_3346, g5802, n_9257);
  nand g180077 (n_3345, g4455, n_9257);
  nand g180082 (n_3344, n_1464, n_6177);
  nand g180083 (n_3343, n_606, n_5660);
  nand g180104 (n_3342, n_2509, n_4952);
  nand g180106 (n_3341, n_2515, n_5128);
  nand g180107 (n_3340, n_2512, n_5130);
  nand g180108 (n_3339, n_2367, n_4922);
  nand g180109 (n_3338, n_2511, n_4168);
  nand g180110 (n_3337, n_1909, n_10393);
  nand g180111 (n_3336, n_2369, g25114);
  nand g180112 (n_3335, g269, n_3333);
  nand g180113 (n_3334, g246, n_3333);
  fflopd g203_reg(.CK (clock), .D (n_2402), .Q (g203));
  nor g180122 (n_3332, g5802, n_2180);
  nor g180125 (n_3331, g6148, n_2168);
  nor g180126 (n_3330, g6494, n_2175);
  nor g180129 (n_3328, g3100, n_2320);
  nand g180133 (n_3327, n_2281, n_2364);
  nor g180134 (n_3326, g3451, n_2179);
  nor g180139 (n_3325, g3802, n_2173);
  nor g180141 (n_3324, g4087, n_2556);
  nor g180143 (n_3323, n_620, n_2554);
  nand g180145 (n_3322, n_2286, n_2669);
  nor g180150 (n_3321, n_3320, n_2877);
  nor g180151 (n_3319, g1710, n_10397);
  nor g180155 (n_3318, g2269, n_10387);
  nor g180157 (n_3317, g1913, n_10389);
  nor g180158 (n_3316, g5456, n_2178);
  nand g180161 (n_3315, n_1823, n_6177);
  nand g180163 (n_3314, n_2128, n_2685);
  nand g180164 (n_3313, n_2386, n_2661);
  nand g180165 (n_3312, n_2467, n_2656);
  nand g180166 (n_3311, n_2401, n_2657);
  nand g180170 (n_3310, n_384, n_2549);
  nand g180176 (n_3309, n_3308, n_2424);
  nor g180182 (n_3307, g1389, n_3130);
  nand g180188 (n_3306, n_1149, n_3305);
  nand g180196 (n_3304, g1442, n_3302);
  nand g180197 (n_3303, g1484, n_3302);
  nand g180198 (n_3301, g1495, n_3302);
  nand g180199 (n_3300, n_3290, n_1517);
  nand g180200 (n_3299, n_3283, n_1595);
  nand g180202 (n_3297, n_3296, n_1594);
  nand g180495 (n_3295, n_387, n_2651);
  nor g180203 (n_3294, g17580, n_2541);
  nor g180204 (n_3293, g17607, n_2542);
  nor g180205 (n_3292, g17649, n_2543);
  nor g180206 (n_3291, n_3290, n_2278);
  nand g180207 (n_3289, n_2508, n_1945);
  nor g180209 (n_3288, n_3290, n_3001);
  nand g180210 (n_3287, n_2361, n_3627);
  nand g180211 (n_3286, g16627, n_2352);
  nor g180212 (n_3285, g16627, n_2540);
  nor g180213 (n_3284, n_3283, n_2264);
  nand g180214 (n_3282, g17649, n_2363);
  nor g180216 (n_3281, n_3283, n_3003);
  nor g180217 (n_3280, n_2686, n_2267);
  nor g180218 (n_3279, n_3296, n_2999);
  nor g180219 (n_3278, g17688, n_2368);
  nand g180221 (n_3277, n_2365, n_5152);
  nand g180222 (n_3276, n_2514, n_5150);
  nand g180223 (n_3275, n_2366, n_5148);
  nor g180224 (n_3274, n_2362, n_2273);
  nand g180225 (n_3273, n_2692, n_3272);
  nor g180227 (n_3271, n_2684, n_2262);
  nand g180494 (n_3270, g6649, n_2412);
  nand g180244 (n_3269, g225, n_3333);
  nand g180245 (n_3268, g232, n_3333);
  nand g180246 (n_3267, g239, n_3333);
  nand g180250 (n_3266, g262, n_3333);
  nand g180259 (n_3265, n_1908, n_2484);
  nand g180260 (n_3264, g255, n_3333);
  nand g180267 (n_3263, g446, n_3333);
  nand g180493 (n_3262, g5575, n_2489);
  nand g180492 (n_3261, g6613, n_2711);
  nand g180489 (n_3260, g35, n_2418);
  nand g180488 (n_3259, g6629, n_2574);
  nand g180487 (n_3258, g6625, n_2571);
  nand g180304 (n_3257, n_3256, n_5660);
  nand g180305 (n_3255, n_8069, n_5660);
  nand g180485 (n_3254, g6617, n_2408);
  nand g180484 (n_3253, g6605, n_2599);
  nand g180483 (n_3252, g6633, n_2398);
  nand g180482 (n_3251, g6589, n_2618);
  nand g180481 (n_3250, g5142, n_3135);
  nand g180479 (n_3249, g5835, n_3222);
  nand g180478 (n_3248, g6621, n_2391);
  nand g180476 (n_3247, g6299, n_2417);
  not g180364 (n_3246, n_2928);
  not g180368 (n_3245, n_2913);
  not g180370 (n_3244, n_2908);
  not g180371 (n_3243, n_2907);
  not g180377 (n_3242, n_2904);
  not g180379 (n_3241, n_2900);
  not g180380 (n_3240, n_2898);
  nand g180475 (n_3239, g6295, n_2713);
  nor g180474 (n_3238, n_3237, n_6019);
  nand g180473 (n_3236, g6287, n_2395);
  nand g180402 (n_3235, g6494, n_9257);
  nand g180403 (n_3234, g5109, n_9257);
  nand g180404 (n_3233, g5456, n_9257);
  nand g180407 (n_3232, g35, n_2374);
  nor g180414 (n_3231, n_2814, n_3230);
  nand g180431 (n_3229, g14201, n_5795);
  nand g180432 (n_3228, g5489, n_3218);
  nand g180434 (n_3227, g5925, n_2399);
  nand g180437 (n_3226, g5571, n_2583);
  nand g180438 (n_3225, g5587, n_2552);
  nand g180439 (n_3224, g5252, n_2678);
  nand g180440 (n_3223, g5849, n_3222);
  nand g180441 (n_3221, g5607, n_2694);
  nand g180442 (n_3220, g6279, n_2577);
  nand g180443 (n_3219, g5503, n_3218);
  nand g180444 (n_3217, n_346, n_2655);
  nand g180445 (n_3216, g5204, n_2630);
  nand g180446 (n_3215, g5611, n_2390);
  nand g180449 (n_3214, g6259, n_2459);
  nand g180450 (n_3213, g5917, n_2562);
  nand g180451 (n_3212, g5921, n_2706);
  nand g180452 (n_3211, g3929, n_2523);
  nand g180454 (n_3210, g5941, n_2425);
  nand g180455 (n_3209, g5949, n_2563);
  nand g180456 (n_3208, g5953, n_2393);
  nand g180459 (n_3207, g6181, n_3167);
  nand g180460 (n_3206, g3917, n_2558);
  nand g180465 (n_3205, g6243, n_2616);
  nand g180467 (n_3204, g5583, n_2481);
  nand g180468 (n_3203, g6263, n_2569);
  nand g180469 (n_3202, n_2589, n_2430);
  nand g180470 (n_3201, g6267, n_2383);
  nand g180471 (n_3200, g6271, n_2454);
  nand g180472 (n_3199, g6275, n_2415);
  nand g180300 (n_3502, g847, n_3497);
  not g180046 (n_3737, n_3198);
  not g180060 (n_3795, g16693);
  not g180061 (n_3784, g17685);
  not g180062 (n_3786, g17604);
  not g180063 (n_3858, g16624);
  not g180066 (n_3788, g17722);
  not g180068 (n_3755, n_3538);
  nand g180316 (n_3501, g7916, n_2546);
  nand g180315 (n_3506, g7946, n_2548);
  nand g180309 (n_3505, g518, n_2397);
  nand g180302 (n_3740, g817, n_3497);
  not g180067 (n_3791, g17646);
  nand g180294 (n_3517, g4975, n_2645);
  nand g180288 (n_3519, g4785, n_2647);
  fflopd g5112_reg(.CK (clock), .D (g9553), .Q (g5112));
  nand g180336 (n_3630, n_2642, n_6019);
  nor g180321 (n_3811, n_2290, n_2591);
  not g180396 (n_3822, n_2886);
  nand g180322 (n_3775, g4669, n_3834);
  not g180399 (n_3779, n_3562);
  fflopd g5176_reg(.CK (clock), .D (n_2380), .Q (new_g7704_));
  nor g180342 (n_7347, new_g7753_, n_3197);
  fflopd g6561_reg(.CK (clock), .D (n_2703), .Q (new_g7812_));
  not g180400 (n_3845, n_3570);
  nand g180519 (n_3196, g3215, n_2379);
  nand g180521 (n_3195, g3223, n_2472);
  nand g180522 (n_3194, n_1978, n_3185);
  nand g180524 (n_3193, g3231, n_2470);
  nand g180525 (n_3192, g3235, n_2469);
  nand g180526 (n_3191, g3239, n_2392);
  nand g180527 (n_3190, g3243, n_2466);
  nand g180528 (n_3189, g3247, n_2464);
  nand g180529 (n_3188, g3251, n_2463);
  nand g180530 (n_3187, g3255, n_2461);
  nand g180533 (n_3186, n_1348, n_3185);
  nand g180534 (n_3184, g499, n_3185);
  nand g180535 (n_3183, n_2165, n_2535);
  nand g180536 (n_3182, g4459, n_9257);
  nand g180538 (n_3181, g3802, n_9257);
  nand g180541 (n_3180, g5913, n_2360);
  nand g180545 (n_3179, g3498, n_3164);
  nand g180546 (n_3178, g5929, n_2437);
  nand g180547 (n_3177, g5897, n_2635);
  nand g180548 (n_3176, g3546, n_2633);
  nand g180551 (n_3175, g3566, n_2566);
  nand g180552 (n_3174, g35, n_2594);
  nand g180553 (n_3173, g3953, n_2426);
  nand g180554 (n_3172, g3570, n_2491);
  nand g180556 (n_3171, g6291, n_2420);
  nand g180557 (n_3170, g3578, n_2683);
  nand g180558 (n_3169, g3582, n_2565);
  nand g180559 (n_3168, g6195, n_3167);
  nand g180560 (n_3166, g3586, n_2443);
  nand g180562 (n_3165, g3484, n_3164);
  nand g180563 (n_3163, g3594, n_2442);
  nand g180564 (n_3162, g3598, n_2560);
  nand g180565 (n_3161, g3602, n_2406);
  nand g180568 (n_3160, g5957, n_2446);
  nand g180569 (n_3159, n_1907, n_2377);
  nand g180570 (n_3158, g5599, n_2389);
  nand g180571 (n_3157, g686, n_3185);
  nand g180572 (n_3156, g5551, n_2625);
  nand g180573 (n_3155, g35, n_3019);
  nand g180574 (n_3154, g3227, n_2441);
  nand g180576 (n_3153, g3849, n_3151);
  nand g180577 (n_3152, g3835, n_3151);
  nand g180518 (n_3150, g3211, n_2477);
  nand g180579 (n_3149, g5232, n_2680);
  nand g180582 (n_3148, g3897, n_2628);
  nand g180583 (n_3147, n_2592, n_2487);
  nand g180585 (n_3146, g3913, n_2691);
  nand g180586 (n_3145, g3921, n_2428);
  nand g180587 (n_3144, g3925, n_2521);
  nand g180589 (n_3143, g3933, n_2579);
  nand g180590 (n_3142, g3937, n_2671);
  nand g180592 (n_3141, g3941, n_2427);
  nand g180594 (n_3140, g3945, n_2668);
  nand g180595 (n_3139, g3949, n_2557);
  nand g180596 (n_3138, g3957, n_2500);
  nand g180598 (n_3137, n_2271, n_2604);
  nand g180600 (n_3136, g5156, n_3135);
  nand g180603 (n_3134, g6637, n_2414);
  nand g180606 (n_3133, n_2584, n_2422);
  nand g180607 (n_3132, n_2265, n_2603);
  nand g180609 (n_3131, g1312, n_3130);
  nand g180612 (n_3129, n_2640, n_2519);
  nand g180613 (n_3128, g5579, n_2674);
  nand g180614 (n_3127, g5595, n_2404);
  nand g180616 (n_3126, g6641, n_2551);
  nand g180619 (n_3125, g6609, n_2576);
  nand g180623 (n_3124, n_3122, n_3123);
  nand g180626 (n_3121, n_2016, n_2595);
  nand g180627 (n_3120, g5937, n_2405);
  nand g180630 (n_3119, g5260, n_2385);
  nand g180631 (n_3118, n_2449, n_259);
  nand g180633 (n_3117, g5603, n_2581);
  nand g180634 (n_3116, n_2268, n_2605);
  nand g180635 (n_3115, g6303, n_2407);
  nand g180638 (n_3114, g6527, n_3110);
  nand g180639 (n_3113, g6283, n_2495);
  nand g180640 (n_3112, n_2394, n_275);
  nand g180641 (n_3111, g6541, n_3110);
  nand g180642 (n_3109, g35, g4459);
  nand g180643 (n_3108, g5264, n_2378);
  nand g180644 (n_3107, g1008, n_2643);
  nand g180645 (n_3106, n_3104, n_3105);
  nand g180646 (n_3103, n_2638, n_2517);
  nand g180647 (n_3102, g5220, n_2498);
  nor g180649 (n_3101, g1221, n_2456);
  nand g180650 (n_3100, g5567, n_2672);
  nand g180652 (n_3099, g5933, n_2578);
  nand g180653 (n_3098, g1351, n_2637);
  nand g180655 (n_3097, g5591, n_2388);
  nand g180656 (n_3096, g5224, n_2573);
  nand g180657 (n_3095, g5228, n_2371);
  nand g180658 (n_3094, n_2269, n_2588);
  nand g180659 (n_3093, g5236, n_2447);
  nand g180660 (n_3092, g5240, n_2550);
  nand g180661 (n_3091, g5244, n_2700);
  nand g180662 (n_3090, g5248, n_2689);
  nand g180663 (n_3089, g5256, n_2555);
  nand g180664 (n_3088, g5945, n_2435);
  nand g180666 (n_3087, g35, n_2602);
  nand g180667 (n_3086, g6645, n_2410);
  not g180696 (n_3085, n_2885);
  not g180699 (n_3084, n_2959);
  not g180700 (n_3083, n_2961);
  not g180704 (n_3081, n_2855);
  not g180708 (n_3079, n_2844);
  not g180716 (n_3076, g11678);
  not g180702 (g21727, n_2967);
  nand g180790 (n_3074, g12238, n_2349);
  nand g180793 (n_3073, g11349, n_2350);
  nand g180803 (n_3072, g12422, n_2704);
  nand g180807 (n_3071, g4643, n_2357);
  nand g180826 (n_3070, g4253, n_2358);
  nand g180839 (n_3069, g1454, n_6441);
  nand g180889 (n_3068, g13895, n_2356);
  nand g180890 (n_3067, g13926, n_2354);
  nand g180891 (n_3066, g16775, n_2351);
  nand g180896 (n_3065, g13966, n_2355);
  not g180366 (n_3064, n_2918);
  not g180381 (n_3063, n_2892);
  not g181031 (n_3062, n_2807);
  not g181033 (n_3060, n_2805);
  not g181036 (n_3058, n_2795);
  not g181039 (n_3057, n_2792);
  not g181040 (n_3056, n_2790);
  not g181043 (n_3055, n_2788);
  not g181044 (n_3054, n_2785);
  not g181046 (n_3053, n_2780);
  not g181048 (n_3052, n_2779);
  not g181051 (n_3051, n_2776);
  not g181054 (n_3050, n_2769);
  not g181055 (n_3049, n_2768);
  not g181056 (n_3048, n_2765);
  not g181058 (n_3046, n_2760);
  not g181060 (n_3045, n_2757);
  not g181061 (n_3044, n_2752);
  not g181063 (n_3043, n_2751);
  not g181068 (n_3041, n_2743);
  not g181071 (n_3040, n_2737);
  not g181077 (n_3038, n_2728);
  not g181078 (n_3037, n_2727);
  not g181080 (n_3035, n_2849);
  not g181081 (n_3034, n_2864);
  not g181082 (n_3033, n_2810);
  not g181085 (n_3032, n_3031);
  not g181035 (n_3026, n_2799);
  not g181083 (n_3023, n_2817);
  not g180718 (n_3022, n_3379);
  not g181059 (n_3021, n_2759);
  nand g180520 (n_3020, g3219, n_2474);
  not g181097 (n_3631, n_3510);
  fflopd g218_reg(.CK (clock), .D (g8291), .Q (g218));
  nand g180684 (n_3377, n_2888, n_3019);
  fflopd g550_reg(.CK (clock), .D (n_2451), .Q (g550));
  fflopd g2980_reg(.CK (clock), .D (n_2492), .Q (g2980));
  nand g180690 (n_3372, g35, n_3497);
  fflopd g2984_reg(.CK (clock), .D (n_2679), .Q (g2984));
  nand g180674 (n_3410, g35, n_10391);
  nand g180676 (n_3408, g35, n_10395);
  nand g180683 (n_3732, g35, n_3130);
  fflopd g875_reg(.CK (clock), .D (g14201), .Q (g14217));
  nand g180682 (n_3718, g218, g8291);
  not g180717 (n_3632, n_3018);
  fflopd g4277_reg(.CK (clock), .D (n_2375), .Q (g8839));
  not g180719 (n_4854, n_3017);
  fflopd g376_reg(.CK (clock), .D (n_2698), .Q (g376));
  fflopd g5523_reg(.CK (clock), .D (n_2662), .Q (new_g7738_));
  fflopd g3869_reg(.CK (clock), .D (n_2431), .Q (new_g7121_));
  fflopd g3518_reg(.CK (clock), .D (n_2450), .Q (new_g10323_));
  fflopd g5869_reg(.CK (clock), .D (n_2675), .Q (new_g7766_));
  fflopd g3167_reg(.CK (clock), .D (n_2486), .Q (new_g10295_));
  nor g180689 (n_7331, new_g7753_, new_g7717_);
  fflopd g6215_reg(.CK (clock), .D (n_2663), .Q (new_g7791_));
  not g180036 (n_3016, n_2701);
  nand g180085 (n_3015, g26801, n_2238);
  nand g180087 (n_3014, n_3013, n_2209);
  nand g180088 (n_3012, n_3011, n_2241);
  nand g180089 (n_3010, n_3009, n_2232);
  nand g180090 (n_3008, n_3007, n_2224);
  nand g180091 (n_3006, n_3005, n_2256);
  nor g180093 (n_3004, n_2621, n_3003);
  nor g180094 (n_3002, n_1516, n_3001);
  nor g180095 (n_3000, n_1593, n_2999);
  nand g180096 (n_2998, n_2863, n_2235);
  nor g180105 (n_2997, n_2239, n_2996);
  nand g180123 (n_2995, n_176, n_2284);
  nand g180148 (n_2994, n_2053, n_3364);
  nand g180156 (n_2993, n_224, n_2287);
  nand g180167 (n_2992, n_2624, n_2950);
  nand g180168 (n_2991, n_2634, n_2937);
  nand g180171 (n_2990, n_2632, n_2988);
  nand g180172 (n_2989, n_2971, n_2988);
  nand g180173 (n_2987, n_2617, n_2947);
  nand g180174 (n_2986, n_2627, n_2910);
  nand g180175 (n_2985, n_2712, n_2942);
  nand g180179 (n_2984, n_2629, n_2954);
  nor g180187 (n_2983, new_g8038_, n_2220);
  nand g180194 (n_2982, n_1381, n_2280);
  nor g180195 (n_2981, n_210, n_2980);
  nand g180208 (n_2979, g262, n_2276);
  nand g180804 (n_2978, g12300, n_2169);
  nor g180284 (n_2977, g4527, n_3364);
  nand g180796 (n_2976, n_5346, n_2170);
  nand g180795 (n_2975, g12238, n_2195);
  nand g180792 (n_2974, g11349, n_2309);
  nand g180531 (n_2973, g3259, n_2234);
  nand g180785 (n_2972, n_2631, n_2971);
  nand g180777 (n_2970, n_2800, n_2969);
  nand g180775 (n_2968, n_2753, n_2770);
  nand g180771 (n_2967, g3003, n_9257);
  nand g180765 (n_2966, g7540, n_2050);
  nand g180762 (n_2964, g35, n_2134);
  nand g180757 (n_2963, n_9257, n_2333);
  nand g180755 (n_2962, g35, n_2137);
  nand g180753 (n_2961, n_1129, n_2145);
  nand g180751 (n_2960, n_1525, n_2097);
  nand g180750 (n_2959, n_1387, n_2102);
  nand g180749 (n_2958, n_2957, n_2784);
  nand g180747 (n_2956, n_1690, n_2106);
  nand g180401 (n_2955, n_2677, n_2954);
  nor g180421 (n_2953, n_2291, n_2028);
  nand g180430 (n_2952, g14189, n_5795);
  nand g180435 (n_2951, n_2673, n_2950);
  nand g180436 (n_2949, n_2480, n_2950);
  nand g180447 (n_2948, n_2413, n_2947);
  nand g180457 (n_2946, n_2688, n_2954);
  nand g180458 (n_2945, n_2710, n_2947);
  nand g180461 (n_2944, g5961, n_2213);
  nand g180463 (n_2943, n_2419, n_2942);
  nand g180464 (n_2941, n_2493, n_2942);
  nand g180466 (n_2940, n_2458, n_2942);
  nand g180477 (n_2939, g6307, n_2250);
  nand g180490 (n_2938, n_2705, n_2937);
  nand g180497 (n_2936, g1395, n_2840);
  nand g180499 (n_2935, n_2598, n_2947);
  nand g180501 (n_2934, n_2933, n_2516);
  wire w151, w152, w153, w154;
  nand g180503 (n_2932, w152, w154);
  nand g169 (w154, w153, n_1651);
  not g167 (w153, n_2931);
  nand g166 (w152, w151, n_2931);
  not g165 (w151, n_1651);
  nand g180504 (n_2930, g1495, n_2929);
  nand g180505 (n_2928, g3259, g16603);
  nand g180510 (n_2927, g1489, n_2929);
  nand g180512 (n_2926, n_2482, n_2924);
  nand g180513 (n_2925, n_2473, n_2924);
  nand g180515 (n_2923, n_2476, n_2924);
  nand g180517 (n_2922, n_2465, n_2924);
  wire w155, w156, w157, w158;
  nand g180532 (n_2921, w156, w158);
  nand g173 (w158, w157, n_2920);
  not g172 (w157, n_429);
  nand g171 (w156, w155, n_429);
  not g170 (w155, n_2920);
  wire w159, w160, w161, w162;
  nand g180537 (n_2919, w160, w162);
  nand g178 (w162, w161, n_3512);
  not g177 (w161, n_2042);
  nand g176 (w160, w159, n_2042);
  not g175 (w159, n_3512);
  nand g180540 (n_2918, g3610, g16627);
  nand g180542 (n_2917, n_2693, n_2950);
  wire w163, w164, w165, w166;
  nand g180544 (n_2916, w164, w166);
  nand g183 (w166, w165, n_198);
  not g181 (w165, n_1760);
  nand g180 (w164, w163, n_1760);
  not g179 (w163, n_198);
  nand g180549 (n_2915, n_2681, n_2988);
  nand g180567 (n_2914, g3610, n_2205);
  nand g180575 (n_2913, g3961, g16659);
  nand g180580 (n_2912, n_2490, n_2988);
  nand g180581 (n_2911, n_2670, n_2910);
  nand g180584 (n_2909, n_2666, n_2910);
  nand g180591 (n_2908, g6653, g17688);
  nand g180593 (n_2907, g4669, n_2897);
  nand g180597 (n_2906, g3961, n_2244);
  nand g180599 (n_2905, g5268, n_2246);
  nand g180608 (n_2904, g5268, g17519);
  nand g180615 (n_2903, g5615, n_2226);
  nand g180617 (n_2902, g6653, n_2255);
  nand g180618 (n_2901, n_2445, n_2937);
  nand g180620 (n_2900, g4633, n_2270);
  nand g180621 (n_2899, g35, n_2292);
  nand g180622 (n_2898, g4664, n_2897);
  nand g180624 (n_2896, n_2436, n_2937);
  nand g180625 (n_2895, g854, n_2894);
  nand g180629 (n_2893, g5615, g17580);
  nand g180632 (n_2892, g6307, g17649);
  nand g180636 (n_2891, g5961, g17607);
  nand g180637 (n_2890, n_2699, n_2954);
  nand g180651 (n_2889, g35, n_2888);
  nor g180669 (n_2887, g262, n_2211);
  nand g180686 (n_2886, g4859, n_2288);
  nand g180743 (n_2885, n_1313, n_2254);
  nand g180735 (n_2884, n_1073, n_2152);
  not g180693 (n_2883, n_2676);
  not g180697 (n_2882, n_2665);
  not g180698 (n_2881, n_2664);
  not g180703 (n_2880, n_2370);
  not g180705 (n_2879, n_2538);
  not g180710 (n_2878, n_2877);
  not g180711 (n_2876, n_2875);
  not g180712 (n_2874, g5109);
  not g180713 (n_2873, n_2872);
  nor g180731 (n_2871, g956, n_2781);
  nor g180279 (n_4223, n_1614, n_2307);
  not g180722 (n_3373, new_g7753_);
  not g180720 (n_3375, n_3130);
  nand g180303 (n_3198, n_2870, n_2282);
  fflopd g4284_reg(.CK (clock), .D (n_2221), .Q (new_g8703_));
  nor g180295 (n_3503, n_1599, n_2249);
  nor g180292 (n_3500, n_1601, n_2298);
  nor g180291 (n_3498, n_2614, n_2230);
  nor g180290 (n_3504, n_2609, n_2327);
  fflopd g2946_reg(.CK (clock), .D (n_2216), .Q (g2946));
  fflopd g3976_reg(.CK (clock), .D (g16659), .Q (g16693));
  nand g180340 (n_3538, n_1099, n_2283);
  fflopd g5976_reg(.CK (clock), .D (g17607), .Q (g17646));
  fflopd g6668_reg(.CK (clock), .D (g17688), .Q (g17722));
  fflopd g3274_reg(.CK (clock), .D (g16603), .Q (g16624));
  fflopd g6322_reg(.CK (clock), .D (g17649), .Q (g17685));
  fflopd g5630_reg(.CK (clock), .D (g17580), .Q (g17604));
  nand g180691 (n_3562, g35, n_2980);
  fflopd g5283_reg(.CK (clock), .D (g17519), .Q (g17577));
  fflopd g1589_reg(.CK (clock), .D (n_2218), .Q (new_g6832_));
  fflopd g1246_reg(.CK (clock), .D (n_2231), .Q (new_g6821_));
  fflopd g3625_reg(.CK (clock), .D (g16627), .Q (g16656));
  not g180730 (n_3593, n_3222);
  nand g180692 (n_3570, g35, n_2504);
  nand g180809 (n_2869, g12350, n_2197);
  nand g180812 (n_2868, n_2866, n_2867);
  nand g180816 (n_2865, n_2101, n_1912);
  nand g181360 (n_2864, n_2862, n_2863);
  nand g180840 (n_2861, n_1591, n_2057);
  nand g180851 (n_2860, n_2564, n_2971);
  nand g180857 (n_2859, n_2682, n_2971);
  nand g180860 (n_2858, n_2559, n_2971);
  nand g180874 (n_2857, n_2856, n_2186);
  nand g180877 (n_2855, g817, n_2854);
  nand g180878 (n_2853, n_4343, n_2182);
  nor g180879 (n_2852, g1300, n_2773);
  nand g180883 (n_2851, g1437, n_6350);
  nand g180099 (n_2850, n_2742, n_2258);
  nand g181356 (n_2849, g5212, n_2734);
  nand g180892 (n_2848, g16775, n_2196);
  nand g180901 (n_2847, g1467, n_6352);
  nand g180903 (n_2846, n_1923, n_2126);
  nand g180904 (n_2845, n_2110, n_2140);
  nand g180907 (n_2844, g5037, n_2754);
  fflopd g2932_reg(.CK (clock), .D (n_2215), .Q (g2932));
  nand g180588 (n_2843, n_1582, n_2242);
  nand g181352 (n_2842, n_1903, n_2139);
  nor g180183 (n_2841, g1404, n_2840);
  nand g180453 (n_2839, g35, n_2162);
  nand g180486 (n_2838, n_2690, n_2910);
  nand g181274 (n_2837, n_1905, n_2138);
  not g181042 (n_2836, n_2479);
  not g181030 (n_2834, n_2524);
  not g181038 (n_2833, n_2488);
  not g181041 (n_2832, n_2485);
  not g181052 (n_2830, n_2438);
  not g181064 (n_2829, n_2421);
  not g181074 (n_2828, n_2387);
  nand g180665 (n_2827, n_2826, n_2518);
  not g181088 (n_2825, n_2824);
  not g181093 (n_2822, n_3105);
  not g180706 (n_2821, n_2533);
  not g180714 (n_2820, n_2819);
  not g181094 (n_2818, n_3123);
  nand g181367 (n_2817, n_2816, n_3013);
  nand g181366 (n_2815, n_2813, n_2814);
  nand g181365 (n_2812, n_2811, n_2798);
  nand g181364 (n_2810, n_741, n_2167);
  nand g181359 (n_2809, n_1639, n_2119);
  nand g181122 (n_2808, n_1570, n_2308);
  nand g181123 (n_2807, n_995, n_2092);
  nand g181127 (n_2806, n_2095, n_1965);
  nand g181129 (n_2805, n_544, n_2206);
  nand g181130 (n_2804, n_1072, n_2064);
  nand g181136 (n_2803, n_1275, n_10406);
  nand g181141 (n_2802, n_2098, n_1964);
  nor g181145 (n_2801, n_2800, n_2969);
  nand g181148 (n_2799, g6251, n_2798);
  nand g181336 (n_2797, n_2796, n_2787);
  nand g181152 (n_2795, n_1372, n_2146);
  nand g181160 (n_2794, n_2345, n_2314);
  nand g181163 (n_2793, n_1075, n_2060);
  nand g181169 (n_2792, n_1152, n_2156);
  nand g181171 (n_2791, n_1658, n_2117);
  nand g181172 (n_2790, n_1268, n_2166);
  nand g181177 (n_2789, n_2037, n_2158);
  nand g181181 (n_2788, g3203, n_2787);
  nand g181183 (n_2786, n_1071, n_2176);
  nand g181195 (n_2785, g5559, n_2784);
  nand g181199 (n_2783, n_1644, n_2113);
  nand g181201 (n_2782, g35, n_2781);
  nand g181205 (n_2780, n_1105, n_2150);
  nand g181213 (n_2779, n_794, n_2159);
  nand g181215 (n_2778, n_1578, n_2306);
  nand g181220 (n_2776, g3554, n_2775);
  nand g181223 (n_2774, g35, n_2773);
  nand g181224 (n_2772, n_1068, n_10403);
  nor g181234 (n_2771, g5033, n_2770);
  nand g181242 (n_2769, n_793, n_2072);
  nand g181244 (n_2768, n_536, n_2112);
  nand g181245 (n_2767, n_2766, n_2764);
  nand g181249 (n_2765, g3905, n_2764);
  nand g181256 (n_2763, n_2011, n_2099);
  nand g181257 (n_2762, n_2761, n_2756);
  nand g181258 (n_2760, n_981, n_2153);
  nand g181261 (n_2759, n_2758, n_3011);
  nand g181262 (n_2757, g5905, n_2756);
  nand g181263 (n_2755, n_2753, n_2754);
  nand g181268 (n_2752, g6597, n_2739);
  nand g181270 (n_2751, n_2750, n_3005);
  nand g181275 (n_2749, n_2748, n_2046);
  nand g181278 (n_2747, n_1028, n_2063);
  nand g181294 (n_2746, n_2347, n_2171);
  nand g181297 (n_2745, n_795, n_2071);
  nand g181309 (n_2743, n_2741, n_2742);
  nand g181312 (n_2740, n_2738, n_2739);
  nand g181315 (n_2737, n_2736, g26801);
  nand g181317 (n_2735, n_2733, n_2734);
  nand g181325 (n_2732, n_1904, n_2135);
  nand g181326 (n_2731, n_1140, n_10409);
  nand g181332 (n_2730, g35, n_2770);
  nand g181340 (n_2729, n_1503, n_2115);
  nand g181346 (n_2728, n_723, n_2066);
  nand g181349 (n_2727, n_2726, n_3009);
  nand g181355 (n_2725, n_1585, n_2094);
  fflopd g4153_reg(.CK (clock), .D (n_2245), .Q (g4153));
  nand g181370 (n_3031, n_2455, n_2184);
  nand g181371 (n_3423, n_2723, n_2724);
  nand g181378 (n_3027, n_2039, n_2720);
  nor g181381 (n_3425, n_9257, n_2718);
  nand g181382 (n_3024, n_2202, n_2722);
  nor g180278 (n_3499, n_2612, n_2248);
  nand g180955 (n_3376, n_2721, n_2722);
  nand g180956 (n_3077, n_2719, n_2720);
  nand g181000 (n_3018, n_2717, n_2718);
  not g181095 (n_3472, n_2716);
  nand g181004 (n_3017, g35, n_2854);
  not g181087 (n_3403, n_2501);
  not g181092 (n_3476, n_2715);
  fflopd g996_reg(.CK (clock), .D (n_2228), .Q (g996));
  fflopd g4294_reg(.CK (clock), .D (n_2247), .Q (g10122));
  nand g181396 (n_3510, n_2174, n_2714);
  nand g180973 (n_3374, g4859, n_2969);
  nand g181002 (n_3379, g4340, n_2714);
  fflopd g4467_reg(.CK (clock), .D (n_2143), .Q (g4467));
  fflopd g1339_reg(.CK (clock), .D (n_2229), .Q (g1339));
  fflopd g802_reg(.CK (clock), .D (g12184), .Q (g11678));
  fflopd g4264_reg(.CK (clock), .D (n_2219), .Q (g4264));
  fflopd g896_reg(.CK (clock), .D (n_2233), .Q (g896));
  not g181108 (n_3523, n_3185);
  not g181104 (n_3595, n_3135);
  not g181101 (n_3590, n_3218);
  not g181106 (n_3437, n_3164);
  not g181102 (n_3470, n_3151);
  not g181107 (n_3456, n_3167);
  not g181100 (n_3445, n_3357);
  not g181105 (n_3598, n_3110);
  nand g180850 (n_2713, n_2416, n_2712);
  nand g181143 (n_2711, n_2710, n_2575);
  nand g181140 (n_2709, g35, n_1924);
  not g181468 (n_2708, n_2784);
  nand g180084 (n_2707, n_2127, n_1988);
  nand g181139 (n_2706, n_2705, n_2561);
  not g181423 (n_2704, n_2305);
  nand g181138 (n_2703, n_1016, n_1841);
  nand g180162 (n_2702, n_218, n_2005);
  nand g180262 (n_2701, n_1989, n_1910);
  nand g181135 (n_2700, n_2699, n_2687);
  nand g180496 (n_2698, n_523, n_1993);
  nand g180516 (n_2697, g35, n_1987);
  nand g180602 (n_2696, g35, n_1990);
  nand g180628 (n_2695, g392, n_2006);
  nand g181133 (n_2694, n_2580, n_2693);
  not g180694 (n_2692, n_2302);
  nand g181128 (n_2691, n_2626, n_2690);
  nand g181126 (n_2689, n_2687, n_2688);
  not g180725 (n_2686, g17580);
  nand g181121 (n_2685, new_g10795_, n_1974);
  not g180729 (n_2684, g17607);
  nand g181235 (n_2683, n_2681, n_2682);
  nand g180732 (n_2680, n_2572, n_2688);
  nand g180733 (n_2679, n_1321, n_1847);
  nand g180734 (n_2678, n_2677, n_2687);
  nand g180736 (n_2676, g4854, n_2038);
  nand g180738 (n_2675, n_725, n_1865);
  nand g180739 (n_2674, n_2582, n_2673);
  nand g180740 (n_2672, n_2623, n_2673);
  nand g180741 (n_2671, n_2670, n_2667);
  nand g180744 (n_2669, g4269, n_1785);
  nand g180745 (n_2668, n_2666, n_2667);
  nand g180746 (n_2665, n_737, n_1959);
  nand g180748 (n_2664, g5033, n_2648);
  nand g181120 (n_2663, n_1360, n_1810);
  nand g180752 (n_2662, n_712, n_1800);
  nor g180754 (n_2661, n_1597, n_2027);
  nand g180756 (n_2660, g35, n_1962);
  nand g180758 (n_2659, g35, n_1963);
  nand g180759 (n_2658, g35, n_1826);
  nor g180760 (n_2657, n_1607, n_2023);
  nor g180761 (n_2656, n_1612, n_1979);
  nand g180766 (n_2655, g305, n_9257);
  nand g180767 (n_2654, g2965, n_9257);
  nand g180768 (n_2653, g2927, n_9257);
  nand g180769 (n_2652, g2878, n_9257);
  nand g180770 (n_2651, g2890, n_9257);
  nand g180776 (n_2650, n_2648, n_2649);
  nor g180778 (n_2647, n_485, n_2646);
  nor g180779 (n_2645, n_912, n_2644);
  nor g180780 (n_2643, n_3104, n_2642);
  nand g180781 (n_2641, n_2640, n_2642);
  nand g180782 (n_2639, n_2638, n_2636);
  nor g180783 (n_2637, n_3122, n_2636);
  nand g180784 (n_2635, n_2359, n_2634);
  nand g180786 (n_2633, n_2631, n_2632);
  nand g180787 (n_2630, n_2497, n_2629);
  nand g180788 (n_2628, n_2626, n_2627);
  nand g180789 (n_2625, n_2623, n_2624);
  nor g180791 (n_2622, n_2621, n_1939);
  nor g180794 (n_2620, n_2619, n_2199);
  nand g180797 (n_2618, n_2597, n_2617);
  nand g180798 (n_2616, n_2457, n_2712);
  nor g180799 (n_2615, n_2614, n_1933);
  fflopd g4455_reg(.CK (clock), .D (g4456), .Q (g4455));
  nor g180802 (n_2613, n_2612, n_1947);
  nor g180805 (n_2611, g4966, n_1953);
  nor g180808 (n_2610, n_2609, n_1930);
  nor g180810 (n_2608, g4826, n_2920);
  nand g181361 (n_2607, n_686, n_1951);
  nor g180811 (n_2606, g4776, n_1954);
  nand g180813 (n_2605, n_8824, n_1765);
  nand g180814 (n_2604, n_8825, n_1801);
  nand g180815 (n_2603, n_8823, n_1839);
  nor g180817 (n_2602, g2370, n_2601);
  nand g181363 (n_2599, n_2597, n_2598);
  nand g180821 (n_2595, n_2505, n_10228);
  nor g180822 (n_2594, g1677, n_2593);
  nand g180823 (n_2592, n_8826, n_1796);
  nand g180824 (n_2591, g4669, n_2015);
  nand g180829 (n_2589, n_8829, n_1869);
  nand g180831 (n_2588, n_8822, n_1838);
  nand g180843 (n_2584, n_1777, n_2001);
  nand g180844 (n_2583, n_2624, n_2582);
  nand g180845 (n_2581, n_2580, n_2624);
  nand g180846 (n_2579, n_2627, n_2667);
  nand g180847 (n_2578, n_2634, n_2434);
  nand g180848 (n_2577, n_2712, n_2494);
  nand g180849 (n_2576, n_2617, n_2575);
  nand g181114 (n_2574, n_2710, n_2570);
  nand g180852 (n_2573, n_2629, n_2572);
  nand g180853 (n_2571, n_2617, n_2570);
  nand g180854 (n_2569, n_2712, n_2453);
  nand g180855 (n_2568, g1495, n_2567);
  nand g180856 (n_2566, n_2632, n_2682);
  nand g180858 (n_2565, n_2632, n_2564);
  nand g180859 (n_2563, n_2444, n_2634);
  nand g180861 (n_2562, n_2634, n_2561);
  nand g180862 (n_2560, n_2559, n_2632);
  nand g180863 (n_2558, n_2627, n_2522);
  nand g180864 (n_2557, n_2499, n_2627);
  nand g180865 (n_2556, g4112, n_2553);
  nand g180866 (n_2555, n_2384, n_2629);
  nand g180867 (n_2554, n_1573, n_2553);
  nand g180868 (n_2552, n_2624, n_2403);
  nand g180869 (n_2551, n_2411, n_2617);
  nand g180871 (n_2550, n_2629, n_2687);
  nand g180872 (n_2549, n_2004, n_2567);
  nor g180875 (n_2548, n_1850, n_2547);
  nor g180876 (n_2546, n_2544, n_2545);
  nand g180882 (n_2543, n_1745, n_1603);
  nand g180884 (n_2542, n_1982, n_1602);
  nand g180885 (n_2541, n_1744, n_1600);
  nand g180887 (n_2540, n_2021, n_1669);
  nand g180893 (n_2539, g14662, n_2010);
  nand g180894 (n_2538, n_849, n_2537);
  nand g180895 (n_2536, g14779, n_1743);
  nand g180900 (n_2535, n_2534, n_1872);
  nand g180902 (n_2533, n_1981, n_1919);
  nand g180912 (n_2532, n_1929, n_6454);
  nand g180913 (n_2531, n_1752, n_3773);
  nand g180914 (n_2530, n_1754, n_5760);
  nand g180915 (n_2529, n_1899, n_3767);
  nand g180916 (n_2528, n_1901, n_6450);
  nand g180917 (n_2527, n_1902, n_6456);
  nand g180918 (n_2526, n_1756, n_3769);
  nand g180919 (n_2525, n_1898, n_5758);
  nand g181113 (n_2524, n_1282, n_1973);
  nand g181112 (n_2523, n_2666, n_2522);
  nand g181111 (n_2521, n_2522, n_2690);
  not g181091 (n_2519, n_2518);
  not g181084 (n_2517, n_2516);
  not g181076 (n_2515, n_2240);
  not g181073 (n_2514, n_2322);
  not g181069 (n_2513, n_2316);
  not g181066 (n_2512, n_2279);
  not g181053 (n_2511, n_2300);
  not g181047 (n_2510, n_2212);
  not g181045 (n_2509, n_2214);
  not g181037 (n_2508, n_2222);
  nand g181348 (n_2507, n_174, n_2567);
  fflopd g2873_reg(.CK (clock), .D (n_1799), .Q (g2873));
  nor g180954 (n_2819, n_2506, n_2644);
  fflopd g5452_reg(.CK (clock), .D (n_1782), .Q (g9615));
  fflopd g3100_reg(.CK (clock), .D (g8215), .Q (g3100));
  nor g180953 (n_2872, n_1892, n_2646);
  fflopd g4157_reg(.CK (clock), .D (n_1791), .Q (g4157));
  fflopd g2868_reg(.CK (clock), .D (n_1769), .Q (g2868));
  fflopd g3802_reg(.CK (clock), .D (g8344), .Q (g3802));
  fflopd g4249_reg(.CK (clock), .D (n_1833), .Q (g4249));
  fflopd g2988_reg(.CK (clock), .D (n_1846), .Q (g2988));
  nand g180922 (n_2877, n_2505, n_2017);
  nand g180923 (n_2875, n_914, n_1753);
  fflopd g5109_reg(.CK (clock), .D (g9497), .Q (g5109));
  fflopd g6494_reg(.CK (clock), .D (g9743), .Q (g6494));
  not g181098 (n_3305, n_2980);
  fflopd g6490_reg(.CK (clock), .D (n_1834), .Q (g9817));
  fflopd g3447_reg(.CK (clock), .D (n_1821), .Q (g8342));
  fflopd g6148_reg(.CK (clock), .D (g9682), .Q (g6148));
  nand g180944 (n_3019, g5052, n_1917);
  fflopd g4459_reg(.CK (clock), .D (n_1749), .Q (g4459));
  fflopd g4245_reg(.CK (clock), .D (n_1835), .Q (g4245));
  fflopd g5802_reg(.CK (clock), .D (g9617), .Q (g5802));
  fflopd g3798_reg(.CK (clock), .D (n_1808), .Q (g8398));
  fflopd g5798_reg(.CK (clock), .D (n_2036), .Q (g9680));
  fflopd g5456_reg(.CK (clock), .D (g9555), .Q (g5456));
  fflopd g2491_reg(.CK (clock), .D (n_1828), .Q (g2491));
  fflopd g215_reg(.CK (clock), .D (n_2030), .Q (g8291));
  nand g181028 (n_3222, g35, n_2439);
  fflopd g869_reg(.CK (clock), .D (g14189), .Q (g14201));
  fflopd g2960_reg(.CK (clock), .D (n_1849), .Q (g2960));
  fflopd g2970_reg(.CK (clock), .D (n_1848), .Q (g2970));
  not g180723 (n_3283, g16659);
  not g180727 (n_3290, g16603);
  not g181099 (n_3302, n_2929);
  nor g180994 (n_6177, n_9257, n_2396);
  fflopd g5105_reg(.CK (clock), .D (n_1816), .Q (g9553));
  nand g181005 (n_3130, n_2636, n_6011);
  fflopd g2719_reg(.CK (clock), .D (n_1879), .Q (new_g7753_));
  fflopd g4253_reg(.CK (clock), .D (n_1786), .Q (g4253));
  not g180724 (n_3497, n_2504);
  nand g181014 (n_6019, n_2019, n_2503);
  nor g181027 (n_5660, n_1432, n_2502);
  not g181103 (n_3333, n_2330);
  nand g181373 (n_2501, n_2191, n_2189);
  nand g181149 (n_2500, n_2499, n_2690);
  nand g181150 (n_2498, n_2497, n_2688);
  nand g181155 (n_2496, g376, n_1860);
  nand g181156 (n_2495, n_2493, n_2494);
  nand g181157 (n_2492, n_634, n_1761);
  nand g181159 (n_2491, n_2490, n_2682);
  nand g181162 (n_2489, n_2693, n_2582);
  nand g181166 (n_2488, g1306, n_1983);
  nand g181250 (n_2487, g1760, n_1874);
  nand g181170 (n_2486, n_953, n_1818);
  nand g181175 (n_2485, n_724, n_1730);
  nand g181176 (n_2484, g2485, n_2009);
  nand g181178 (n_2483, n_2475, n_2482);
  nand g181179 (n_2481, n_2480, n_2582);
  nand g181180 (n_2479, n_694, n_1971);
  nand g181182 (n_2478, n_1352, n_1944);
  nand g181184 (n_2477, n_2475, n_2476);
  nand g181185 (n_2474, n_2473, n_2471);
  nand g181186 (n_2472, n_2471, n_2476);
  nand g181187 (n_2470, n_2482, n_2468);
  nand g181188 (n_2469, n_2473, n_2468);
  nand g181189 (n_2467, g1548, n_1830);
  nand g181190 (n_2466, n_2465, n_2468);
  nand g181191 (n_2464, n_2462, n_2482);
  nand g181192 (n_2463, n_2462, n_2473);
  nand g181193 (n_2461, n_2462, n_2476);
  nand g181200 (n_2460, g35, n_1827);
  nand g181202 (n_2459, n_2457, n_2458);
  nand g181207 (n_2456, n_2455, n_1809);
  nand g181209 (n_2454, n_2453, n_2458);
  nand g181211 (n_2452, g3498, n_2335);
  nand g181212 (n_2451, n_987, n_1811);
  nand g181214 (n_2450, n_1179, n_1829);
  nand g181260 (n_2449, g2927, g2922);
  nand g181216 (n_2448, g1657, n_1779);
  nand g181221 (n_2447, n_2677, n_2572);
  nand g181222 (n_2446, n_2444, n_2445);
  nand g181225 (n_2443, n_2490, n_2564);
  nand g181226 (n_2442, n_2681, n_2564);
  nand g181229 (n_2441, n_2465, n_2471);
  nand g181230 (n_2440, g5849, n_2439);
  nand g181232 (n_2438, n_1806, n_1927);
  nand g181236 (n_2437, n_2436, n_2561);
  nand g181238 (n_2435, n_2436, n_2434);
  nand g181239 (n_2433, g3147, n_2336);
  nand g181241 (n_2432, g3849, n_2338);
  nand g181243 (n_2431, n_543, n_1837);
  nand g181246 (n_2430, g2587, n_1787);
  nand g181248 (n_2429, g324, g305);
  nand g181251 (n_2428, n_2670, n_2522);
  nand g181253 (n_2427, n_2667, n_2690);
  nand g181254 (n_2426, n_2499, n_2670);
  nand g181267 (n_2425, n_2434, n_2445);
  nand g181271 (n_2424, n_2423, n_1731);
  nand g181272 (n_2422, g4593, n_1986);
  nand g181273 (n_2421, g962, n_2008);
  nand g181279 (n_2420, n_2419, n_2494);
  nand g181283 (n_2418, g19357, n_1922);
  nand g181284 (n_2417, n_2416, n_2493);
  nand g181285 (n_2415, n_2419, n_2453);
  nand g181286 (n_2414, n_2413, n_2570);
  nand g181288 (n_2412, n_2411, n_2598);
  nand g181289 (n_2410, n_2411, n_2710);
  nand g181290 (n_2409, g336, g305);
  nand g181291 (n_2408, n_2575, n_2598);
  nand g181292 (n_2407, n_2416, n_2458);
  nand g181296 (n_2406, n_2559, n_2490);
  nand g181298 (n_2405, n_2705, n_2434);
  nand g181301 (n_2404, n_2403, n_2673);
  nand g181302 (n_2402, n_936, n_2931);
  nand g181304 (n_2401, g1205, n_1840);
  nand g181307 (n_2400, g5016, n_1766);
  nand g181308 (n_2399, n_2561, n_2445);
  nand g181313 (n_2398, n_2570, n_2598);
  nor g181318 (n_2397, g513, n_2396);
  nand g181319 (n_2395, n_2494, n_2458);
  nand g181321 (n_2394, g2965, g2960);
  nand g181323 (n_2393, n_2444, n_2705);
  nand g181324 (n_2392, n_2468, n_2476);
  nand g181328 (n_2391, n_2413, n_2575);
  nand g181329 (n_2390, n_2580, n_2673);
  nand g181330 (n_2389, n_2480, n_2403);
  nand g181331 (n_2388, n_2693, n_2403);
  nand g181334 (n_2387, g5029, n_1876);
  nand g181335 (n_2386, g4843, n_1737);
  nand g181337 (n_2385, n_2384, n_2699);
  nand g181338 (n_2383, n_2493, n_2453);
  nand g181342 (n_2382, n_775, n_1925);
  nand g181343 (n_2381, g5503, n_2337);
  nand g181347 (n_2380, n_860, n_1878);
  nand g181350 (n_2379, n_2482, n_2471);
  nand g181358 (n_2378, n_2384, n_2688);
  nand g181362 (n_2377, n_2376, n_2007);
  nand g181265 (n_2375, n_1349, n_2013);
  nor g181368 (n_2374, g5821, n_2439);
  nand g181147 (n_2373, g5156, n_2339);
  not g181463 (n_2372, n_2775);
  nand g181276 (n_2371, n_2699, n_2572);
  nand g180870 (n_2370, n_985, n_1949);
  not g181062 (n_2369, n_2164);
  nand g180886 (n_2368, n_2020, n_1666);
  not g181070 (n_2367, n_2319);
  not g180695 (n_2366, n_2301);
  not g181067 (n_2365, n_2120);
  nand g181341 (n_2364, g5097, n_1762);
  not g180709 (n_2363, n_2260);
  not g180726 (n_2362, g17688);
  not g181050 (n_2361, n_2207);
  nand g181282 (n_2360, n_2359, n_2445);
  not g181408 (n_2358, new_g6888_);
  not g181410 (n_2357, n_2141);
  not g181412 (n_2356, n_2130);
  not g181413 (n_2355, n_2129);
  not g181415 (n_2354, n_2123);
  not g181466 (n_2353, n_2764);
  not g181416 (n_2352, n_2121);
  not g181422 (n_2351, n_2289);
  not g181425 (n_2350, n_2084);
  not g181426 (n_2349, n_2083);
  not g181438 (n_2348, n_2347);
  not g181439 (n_2346, n_2345);
  not g181465 (n_2344, n_2787);
  not g181450 (n_2343, n_2756);
  not g181454 (n_2342, n_2734);
  not g181461 (n_2341, n_2739);
  not g181462 (n_2340, n_2798);
  fflopd g2860_reg(.CK (clock), .D (n_1820), .Q (g2860));
  fflopd g3451_reg(.CK (clock), .D (g8279), .Q (g3451));
  fflopd g6144_reg(.CK (clock), .D (n_1836), .Q (g9741));
  fflopd g2894_reg(.CK (clock), .D (n_1863), .Q (g2894));
  fflopd g2852_reg(.CK (clock), .D (n_1802), .Q (g2852));
  fflopd g3096_reg(.CK (clock), .D (n_1844), .Q (g8277));
  nand g181388 (n_2716, g35, n_2183);
  nand g181376 (n_3230, n_2047, n_2193);
  nand g181385 (n_2715, g35, n_2317);
  fflopd g2994_reg(.CK (clock), .D (n_1783), .Q (g2994));
  fflopd g4489_reg(.CK (clock), .D (n_1776), .Q (g4489));
  fflopd g4239_reg(.CK (clock), .D (n_1788), .Q (g4239));
  nand g181384 (n_6494, g35, g305);
  nand g181377 (n_2824, g35, n_2502);
  fflopd g4492_reg(.CK (clock), .D (n_1774), .Q (g4492));
  fflopd g4486_reg(.CK (clock), .D (n_1882), .Q (g4486));
  not g180721 (n_3834, n_2897);
  nand g181404 (n_3110, g35, n_2043);
  nand g181403 (n_3135, g35, n_2339);
  nand g181401 (n_3151, g35, n_2338);
  nand g181400 (n_3218, g35, n_2337);
  fflopd g37_reg(.CK (clock), .D (n_1871), .Q (g37));
  fflopd g2047_reg(.CK (clock), .D (n_1832), .Q (g2047));
  nand g181399 (n_3357, g35, n_2336);
  fflopd g2606_reg(.CK (clock), .D (n_1789), .Q (g2606));
  fflopd g2936_reg(.CK (clock), .D (n_1855), .Q (g2936));
  nand g181387 (n_3123, g1389, n_2636);
  fflopd g2922_reg(.CK (clock), .D (n_1857), .Q (g2922));
  nand g181386 (n_3105, g1046, n_2642);
  fflopd g2223_reg(.CK (clock), .D (n_1771), .Q (g2223));
  fflopd g2950_reg(.CK (clock), .D (n_1852), .Q (g2950));
  fflopd g2472_reg(.CK (clock), .D (n_1819), .Q (g2472));
  fflopd g2204_reg(.CK (clock), .D (n_1767), .Q (g2204));
  fflopd g1779_reg(.CK (clock), .D (n_1812), .Q (g1779));
  fflopd g2625_reg(.CK (clock), .D (n_1866), .Q (g2625));
  not g181446 (n_6441, n_2067);
  fflopd g2912_reg(.CK (clock), .D (n_1858), .Q (g2912));
  fflopd g4146_reg(.CK (clock), .D (n_1794), .Q (g4146));
  fflopd g2357_reg(.CK (clock), .D (n_1843), .Q (g2357));
  fflopd g1913_reg(.CK (clock), .D (n_1807), .Q (g1913));
  fflopd g2066_reg(.CK (clock), .D (n_1748), .Q (g2066));
  nand g181406 (n_3167, g35, n_2044);
  fflopd g1798_reg(.CK (clock), .D (n_1798), .Q (g1798));
  not g180728 (n_3296, g17519);
  nand g181405 (n_3164, g35, n_2335);
  fflopd g2338_reg(.CK (clock), .D (n_2031), .Q (g2338));
  fflopd g1664_reg(.CK (clock), .D (n_1778), .Q (g1664));
  fflopd g1644_reg(.CK (clock), .D (n_1815), .Q (g1644));
  fflopd g2907_reg(.CK (clock), .D (n_1859), .Q (g2907));
  fflopd g1932_reg(.CK (clock), .D (n_1861), .Q (g1932));
  fflopd g94_reg(.CK (clock), .D (n_1856), .Q (g20652));
  fflopd g4639_reg(.CK (clock), .D (n_1740), .Q (new_g10795_));
  fflopd g4843_reg(.CK (clock), .D (n_1995), .Q (g4843));
  fflopd g136_reg(.CK (clock), .D (n_1784), .Q (g21292));
  fflopd g365_reg(.CK (clock), .D (n_2024), .Q (g8719));
  fflopd g1205_reg(.CK (clock), .D (n_1991), .Q (g1205));
  fflopd g1548_reg(.CK (clock), .D (n_1992), .Q (g1548));
  nand g181407 (n_3185, g35, n_2396);
  fflopd g6549_reg(.CK (clock), .D (n_1817), .Q (g6549));
  fflopd g3155_reg(.CK (clock), .D (n_1870), .Q (g3155));
  fflopd g5164_reg(.CK (clock), .D (n_1877), .Q (g5164));
  fflopd g3857_reg(.CK (clock), .D (n_1831), .Q (g3857));
  fflopd g6203_reg(.CK (clock), .D (n_1814), .Q (g6203));
  fflopd g5511_reg(.CK (clock), .D (n_1873), .Q (g5511));
  fflopd g3506_reg(.CK (clock), .D (n_1824), .Q (g3506));
  fflopd g5857_reg(.CK (clock), .D (n_1842), .Q (g5857));
  not g181409 (n_2333, g4108);
  nand g181949 (g28042, n_2331, n_1589);
  nand g181402 (n_2330, g35, n_2198);
  nand g181502 (n_2329, g35, n_5760);
  nand g181320 (n_2328, n_375, n_1502);
  nand g181322 (n_2327, g16744, g13926);
  nor g180772 (n_2326, n_1565, n_2325);
  nand g181333 (n_2324, n_422, n_1686);
  nand g181327 (n_2322, g6283, g17760);
  nand g181316 (n_2321, n_437, n_1687);
  not g181447 (n_2320, g8215);
  nand g181314 (n_2319, g5252, g17674);
  nand g181311 (n_2316, g6291, g17760);
  not g181434 (n_2315, n_2314);
  not g181431 (n_2313, n_2312);
  not g181427 (n_2311, n_2310);
  not g181417 (n_2309, n_1946);
  nand g181679 (n_2308, g6219, n_2091);
  nand g181306 (n_2307, n_254, n_1656);
  nand g181643 (n_2306, g3522, n_2100);
  nand g181636 (n_2305, g6239, n_4988);
  wire w167, w168, w169, w170;
  nand g180677 (n_2304, w168, w170);
  nand g187 (w170, w169, g255);
  not g186 (w169, n_1284);
  nand g185 (w168, w167, n_1284);
  not g184 (w167, g255);
  wire w171, w172, w173, w174;
  nand g180678 (n_2303, w172, w174);
  nand g192 (w174, w173, g246);
  not g190 (w173, n_505);
  nand g189 (w172, w171, n_505);
  not g188 (w171, g246);
  nand g180737 (n_2302, g6629, g17778);
  nand g180742 (n_2301, g5937, g17739);
  nand g181233 (n_2300, g3243, g16718);
  nand g180764 (n_2299, g4477, n_9257);
  nand g181231 (n_2298, g17739, g14738);
  nor g180773 (n_2297, n_1515, n_2296);
  nor g180774 (n_2295, n_1664, n_2294);
  nand g181351 (n_2293, n_315, n_1504);
  nand g180800 (n_2292, g4688, n_143);
  nor g180806 (n_2291, g4688, n_2290);
  nand g181635 (n_2289, g3945, n_5250);
  nor g180820 (n_2288, n_1596, n_2252);
  nor g180827 (n_2287, g8785, n_1621);
  nor g180828 (n_2286, n_1678, n_1626);
  nand g180830 (n_2285, n_58, n_1623);
  nor g180832 (n_2284, g2357, n_1505);
  nor g180833 (n_2283, g4411, n_1631);
  nor g180835 (n_2282, g4087, n_1574);
  nor g180838 (n_2281, n_1647, n_1482);
  nor g180873 (n_2280, g1554, n_1590);
  nand g181303 (n_2279, g5599, g17711);
  nand g180881 (n_2278, g3251, n_2277);
  nor g180888 (n_2276, n_2210, n_1685);
  nand g180897 (n_2275, g5260, n_2274);
  nand g180898 (n_2273, g6645, n_2272);
  nand g180899 (n_2271, n_203, n_1643);
  nand g181300 (n_2270, n_625, n_1528);
  nand g180905 (n_2269, n_117, n_1660);
  nand g180906 (n_2268, n_171, n_1635);
  nand g180908 (n_2267, g5607, n_2266);
  nand g180909 (n_2265, n_188, n_1701);
  nand g180910 (n_2264, g3953, n_2263);
  nand g180911 (n_2262, g5953, n_2261);
  nand g180920 (n_2260, g6299, n_2259);
  nand g181354 (n_2258, n_403, n_1538);
  nand g181299 (n_2257, n_336, n_1688);
  nand g181295 (n_2256, n_287, n_1572);
  nand g181353 (n_2255, n_2413, n_2411);
  nand g181614 (n_2254, g5188, n_2105);
  nand g181293 (n_2253, n_1261, n_2252);
  nand g181287 (n_2251, n_310, n_1449);
  nand g181281 (n_2250, n_2419, n_2416);
  nand g181280 (n_2249, g17711, g14694);
  nand g181277 (n_2248, g17778, g14828);
  nand g181266 (n_2247, n_837, n_1571);
  nand g181264 (n_2246, n_2677, n_2384);
  nand g181259 (n_2245, n_749, n_1533);
  nand g181255 (n_2244, n_2666, n_2499);
  nand g181252 (n_2243, n_299, n_1649);
  nand g181247 (n_2242, n_858, n_1583);
  nand g181240 (n_2241, n_268, n_1670);
  nand g181345 (n_2240, g5945, g17739);
  nand g181237 (n_2239, g6637, g17778);
  nand g181109 (n_2238, n_405, n_1696);
  nand g181110 (n_2237, n_374, n_1640);
  nand g181115 (n_2236, n_307, n_1523);
  nand g181116 (n_2235, n_296, n_1638);
  nand g181117 (n_2234, n_2465, n_2462);
  wire w175, w176, w177, w178;
  nand g181118 (n_2233, w176, w178);
  nand g196 (w178, w177, g862);
  not g195 (w177, n_1984);
  nand g194 (w176, w175, n_1984);
  not g193 (w175, g862);
  nand g181119 (n_2232, n_302, n_1653);
  nand g181124 (n_2231, n_2227, n_1628);
  nand g181131 (n_2230, g17760, g14779);
  nand g181132 (n_2229, n_2217, n_1526);
  nand g181339 (n_2228, n_2227, n_1634);
  nand g181137 (n_2226, n_2480, n_2580);
  nand g181142 (n_2225, n_248, n_1534);
  nand g181146 (n_2224, n_335, n_1587);
  nand g181164 (n_2223, n_270, n_1536);
  nand g181165 (n_2222, g3235, g16718);
  wire w179, w180, w181, w182;
  nand g181167 (n_2221, w180, w182);
  nand g200 (w182, w181, g4281);
  not g199 (w181, n_806);
  nand g198 (w180, w179, n_806);
  not g197 (w179, g4281);
  nand g181168 (n_2220, g499, n_1629);
  wire w183, w184, w185, w186;
  nand g181173 (n_2219, w184, w186);
  nand g205 (w186, w185, g4258);
  not g204 (w185, n_1185);
  nand g202 (w184, w183, n_1185);
  not g201 (w183, g4258);
  nand g181194 (n_2218, n_2217, n_1630);
  wire w187, w188, w189, w190;
  nand g181196 (n_2216, w188, w190);
  nand g210 (w190, w189, g4291);
  not g208 (w189, n_813);
  nand g207 (w188, w187, n_813);
  not g206 (w187, g4291);
  wire w191, w192, w193, w194;
  nand g181197 (n_2215, w192, w194);
  nand g214 (w194, w193, g4308);
  not g213 (w193, n_589);
  nand g212 (w192, w191, n_589);
  not g211 (w191, g4308);
  nand g181203 (n_2214, g3594, g16744);
  nand g181204 (n_2213, n_2436, n_2444);
  nand g181206 (n_2212, n_1522, n_839);
  nand g181208 (n_2211, n_2210, n_1609);
  nand g181210 (n_2209, n_332, n_1532);
  nand g181217 (n_2208, n_1300, n_2014);
  nand g181219 (n_2207, g3586, g16744);
  nand g181664 (n_2206, g5881, n_2118);
  nand g181227 (n_2205, n_2681, n_2559);
  nand g181228 (n_2204, n_351, n_1681);
  nand g181374 (n_2999, g17674, g14662);
  fflopd g4417_reg(.CK (clock), .D (n_1471), .Q (g4417));
  not g181469 (n_2814, n_2203);
  not g181483 (n_2722, n_2644);
  nand g181011 (n_2504, g358, n_1652);
  nand g181383 (n_2518, n_1887, n_1620);
  nand g181380 (n_3003, g16775, g13966);
  nand g181379 (n_2894, n_957, n_1615);
  nand g181375 (n_3001, g16718, g13895);
  nand g181724 (n_2347, g4888, n_2202);
  fflopd g538_reg(.CK (clock), .D (n_1636), .Q (g538));
  nand g180933 (n_2888, n_5549, n_1604);
  not g181475 (n_2720, n_2646);
  fflopd g4141_reg(.CK (clock), .D (n_1467), .Q (g4141));
  not g181449 (n_2718, n_2201);
  not g181460 (n_2813, n_2200);
  fflopd g4172_reg(.CK (clock), .D (n_1693), .Q (g4172));
  not g181459 (n_2867, n_2199);
  nand g181369 (n_2516, n_1719, n_1619);
  nand g181389 (n_2840, g12923, n_1513);
  nand g181007 (n_2897, g4688, n_1003);
  nand g181745 (n_2734, new_g7704_, n_1689);
  fflopd g4087_reg(.CK (clock), .D (n_1477), .Q (g4087));
  not g181445 (n_6350, n_1895);
  nand g180992 (n_3364, g4489, n_1627);
  nand g180993 (n_2947, g35, n_1885);
  nand g180999 (n_2950, g35, n_1725);
  fflopd g3969_reg(.CK (clock), .D (g16775), .Q (g16659));
  nand g181390 (n_2910, g35, n_1717);
  nand g181391 (n_2954, g35, n_1884);
  fflopd g4057_reg(.CK (clock), .D (n_1468), .Q (g4057));
  nand g181392 (n_2988, g35, n_1883);
  nand g181393 (n_2924, g35, n_1718);
  nand g181395 (n_2937, g35, n_1888);
  nand g181398 (n_2929, g35, n_1712);
  fflopd g3267_reg(.CK (clock), .D (g16718), .Q (g16603));
  fflopd g5276_reg(.CK (clock), .D (g17674), .Q (g17519));
  fflopd g3618_reg(.CK (clock), .D (g16744), .Q (g16627));
  fflopd g6315_reg(.CK (clock), .D (g17760), .Q (g17649));
  fflopd g6661_reg(.CK (clock), .D (g17778), .Q (g17688));
  fflopd g5623_reg(.CK (clock), .D (g17711), .Q (g17580));
  nor g181029 (n_5795, n_9257, n_2198);
  not g181418 (n_2197, n_1942);
  not g181420 (n_2196, n_1940);
  not g181424 (n_2195, n_1913);
  not g181432 (n_2188, n_2187);
  not g181436 (n_2186, n_2185);
  not g181442 (n_2184, n_2183);
  not g181440 (n_2182, n_2181);
  not g181448 (n_2180, g9617);
  not g181451 (n_2179, g8279);
  not g181452 (n_2178, g9555);
  not g181798 (n_2177, n_1862);
  nand g181494 (n_2176, g35, n_1496);
  not g181457 (n_2175, g9743);
  not g181458 (n_2174, n_2619);
  not g181464 (n_2173, g8344);
  not g181433 (n_2172, n_2171);
  not g181473 (n_2170, n_2396);
  not g181419 (n_2169, n_1941);
  not g181453 (n_2168, g9682);
  nand g181682 (n_2167, g6573, n_2093);
  nand g181641 (n_2166, g3179, n_2116);
  nand g181563 (n_2165, g2429, n_2133);
  nand g181269 (n_2164, g5244, g17674);
  not g181486 (n_2163, g305);
  nand g180880 (n_2162, n_2866, n_1478);
  nand g181496 (n_2160, g35, n_6456);
  nand g181497 (n_2159, g35, n_5157);
  fflopd g3003_reg(.CK (clock), .D (n_1672), .Q (g3003));
  nand g181501 (n_2158, g35, n_2157);
  nand g181504 (n_2156, g35, n_5145);
  nand g181507 (n_2155, g35, n_6454);
  fflopd g4164_reg(.CK (clock), .D (n_1677), .Q (new_g6888_));
  nand g181510 (n_2154, g35, n_3767);
  nand g181512 (n_2153, g35, n_5089);
  nand g181513 (n_2152, g35, n_1668);
  nand g181516 (n_2151, g35, n_3773);
  nand g181519 (n_2150, g35, n_5039);
  nand g181521 (n_2148, g35, n_6450);
  nand g181523 (n_2147, g35, n_1495);
  nand g181524 (n_2146, g35, n_5047);
  nand g181526 (n_2145, g35, n_5199);
  nand g181530 (n_2144, new_g6961_, n_2142);
  nand g181532 (n_2143, n_246, n_2142);
  nand g181535 (n_2141, g4462, n_2070);
  nand g181544 (n_2140, g1600, n_1476);
  nand g181547 (n_2139, g2295, n_1703);
  nand g181550 (n_2138, g1870, n_2136);
  nor g181553 (n_2137, g1945, n_2136);
  nand g181560 (n_2135, g2161, n_1691);
  nor g181564 (n_2134, g2504, n_2133);
  nand g181565 (n_2132, n_1972, n_2131);
  nand g181567 (n_2130, g3227, n_6884);
  nand g181568 (n_2129, g3929, n_5789);
  nand g181576 (n_2128, n_2127, n_1894);
  nand g181578 (n_2126, g1620, g25167);
  nor g181579 (n_2125, n_1426, n_2124);
  nand g181581 (n_2123, g3578, n_4646);
  nand g181310 (n_2122, n_318, n_1637);
  nand g181583 (n_2121, g3602, n_4646);
  nand g181305 (n_2120, g5591, g17711);
  nand g181617 (n_2119, g5873, n_2118);
  nand g181625 (n_2117, g3171, n_2116);
  nand g181626 (n_2115, g5092, n_1463);
  nand g181630 (n_2114, g2093, n_8568);
  nand g181639 (n_2113, g3873, n_2111);
  nand g181640 (n_2112, g3881, n_2111);
  nand g181644 (n_2110, n_2109, n_1673);
  nand g181647 (n_2108, n_2107, n_4988);
  nand g181648 (n_2106, g5180, n_2105);
  nand g181651 (n_2104, n_2103, n_5250);
  nand g181654 (n_2102, g5535, n_2096);
  nand g181656 (n_2101, g3530, n_2100);
  nand g181582 (n_2099, g2004, n_8568);
  nand g181663 (n_2098, g1792, n_1492);
  nand g181669 (n_2097, g5527, n_2096);
  nand g181680 (n_2095, g2619, n_1704);
  nand g181681 (n_2094, g6565, n_2093);
  nand g181683 (n_2092, g6227, n_2091);
  nand g181684 (n_2090, n_1139, n_4952);
  nand g181685 (n_2089, n_2088, n_4952);
  nand g181686 (n_2087, n_2086, n_5126);
  nand g181688 (n_2085, n_811, n_5128);
  nand g181691 (n_2084, g3191, n_4168);
  nand g181692 (n_2083, g5200, n_4922);
  nand g181693 (n_2082, n_2081, n_4922);
  nand g181694 (n_2080, n_2079, n_4168);
  nand g181695 (n_2078, n_807, n_5126);
  nand g181696 (n_2077, n_884, n_5130);
  nand g181697 (n_2076, n_2075, n_5130);
  nand g181698 (n_2074, n_2073, n_5128);
  nand g181955 (n_2072, g35, n_5186);
  nand g181906 (n_2071, n_226, n_2070);
  nand g181872 (n_2069, g35, n_5758);
  nand g181871 (n_2068, g35, n_3769);
  nand g181735 (n_2067, g13272, n_2157);
  nand g181870 (n_2066, g35, n_5098);
  nand g181867 (n_2064, g35, n_1667);
  nand g181861 (n_2063, g35, n_1494);
  nand g181860 (n_2062, g35, n_1485);
  nand g181859 (n_2061, g35, n_1674);
  nand g181858 (n_2060, g35, n_1514);
  not g181797 (n_2059, n_1864);
  not g181799 (n_2058, n_1854);
  not g181803 (n_2057, n_1813);
  not g181806 (n_2055, n_1790);
  not g181809 (n_2054, n_1781);
  not g181810 (n_2053, n_1772);
  not g181811 (n_2052, n_1768);
  not g181813 (n_2051, n_1739);
  not g181816 (n_2050, n_2049);
  nand g181856 (n_2046, g35, n_1497);
  not g181455 (n_2742, n_2044);
  not g181823 (n_2724, n_1755);
  not g181456 (n_2863, n_2043);
  not g181470 (n_2714, n_2042);
  not g181471 (n_2754, n_2648);
  not g181478 (n_3007, n_2439);
  not g181834 (n_7413, n_2041);
  nand g181699 (n_2773, g1484, n_1474);
  nand g181712 (n_2748, g4375, n_2040);
  nand g181725 (n_2345, g4698, n_2039);
  nand g181719 (n_2781, g1141, n_1473);
  nand g181754 (n_2798, new_g7791_, n_1650);
  nand g181760 (n_2784, new_g7738_, n_1483);
  nand g181741 (n_2756, new_g7766_, n_1508);
  not g181482 (n_3005, n_2337);
  not g181480 (n_3009, n_2336);
  not g181444 (n_6352, n_2025);
  nand g181753 (n_2739, new_g7812_, n_1484);
  not g181477 (n_3013, n_2335);
  not g181833 (n_2854, n_1750);
  fflopd g799_reg(.CK (clock), .D (n_1470), .Q (g12184));
  nand g181755 (n_2775, new_g10323_, n_1682);
  not g181474 (n_2770, n_2649);
  not g181479 (n_3011, n_2338);
  nand g181757 (n_2787, new_g10295_, n_1683);
  nand g181758 (n_2764, new_g7121_, n_1679);
  fflopd g4304_reg(.CK (clock), .D (n_1568), .Q (g9251));
  nand g181394 (n_2942, g35, n_1714);
  not g181476 (n_2969, n_2038);
  nand g181397 (n_2980, g358, n_1611);
  not g181490 (g26801, n_2339);
  not g181835 (n_2971, n_1729);
  fflopd g5969_reg(.CK (clock), .D (g17739), .Q (g17607));
  nand g181621 (n_2037, g1526, n_1980);
  nand g181882 (n_2036, n_372, n_1333);
  nand g181973 (n_2035, g1404, n_821);
  nand g181877 (n_2034, g35, n_1519);
  fflopd g2878_reg(.CK (clock), .D (n_610), .Q (g2878));
  nand g181876 (n_2033, g4375, n_2032);
  nand g181976 (n_2031, n_350, n_683);
  nand g181873 (n_2030, n_974, n_614);
  fflopd g4456_reg(.CK (clock), .D (n_1251), .Q (g4456));
  nand g181868 (n_2029, g35, n_1093);
  nor g181866 (n_2028, n_9257, n_1092);
  nor g181865 (n_2027, n_9257, n_1101);
  nand g181864 (n_2026, g35, n_1210);
  nand g181732 (n_2025, g13272, n_2856);
  nor g181506 (n_2024, n_9257, n_525);
  nor g181863 (n_2023, n_9257, n_501);
  nand g181857 (n_2022, g35, n_1926);
  not g181488 (n_2021, g16744);
  not g181485 (n_2020, g17778);
  not g181472 (n_2019, g990);
  nand g181855 (n_2018, g35, n_1395);
  not g181818 (n_2017, n_2016);
  not g181437 (n_2015, n_2014);
  nand g181854 (n_2013, g35, n_1374);
  nand g181687 (n_2011, g2060, n_1064);
  not g181411 (n_2010, n_1622);
  nand g181853 (n_2009, n_308, n_976);
  nand g181670 (n_2008, g7916, n_4343);
  nand g181593 (n_2007, n_1059, n_1174);
  nand g180841 (n_2006, n_113, n_1172);
  nor g180842 (n_2005, n_1157, n_1164);
  not g181832 (n_2004, n_5035);
  not g181819 (n_2001, n_2000);
  nand g181615 (n_1997, g3698, n_3627);
  wire w195, w196, w197, w198;
  nand g181125 (n_1996, w196, w198);
  nand g219 (w198, w197, g979);
  not g217 (w197, g1236);
  nand g216 (w196, w195, g1236);
  not g215 (w195, g979);
  wire w199, w200, w201, w202;
  nand g181144 (n_1995, w200, w202);
  nand g224 (w202, w201, n_1994);
  not g223 (w201, n_279);
  nand g221 (w200, w199, n_279);
  not g220 (w199, n_1994);
  nand g181151 (n_1993, g35, n_1162);
  wire w203, w204, w205, w206;
  nand g181153 (n_1992, w204, w206);
  nand g229 (w206, w205, n_5);
  not g228 (w205, n_402);
  nand g227 (w204, w203, n_402);
  not g226 (w203, n_5);
  wire w207, w208, w209, w210;
  nand g181154 (n_1991, w208, w210);
  nand g234 (w210, w209, n_56);
  not g233 (w209, n_247);
  nand g231 (w208, w207, n_247);
  not g230 (w207, n_56);
  wire w211, w212, w213, w214;
  nand g181158 (n_1990, w212, w214);
  nand g238 (w214, w213, g4273);
  not g237 (w213, n_1625);
  nand g236 (w212, w211, n_1625);
  not g235 (w211, g4273);
  nand g181161 (n_1989, g437, n_1161);
  wire w215, w216, w217, w218;
  nand g181198 (n_1988, w216, w218);
  nand g243 (w218, w217, n_624);
  not g242 (w217, n_1527);
  nand g241 (w216, w215, n_1527);
  not g240 (w215, n_624);
  wire w219, w220, w221, w222;
  nand g181174 (n_1987, w220, w222);
  nand g248 (w222, w221, g20557);
  not g247 (w221, n_1481);
  nand g245 (w220, w219, n_1481);
  not g244 (w219, g20557);
  nor g181598 (n_1986, g4601, n_963);
  nand g181596 (n_1985, g896, n_1984);
  nand g181592 (n_1983, g7946, n_2856);
  not g181484 (n_1982, g17739);
  nand g181492 (n_1981, g1514, n_1980);
  nor g181498 (n_1979, n_9257, n_1065);
  nand g181499 (n_1978, g35, n_956);
  nand g181503 (n_1977, g35, n_1218);
  nand g181511 (n_1976, g35, n_1886);
  fflopd g2890_reg(.CK (clock), .D (n_1344), .Q (g2890));
  nand g181517 (n_1975, g35, n_1056);
  fflopd g4108_reg(.CK (clock), .D (n_628), .Q (g4108));
  nand g181522 (n_1974, g35, n_1212);
  nand g181531 (n_1973, g1178, n_1972);
  nand g181540 (n_1971, g1521, n_1918);
  nand g181562 (n_1967, n_1966, n_865);
  nand g181566 (n_1965, g2563, n_8577);
  nand g181569 (n_1964, g1736, n_8579);
  nor g181570 (n_1963, g1811, n_8579);
  nor g181571 (n_1962, g2638, n_8577);
  nand g181573 (n_1961, g1532, n_1980);
  nand g181574 (n_1960, g1189, n_1958);
  nand g181575 (n_1959, g1178, n_1958);
  nand g181585 (n_1957, n_81, n_1424);
  nand g181587 (n_1956, n_1955, n_834);
  nand g181589 (n_1954, n_1558, n_1436);
  nand g181590 (n_1953, n_1559, n_1435);
  nand g181591 (n_1952, g4040, n_809);
  nand g181594 (n_1951, g7946, n_1950);
  nand g181597 (n_1949, n_167, n_1948);
  nand g181599 (n_1947, g6601, n_3272);
  nand g181600 (n_1946, g3207, n_1945);
  nand g181601 (n_1944, g168, n_1376);
  nand g181602 (n_1943, g4049, n_5154);
  nand g181603 (n_1942, g5909, n_5148);
  nand g181604 (n_1941, g5563, n_5152);
  nand g181605 (n_1940, g3937, n_5154);
  nand g181606 (n_1939, g3909, n_5154);
  nand g181607 (n_1938, g5698, n_5152);
  nand g181608 (n_1937, g6044, n_5148);
  nand g181609 (n_1936, g6390, n_5150);
  nand g181611 (n_1933, g6255, n_5150);
  nand g181612 (n_1932, g6736, n_3272);
  nand g181613 (n_1931, g3347, n_1945);
  nand g181616 (n_1930, g3558, n_3627);
  not g181815 (n_1929, n_1486);
  nand g181623 (n_1928, g17400, n_1732);
  nand g181627 (n_1927, g4311, n_1926);
  nand g181628 (n_1925, g1183, n_1958);
  nor g181633 (n_1924, g5022, n_1875);
  nand g181637 (n_1923, n_1009, n_1090);
  nand g181638 (n_1922, n_222, n_992);
  nand g181642 (n_1921, g4358, n_1920);
  nand g181645 (n_1919, n_472, n_1918);
  nor g181646 (n_1917, n_1916, n_602);
  nand g181650 (n_1915, g1171, n_1958);
  nand g181653 (n_1914, g5352, g25114);
  nand g181660 (n_1913, g5216, g25114);
  nand g181662 (n_1912, n_968, n_1890);
  nand g181666 (n_1911, g392, n_935);
  nand g181667 (n_1910, n_1909, n_1060);
  nand g181668 (n_1908, n_975, n_808);
  nand g181671 (n_1907, g691, n_850);
  nand g181672 (n_1906, n_524, n_1889);
  nand g181676 (n_1905, g1926, n_810);
  nand g181689 (n_1904, g2217, n_812);
  nand g181690 (n_1903, g2351, n_1236);
  not g181814 (n_1902, n_1586);
  not g181807 (n_1901, n_1697);
  not g181801 (n_1899, n_1654);
  not g181795 (n_1898, n_1576);
  not g181794 (n_1897, n_1575);
  nand g181734 (n_1895, g13272, n_1950);
  fflopd g4098_reg(.CK (clock), .D (n_627), .Q (g4098));
  nand g181717 (n_2314, g4743, n_2719);
  nor g181722 (n_2547, n_1433, n_1103);
  nand g181728 (n_2181, g996, n_1972);
  nand g181730 (n_2183, g1087, n_1167);
  nand g181731 (n_2317, g1430, n_1156);
  nand g181713 (n_2187, g4785, n_971);
  nand g181751 (n_2199, g4633, n_1894);
  nand g181752 (n_2200, g35, n_10238);
  nand g181762 (n_2203, g35, n_10240);
  nand g181763 (n_2042, g4628, n_1894);
  nand g181714 (n_4153, n_820, n_300);
  nor g181726 (n_2545, n_1434, n_1288);
  nand g181774 (n_2038, g4878, n_1219);
  nand g181747 (n_2043, new_g7812_, n_1345);
  nand g181746 (n_2044, new_g7791_, n_1208);
  nand g181711 (n_2312, n_120, n_1893);
  nor g181710 (n_3491, n_128, n_1892);
  nor g181709 (n_3493, n_22, n_2506);
  fflopd g2965_reg(.CK (clock), .D (n_632), .Q (g2965));
  fflopd g2927_reg(.CK (clock), .D (n_1397), .Q (g2927));
  nand g181704 (n_2191, g35, n_10244);
  nand g181702 (n_2193, g35, n_10242);
  nand g181700 (n_2310, g4975, n_1211);
  fflopd g4082_reg(.CK (clock), .D (n_622), .Q (g4082));
  nand g181705 (n_2189, g35, n_10250);
  not g181441 (n_2537, n_1676);
  nand g181716 (n_2171, g4933, n_2721);
  nand g181749 (n_2619, g4340, n_509);
  nand g181772 (n_2649, n_1891, n_1041);
  nand g181777 (n_2338, new_g7121_, n_800);
  fflopd g6140_reg(.CK (clock), .D (n_856), .Q (g9682));
  nand g181775 (n_2335, new_g10323_, n_875);
  fflopd g3794_reg(.CK (clock), .D (n_1159), .Q (g8344));
  nand g181778 (n_2336, new_g10295_, n_1186);
  fflopd g3443_reg(.CK (clock), .D (n_1890), .Q (g8279));
  fflopd g5448_reg(.CK (clock), .D (n_746), .Q (g9555));
  fflopd g3092_reg(.CK (clock), .D (n_817), .Q (g8215));
  nand g181781 (n_2337, new_g7738_, n_1320);
  fflopd g5794_reg(.CK (clock), .D (n_1310), .Q (g9617));
  fflopd g6486_reg(.CK (clock), .D (n_1379), .Q (g9743));
  not g181491 (n_2920, g4688);
  nand g181740 (n_2502, g1193, n_1429);
  nand g181764 (n_2648, g5062, n_492);
  nand g181768 (n_2931, g8719, n_1889);
  not g181846 (n_5094, n_1888);
  not g181847 (n_2642, n_1887);
  nand g181770 (n_2396, g358, n_1886);
  nand g181773 (n_2646, g4776, n_990);
  nand g181776 (n_2439, new_g7766_, n_1357);
  fflopd g5101_reg(.CK (clock), .D (n_881), .Q (g9497));
  not g181842 (n_5056, n_1885);
  nand g181782 (n_2644, g4966, n_999);
  not g181839 (n_5201, n_1884);
  not g181837 (n_5190, n_1883);
  nand g182144 (n_2458, g35, n_2811);
  nand g182154 (n_2598, g35, n_2738);
  not g181851 (n_2624, n_1501);
  not g181838 (n_2627, n_1510);
  not g181841 (n_2629, n_1507);
  not g181843 (n_2634, n_1531);
  not g181845 (n_2712, n_1702);
  nand g182147 (n_2445, g35, n_2761);
  nand g182131 (n_2688, g35, n_2733);
  fflopd g305_reg(.CK (clock), .D (n_558), .Q (g305));
  nand g182030 (n_1882, n_1881, n_986);
  nand g181885 (n_1880, g1193, n_2544);
  nand g181892 (n_1879, n_9257, n_3197);
  nand g181893 (n_1878, n_1549, n_5216);
  nor g181894 (n_1877, g5164, n_2497);
  nand g181895 (n_1876, n_612, n_1875);
  nand g181896 (n_1874, n_283, n_677);
  nor g181899 (n_1873, g5511, n_2623);
  nand g181901 (n_1872, n_442, n_864);
  nand g181902 (n_1871, n_380, n_1341);
  nor g181904 (n_1870, g3155, n_2475);
  nand g181907 (n_1869, n_249, n_1052);
  nand g181908 (n_1868, g35, n_1867);
  nand g181909 (n_1866, n_272, n_824);
  nand g181911 (n_1865, n_1438, n_5197);
  nand g181912 (n_1864, n_311, n_1123);
  nand g181913 (n_1863, n_385, n_696);
  nand g181914 (n_1862, n_295, n_1062);
  nand g181915 (n_1861, n_338, n_690);
  nand g181916 (n_1860, g35, n_958);
  nand g181917 (n_1859, n_298, n_716);
  nand g181918 (n_1858, n_251, n_1224);
  nand g181919 (n_1857, n_371, n_1177);
  nand g181920 (n_1856, n_288, n_1021);
  nand g181921 (n_1855, n_341, n_756);
  nand g181922 (n_1854, n_294, n_1853);
  nand g181923 (n_1852, n_342, n_638);
  nand g181924 (n_1851, g1536, n_1850);
  nand g181925 (n_1849, n_393, n_973);
  nand g181926 (n_1848, n_281, n_1146);
  nand g181927 (n_1847, g35, n_552);
  nand g181928 (n_1846, n_1845, n_830);
  nand g181929 (n_1844, n_1297, n_1035);
  nand g181930 (n_1843, n_280, n_1315);
  nor g181931 (n_1842, g5857, n_2359);
  nand g181932 (n_1841, n_1440, n_5195);
  nand g181933 (n_1840, g35, n_862);
  nand g181934 (n_1839, n_289, n_1018);
  nand g181936 (n_1838, n_321, n_885);
  nand g181937 (n_1837, n_1441, n_5193);
  nand g181938 (n_1836, n_344, n_671);
  nand g181939 (n_1835, n_258, n_1304);
  nand g181941 (n_1834, n_278, n_555);
  nand g181942 (n_1833, n_347, n_533);
  nand g181946 (n_1832, n_409, n_507);
  nor g181948 (n_1831, g3857, n_2626);
  nand g181950 (n_1830, g35, n_1382);
  nand g181951 (n_1829, n_1556, n_5160);
  nand g181952 (n_1828, n_439, n_871);
  nand g181953 (n_1827, n_260, n_1020);
  nor g181954 (n_1826, n_1825, n_6011);
  nor g181956 (n_1824, g3506, n_2631);
  nand g181957 (n_1823, g518, n_5346);
  nand g181958 (n_1822, n_438, n_1143);
  nand g181959 (n_1821, n_426, n_814);
  nand g181960 (n_1820, n_417, n_650);
  nand g181961 (n_1819, n_252, n_1066);
  nand g181963 (n_1818, n_1551, n_5170);
  nor g181964 (n_1817, g6549, n_2597);
  nand g181965 (n_1816, n_804, n_616);
  nand g181967 (n_1815, n_432, n_1215);
  nor g181969 (n_1814, g6203, n_2457);
  nand g181970 (n_1813, n_441, n_604);
  nand g181971 (n_1812, n_420, n_652);
  nand g181972 (n_1811, g35, n_1074);
  nand g181974 (n_1810, n_1442, n_5044);
  nor g181975 (n_1809, g1205, n_1351);
  nand g181980 (n_1808, n_1367, n_1136);
  nand g181982 (n_1807, n_399, n_1057);
  nand g181983 (n_1806, n_1805, n_993);
  nand g181984 (n_1804, g35, n_1803);
  nand g181985 (n_1802, n_391, n_1122);
  nand g181987 (n_1801, n_301, n_1014);
  nand g181988 (n_1800, n_1550, n_5220);
  nand g181990 (n_1799, n_340, n_762);
  nand g181991 (n_1798, n_325, n_570);
  nand g181992 (n_1797, n_354, n_926);
  nand g181993 (n_1796, n_312, n_1053);
  nand g181995 (n_1795, g35, n_1487);
  nand g181996 (n_1794, n_282, n_750);
  nand g181999 (n_1793, g35, n_1489);
  nand g182001 (n_1792, n_428, n_666);
  nand g182004 (n_1791, n_443, n_734);
  nand g182006 (n_1790, n_414, n_1237);
  nand g182008 (n_1789, n_349, n_1358);
  nand g182009 (n_1788, n_1170, n_629);
  nand g182011 (n_1787, n_255, n_980);
  nand g182014 (n_1786, n_253, n_676);
  nand g182015 (n_1785, n_623, n_1067);
  nand g182016 (n_1784, n_430, n_500);
  nand g182022 (n_1783, n_377, n_929);
  nand g182023 (n_1782, n_390, n_1346);
  nand g182024 (n_1781, n_392, n_1780);
  nand g182026 (n_1779, n_411, n_1010);
  nand g182028 (n_1778, n_245, n_1327);
  nand g181883 (n_1777, n_802, n_2423);
  nand g182031 (n_1776, n_1775, n_513);
  nand g182032 (n_1774, n_1773, n_836);
  nand g182036 (n_1772, n_1845, n_585);
  nand g182037 (n_1771, n_309, n_1302);
  wire w223, w224, w225, w226;
  nand g181134 (n_1770, w224, w226);
  nand g252 (w226, w225, g1579);
  not g251 (w225, n_3496);
  nand g250 (w224, w223, n_3496);
  not g249 (w223, g1579);
  nand g182038 (n_1769, n_396, n_1373);
  nand g182039 (n_1768, n_337, n_1287);
  nand g182042 (n_1767, n_267, n_736);
  nand g182045 (n_1766, g35, n_596);
  nand g182047 (n_1765, n_381, n_1017);
  nand g182048 (n_1764, g35, n_1763);
  nand g182055 (n_1762, n_611, n_1027);
  nand g181525 (n_1761, g35, n_539);
  nand g182060 (n_1760, g2250, n_8551);
  nand g182061 (n_1759, g1950, n_1318);
  nand g182067 (n_1758, g1816, n_1452);
  nand g182068 (n_1757, g1682, n_583);
  not g181796 (n_1756, n_1579);
  nand g182075 (n_1755, n_511, n_1920);
  not g181802 (n_1754, n_1663);
  not g181808 (n_1753, n_1700);
  not g181800 (n_1752, n_1648);
  not g181812 (n_1751, n_1537);
  nand g182088 (n_1750, n_1581, n_996);
  nand g182027 (n_1749, n_1555, n_1437);
  nand g182025 (n_1748, n_376, n_841);
  not g181435 (n_1747, n_1746);
  not g181487 (n_1745, g17760);
  not g181489 (n_1744, g17711);
  not g181414 (n_1743, n_1580);
  nor g181577 (n_1740, new_g10795_, n_1439);
  nand g182041 (n_1739, n_333, n_1738);
  nand g182049 (n_1737, g35, n_1401);
  nand g182059 (n_1736, g2241, n_1460);
  nand g182077 (n_1735, g2509, n_1605);
  nand g181559 (n_1733, g1052, n_1732);
  nand g181665 (n_1731, g4584, n_803);
  nand g181572 (n_1730, g1521, n_1980);
  nand g182130 (n_1729, n_1577, n_1165);
  nand g182078 (n_2593, g1691, n_8550);
  nand g182089 (n_2041, g35, n_1728);
  nand g181739 (n_2201, g1536, n_1431);
  nand g182072 (n_2047, g35, n_10232);
  nand g181720 (n_2185, g1339, n_1918);
  nand g182062 (n_2049, g35, n_840);
  nand g182076 (n_2601, g2384, n_8548);
  nor g182058 (n_2723, new_g12440_, n_876);
  fflopd g4093_reg(.CK (clock), .D (n_621), .Q (g4093));
  nor g181727 (n_2553, n_1095, n_954);
  nand g181759 (n_3387, g35, n_10252);
  fflopd g859_reg(.CK (clock), .D (n_1182), .Q (g14189));
  fflopd g4076_reg(.CK (clock), .D (n_590), .Q (g4076));
  nand g182079 (n_4193, g35, n_10254);
  nand g181792 (n_2339, new_g7704_, n_801);
  nand g182118 (n_2453, g35, n_1727);
  nand g182099 (n_2575, g35, n_1726);
  not g181850 (n_5105, n_1725);
  nand g182116 (n_2473, g35, n_1724);
  nand g182113 (n_2561, g35, n_1723);
  nand g182129 (n_2705, g35, n_1722);
  nand g182111 (n_2693, g35, n_1721);
  nand g182108 (n_2494, g35, n_1414);
  nand g182126 (n_2699, g35, n_1720);
  nand g182127 (n_2570, g35, n_1416);
  not g181848 (n_2636, n_1719);
  not g181844 (n_5073, n_1718);
  not g181840 (n_5178, n_1717);
  nand g182107 (n_2522, g35, n_1716);
  nand g182117 (n_2687, g35, n_1546);
  nand g182105 (n_2710, g35, n_1715);
  not g181836 (n_5085, n_1714);
  nand g182104 (n_2572, g35, n_1713);
  not g181481 (n_2567, n_1712);
  nand g182098 (n_2682, g35, n_1711);
  nand g182097 (n_2493, g35, n_1710);
  nand g182101 (n_2667, g35, n_1415);
  nand g182128 (n_2468, g35, n_1412);
  fflopd g4258_reg(.CK (clock), .D (n_597), .Q (g4258));
  nand g182095 (n_2403, g35, n_1542);
  nand g182092 (n_2564, g35, n_1544);
  nand g182090 (n_2582, g35, n_1709);
  nand g182122 (n_2434, g35, n_1541);
  nand g182121 (n_2471, g35, n_1708);
  nand g182124 (n_2670, g35, n_1707);
  nand g182102 (n_2490, g35, n_1706);
  not g181849 (n_2617, n_1659);
  not g181852 (n_2632, n_1499);
  nand g182155 (n_2673, g35, n_2957);
  nand g182146 (n_2476, g35, n_2796);
  nand g182143 (n_2690, g35, n_2766);
  nand g182132 (n_2482, g35, n_1705);
  not g182178 (n_1704, n_979);
  not g182220 (n_1703, n_8548);
  nand g182142 (n_1702, n_855, n_1569);
  nand g182021 (n_1701, n_328, n_304);
  nand g182019 (n_1700, n_1698, n_1699);
  nand g182018 (n_1697, g5575, g14694);
  nand g182013 (n_1696, g35, n_408);
  nand g182005 (n_1693, n_418, n_1692);
  not g182221 (n_1691, n_8551);
  nand g182003 (n_1690, new_g7704_, n_1506);
  not g182203 (n_1689, n_1720);
  nand g182000 (n_1688, g35, n_406);
  nand g181998 (n_1687, g35, n_361);
  nand g181997 (n_1686, g35, n_383);
  nand g181981 (n_1685, n_1608, n_313);
  not g182211 (n_1684, n_1867);
  not g182197 (n_1683, n_1724);
  not g182205 (n_1682, n_1706);
  nand g181979 (n_1681, g35, n_362);
  not g182186 (n_1680, n_1307);
  not g182202 (n_1679, n_1707);
  not g182184 (n_1678, n_1191);
  not g182182 (n_1677, n_1377);
  nand g181729 (n_1676, n_197, n_410);
  not g182183 (n_1675, n_517);
  not g182176 (n_1674, n_1007);
  not g182174 (n_1673, n_1015);
  not g182172 (n_1672, n_1023);
  not g182213 (n_1671, n_1763);
  nand g181978 (n_1670, g35, n_373);
  nand g181661 (n_1669, g13926, n_2609);
  not g182162 (n_1668, n_1086);
  not g182163 (n_1667, n_1084);
  nand g181655 (n_1666, g14828, n_2612);
  not g182156 (n_1665, n_1130);
  nand g181977 (n_1664, g5583, g14694);
  nand g181966 (n_1663, g3570, g13926);
  nor g181649 (n_1662, g1171, n_454);
  not g182157 (n_1661, n_1120);
  nand g181962 (n_1660, n_277, n_434);
  nand g182150 (n_1659, n_1378, n_1584);
  nand g181945 (n_1658, new_g10295_, n_316);
  nand g181631 (n_1656, n_1613, n_261);
  nand g181944 (n_1654, g5228, g14662);
  nand g181943 (n_1653, g35, n_407);
  nor g181620 (n_1652, n_1651, n_1610);
  not g182196 (n_1650, n_1710);
  nand g181940 (n_1649, g35, n_413);
  nand g181935 (n_1648, g3219, g13895);
  not g182181 (n_1647, n_1312);
  not g182170 (n_1646, n_1039);
  nand g181947 (n_1644, new_g7121_, n_1509);
  nand g181910 (n_1643, n_276, n_356);
  not g182969 (n_1642, n_1738);
  not g182891 (n_1641, n_699);
  nand g181968 (n_1640, g35, n_297);
  nand g181905 (n_1639, new_g7766_, n_1530);
  nand g181900 (n_1638, g35, n_353);
  nand g181898 (n_1637, g35, n_369);
  nor g181495 (n_1636, n_9257, n_386);
  nand g181897 (n_1635, n_319, n_293);
  nand g181528 (n_1634, g1236, n_9257);
  nand g181529 (n_1633, g347, n_9257);
  nor g181533 (n_1632, g1041, n_909);
  nand g181534 (n_1631, n_175, n_358);
  nand g181536 (n_1630, g1585, n_9257);
  nor g181539 (n_1629, g504, n_1554);
  nand g181542 (n_1628, g23683, n_9257);
  nor g181546 (n_1627, n_30, n_305);
  nor g181549 (n_1626, g4269, n_1625);
  nor g181552 (n_1623, g4452, g7260);
  nand g181554 (n_1622, g5236, n_6886);
  nand g181561 (n_1621, n_110, n_365);
  nor g181586 (n_1620, n_1055, n_357);
  nor g181588 (n_1619, n_1618, n_343);
  not g182947 (n_1617, n_1616);
  nor g181618 (n_1615, n_123, n_427);
  nor g181619 (n_1614, n_1613, n_364);
  nor g181622 (n_1612, g1430, n_1155);
  nor g181624 (n_1611, g370, n_1610);
  nor g181629 (n_1609, n_1608, n_274);
  nor g181632 (n_1607, g1087, n_1166);
  not g182948 (n_1606, n_1605);
  nor g181652 (n_1604, g5046, n_271);
  nand g181657 (n_1603, g14779, n_2614);
  nand g181658 (n_1602, g14738, n_1601);
  nand g181659 (n_1600, g14694, n_1599);
  nor g181673 (n_1598, g7916, g8416);
  nor g181675 (n_1597, g4878, n_1596);
  nand g181677 (n_1595, g13966, n_2621);
  nand g181678 (n_1594, g14662, n_1593);
  not g182946 (n_1592, n_1591);
  nand g182054 (n_1590, g1404, n_363);
  not g182943 (n_1589, n_1588);
  nand g181890 (n_1587, g35, n_370);
  nand g182052 (n_1586, g6267, g14779);
  nand g182051 (n_1585, new_g7812_, n_1584);
  nor g181584 (n_1583, n_29, n_425);
  nand g181994 (n_1582, g703, n_1581);
  nand g181580 (n_1580, g6275, n_6881);
  nand g181888 (n_1579, g6613, g14828);
  nand g181886 (n_1578, new_g10323_, n_1577);
  nand g181884 (n_1576, g3921, g13966);
  nand g181878 (n_1575, n_329, n_1581);
  nand g182012 (n_1574, n_368, n_1573);
  nand g181875 (n_1572, g35, n_256);
  nand g182017 (n_1571, g35, n_367);
  nand g181986 (n_1570, new_g7791_, n_1569);
  nor g181862 (n_1568, g4308, n_9257);
  not g181821 (n_1567, n_1566);
  nand g181989 (n_1565, g6621, g14828);
  nand g182002 (n_1564, n_345, n_394);
  not g182986 (n_2118, n_2359);
  not g181829 (n_2263, n_1563);
  not g181825 (n_2259, n_1562);
  nand g181780 (n_1712, g13272, n_1561);
  not g182201 (n_2131, n_1560);
  nand g181723 (n_2252, g4966, n_1559);
  nand g181721 (n_2014, g4776, n_1558);
  nand g181715 (n_4017, n_32, n_348);
  nand g182057 (n_2198, g890, n_269);
  not g182210 (n_6017, n_1557);
  nand g182134 (n_1883, n_1556, n_326);
  not g182963 (n_2070, n_1555);
  not g182987 (n_2093, n_2597);
  nand g181718 (n_1746, n_31, n_1554);
  not g181831 (n_2277, n_1553);
  not g182985 (n_2100, n_2631);
  not g182212 (n_5380, n_1552);
  nand g182141 (n_1718, n_1551, n_421);
  nand g182151 (n_1725, n_1550, n_290);
  nand g182136 (n_1884, n_1549, n_404);
  fflopd g990_reg(.CK (clock), .D (g8416), .Q (g990));
  not g182227 (n_2157, n_1850);
  nand g182091 (n_2580, g35, n_894);
  nand g182114 (n_2419, g35, n_1548);
  not g182236 (n_5120, n_1708);
  not g182235 (n_5083, n_1709);
  not g182241 (n_5076, n_1726);
  not g182997 (n_7035, n_2296);
  not g182239 (n_5181, n_1716);
  fflopd g4688_reg(.CK (clock), .D (g4681), .Q (g4688));
  not g182995 (n_6884, n_1547);
  not g182233 (n_5098, n_1546);
  not g182249 (n_5250, n_1545);
  not g182243 (n_5157, n_1544);
  not g182248 (n_4988, n_1543);
  not g182245 (n_5199, n_1542);
  not g182244 (n_5089, n_1541);
  not g182260 (n_5130, n_1540);
  fflopd g6704_reg(.CK (clock), .D (g14828), .Q (g17778));
  fflopd g5320_reg(.CK (clock), .D (g14662), .Q (g17674));
  not g182889 (n_1539, n_752);
  nand g182035 (n_1538, g35, n_379);
  nand g182040 (n_1537, n_431, n_262);
  nand g182044 (n_1536, g35, n_435);
  not g182180 (n_1535, n_653);
  nand g181903 (n_1534, g35, n_388);
  nand g182050 (n_1533, g35, n_389);
  nand g182053 (n_1532, g35, n_401);
  nand g182140 (n_1531, n_1309, n_1530);
  not g182185 (n_1529, n_1265);
  nand g182070 (n_1528, g4628, n_1527);
  fflopd g4477_reg(.CK (clock), .D (new_g12875_), .Q (g4477));
  nand g181537 (n_1526, g1579, n_9257);
  nand g182020 (n_1525, new_g7738_, n_1500);
  nand g181889 (n_1523, g35, n_440);
  nand g181887 (n_1522, g4831, g4681);
  not g182187 (n_1521, n_1362);
  not g182189 (n_1520, n_1519);
  not g182173 (n_1518, n_577);
  nand g181674 (n_1517, g13895, n_1516);
  nand g182029 (n_1515, g5929, g14738);
  not g182165 (n_1514, n_1080);
  nand g181595 (n_1513, n_473, n_1512);
  not g182171 (n_1511, n_848);
  nand g182135 (n_1510, n_1158, n_1509);
  not g182195 (n_1508, n_1722);
  nand g182138 (n_1507, n_880, n_1506);
  nand g181538 (n_1505, n_162, n_366);
  nand g182034 (n_1504, g35, n_320);
  nand g182046 (n_1503, g5084, n_395);
  nand g182043 (n_1502, g35, n_400);
  nand g182152 (n_1501, n_745, n_1500);
  nand g182153 (n_1499, n_910, n_1577);
  not g182158 (n_1498, n_1115);
  not g182160 (n_1497, n_1100);
  not g182164 (n_1496, n_1082);
  not g182168 (n_1495, n_1051);
  not g182169 (n_1494, n_1048);
  not g182175 (n_1493, n_1012);
  not g182177 (n_1492, n_581);
  not g182179 (n_1491, n_977);
  not g182188 (n_1490, n_1489);
  not g182190 (n_1488, n_1487);
  nand g182056 (n_1486, g5921, g14738);
  not g182194 (n_1485, n_1892);
  not g182199 (n_1484, n_1715);
  not g182200 (n_1483, n_1721);
  nor g181545 (n_1482, g5097, n_1481);
  not g182206 (n_1480, n_1803);
  not g182159 (n_1479, n_1111);
  nor g181558 (n_1478, g4633, n_1527);
  not g182886 (n_1477, n_785);
  not g182219 (n_1476, n_8550);
  not g182890 (n_1475, n_744);
  not g182225 (n_1474, n_3378);
  not g182226 (n_1473, n_7970);
  not g182893 (n_1472, n_667);
  not g182892 (n_1471, n_1398);
  not g182894 (n_1470, n_665);
  not g182896 (n_1469, n_519);
  not g182898 (n_1468, n_878);
  not g182888 (n_1467, n_1308);
  not g182887 (n_1466, n_758);
  not g182965 (n_1465, n_1780);
  not g182247 (n_1464, n_5346);
  not g182958 (n_1463, n_8116);
  not g182954 (n_1462, n_1853);
  not g182949 (n_1461, n_1460);
  not g182942 (n_1457, n_1456);
  not g182941 (n_1455, n_1454);
  not g182931 (n_1453, n_1452);
  not g182897 (n_1451, n_654);
  not g182895 (n_1450, n_510);
  nand g182033 (n_1449, g35, n_415);
  not g182885 (n_1448, n_788);
  not g182884 (n_1447, n_613);
  not g181827 (n_2261, n_1446);
  not g182979 (n_2091, n_2457);
  nand g182066 (n_2000, n_1445, n_416);
  nand g182074 (n_2002, g35, n_359);
  not g181826 (n_2266, n_1444);
  not g182223 (n_2136, n_8549);
  not g181828 (n_2272, n_1443);
  nand g182133 (n_1714, n_1442, n_266);
  nand g182137 (n_1717, n_1441, n_286);
  nand g182139 (n_1885, n_1440, n_303);
  not g182962 (n_2127, n_1439);
  nand g182145 (n_1888, n_1438, n_444);
  not g182966 (n_2142, n_1437);
  not g182967 (n_2039, n_1436);
  not g182972 (n_2202, n_1435);
  not g182975 (n_2040, n_2032);
  wire w227, w228, w229, w230;
  nand g182148 (n_1887, w228, w230);
  nand g257 (w230, w229, g979);
  not g256 (w229, n_1434);
  nand g254 (w228, w227, n_1434);
  not g253 (w227, g979);
  not g182981 (n_2096, n_2623);
  not g182982 (n_2105, n_2497);
  not g182984 (n_2111, n_2626);
  not g182983 (n_2116, n_2475);
  wire w231, w232, w233, w234;
  nand g182149 (n_1719, w232, w234);
  nand g261 (w234, w233, g1322);
  not g260 (w233, n_1433);
  nand g259 (w232, w231, n_1433);
  not g258 (w231, g1322);
  not g182204 (n_2717, n_1432);
  nand g182063 (n_1998, g35, n_360);
  nand g182065 (n_2016, n_1324, n_1355);
  not g182208 (n_2933, n_1431);
  not g181830 (n_2274, n_1430);
  not g182209 (n_2826, n_1429);
  not g182214 (n_2124, n_1428);
  not g182216 (n_5379, n_1427);
  not g182228 (n_4319, n_2544);
  not g182222 (n_2133, n_8546);
  nand g182087 (n_5035, g35, n_424);
  not g182230 (g25167, n_1426);
  nand g182094 (n_2677, g35, n_1425);
  not g182231 (n_8568, n_1424);
  nand g182115 (n_2559, g35, n_895);
  not g182238 (n_5163, n_1723);
  not g182240 (n_5051, n_1727);
  not g182242 (n_5208, n_1713);
  nand g182120 (n_2462, g35, n_897);
  nand g182125 (n_2444, g35, n_898);
  not g182994 (n_6888, n_2294);
  not g182257 (n_3767, n_5464);
  not g182992 (n_7031, n_2325);
  not g182980 (n_4646, n_1423);
  nand g182123 (n_2666, g35, n_1422);
  not g182237 (n_5212, n_1711);
  nand g182109 (n_2465, g35, n_1421);
  nand g182093 (n_2480, g35, n_1420);
  not g182256 (n_3769, n_5462);
  nand g182119 (n_2413, g35, n_1419);
  not g182265 (n_3773, n_5466);
  nand g182112 (n_2411, g35, n_449);
  nand g182110 (n_2681, g35, n_1418);
  nand g182106 (n_2384, g35, n_446);
  nand g182096 (n_2436, g35, n_1417);
  nand g182103 (n_2416, g35, n_447);
  nand g182100 (n_2499, g35, n_893);
  not g182234 (n_5039, n_1416);
  not g182264 (n_6450, n_3616);
  not g182259 (n_4168, n_4831);
  not g182258 (n_5126, n_2996);
  not g182246 (n_5186, n_1415);
  not g182252 (n_5047, n_1414);
  not g182266 (n_4952, n_6159);
  not g182263 (n_6454, n_3614);
  not g182996 (n_5789, n_1413);
  not g182250 (n_5145, n_1412);
  not g182254 (n_5758, n_4444);
  not g182261 (n_4922, n_1411);
  fflopd g5666_reg(.CK (clock), .D (g14694), .Q (g17711));
  fflopd g3661_reg(.CK (clock), .D (g13926), .Q (g16744));
  fflopd g6358_reg(.CK (clock), .D (g14779), .Q (g17760));
  fflopd g6012_reg(.CK (clock), .D (g14738), .Q (g17739));
  fflopd g4012_reg(.CK (clock), .D (g13966), .Q (g16775));
  fflopd g3310_reg(.CK (clock), .D (g13895), .Q (g16718));
  not g182262 (n_5128, n_1410);
  not g182253 (n_5760, n_1409);
  not g182255 (n_6456, n_823);
  nand g182737 (n_1408, g25219, n_9257);
  nand g183255 (n_1407, g3965, n_9257);
  nand g183302 (n_1406, g35, n_6357);
  nand g182460 (n_1405, g2629, n_9257);
  nand g182712 (n_1404, g1854, n_9257);
  nand g182661 (n_1403, g5228, n_9257);
  nand g182273 (n_1402, g4417, n_9257);
  nand g182531 (n_1401, g4878, n_181);
  nand g182589 (n_1400, g671, n_9257);
  nand g182345 (n_1399, g4864, n_146);
  nand g183193 (n_1398, g4382, n_9257);
  nand g183294 (n_1397, n_9257, n_72);
  nand g182732 (n_1396, g2495, n_9257);
  not g182198 (n_1395, g4291);
  nand g183119 (n_1394, g703, n_9257);
  nand g182729 (n_1393, g6593, n_9257);
  nand g182594 (n_1392, g6267, n_9257);
  nand g183026 (n_1391, g1632, n_9257);
  nand g182672 (n_1390, g5937, n_9257);
  nand g183259 (n_1389, g6633, n_9257);
  nand g182727 (n_1388, g2269, n_9257);
  nand g183257 (n_1387, g5527, n_9257);
  nand g182427 (n_1386, g3905, n_9257);
  nand g182439 (n_1385, new_g6905_, n_9257);
  nand g182706 (n_1384, g2472, n_9257);
  nand g182596 (n_1383, g2236, n_9257);
  nand g182436 (n_1382, g1430, n_1381);
  nand g182421 (n_1380, g1612, n_9257);
  not g182924 (n_1379, n_1378);
  nand g182597 (n_1377, g4153, n_9257);
  not g182215 (n_1376, n_1934);
  nand g183260 (n_1375, g2012, n_9257);
  not g182207 (n_1374, g4281);
  nand g182683 (n_1373, g2988, n_9257);
  nand g182417 (n_1372, g6203, n_9257);
  nand g183191 (n_1371, g4297, n_9257);
  nand g182725 (n_1370, g1532, n_9257);
  nand g183256 (n_1369, g2066, n_9257);
  not g182920 (n_1368, n_1367);
  nand g182721 (n_1366, g2020, n_9257);
  nand g182591 (n_1365, g6601, n_9257);
  nand g182577 (n_1364, g5893, n_9257);
  nand g182592 (n_1363, new_g6928_, n_9257);
  nand g182717 (n_1362, g153, n_9257);
  nand g182560 (n_1361, g5941, n_9257);
  nand g183112 (n_1360, g6209, n_9257);
  nand g182675 (n_1359, g6259, n_9257);
  nand g183232 (n_1358, g2555, n_9257);
  not g182956 (n_1357, n_1417);
  nand g183074 (n_1354, g4119, n_9257);
  nand g182399 (n_1351, g1061, n_1350);
  nand g183189 (n_1349, g4245, n_9257);
  nand g183338 (n_1348, g35, n_1347);
  nand g182685 (n_1346, g5406, n_9257);
  not g182964 (n_1345, n_1419);
  nand g183334 (n_1344, n_9257, n_52);
  nand g182276 (n_1343, g6533, n_9257);
  nand g183108 (n_1342, g191, n_9257);
  nand g182715 (n_1341, g2894, n_9257);
  nand g183106 (n_1340, g4180, n_9257);
  nand g182315 (n_1339, g269, n_9257);
  nand g183204 (n_1338, g5264, n_9257);
  nand g182666 (n_1337, new_g7028_, n_9257);
  nand g183102 (n_1336, g681, n_9257);
  nand g183181 (n_1335, g3219, n_9257);
  nand g183241 (n_1334, g1825, n_9257);
  nand g183176 (n_1333, g5752, n_9257);
  nand g183177 (n_1332, g6727, n_9257);
  nand g182556 (n_1331, g5240, n_9257);
  nand g182713 (n_1330, g1178, n_9257);
  nand g182736 (n_1329, g2445, n_9257);
  nand g182519 (n_1328, g1936, n_9257);
  nand g183273 (n_1327, g1648, n_9257);
  nand g182413 (n_1326, g3538, n_9257);
  nand g182711 (n_1323, g1744, n_9257);
  nand g183090 (n_1322, g2250, n_9257);
  nand g182709 (n_1321, g2980, n_9257);
  not g182973 (n_1320, n_1420);
  nand g183082 (n_1319, g3115, n_9257);
  nand g183309 (n_1318, n_1030, n_1317);
  nand g182705 (n_1316, g2657, n_9257);
  nand g182731 (n_1315, g2342, n_9257);
  nand g182733 (n_1314, g2518, n_9257);
  nand g182582 (n_1313, g5180, n_9257);
  nand g182576 (n_1312, g5092, n_9257);
  nand g182336 (n_1311, g3462, n_9257);
  not g182928 (n_1310, n_1309);
  nand g183070 (n_1308, g4057, n_9257);
  nand g182701 (n_1307, g772, n_9257);
  nand g182407 (n_1306, g1687, n_9257);
  nand g182699 (n_1305, g6597, n_9257);
  nand g183229 (n_1304, g4249, n_9257);
  nand g182291 (n_1303, g5881, n_9257);
  nand g183277 (n_1302, g2208, n_9257);
  nand g183269 (n_1301, g1752, n_9257);
  nand g182511 (n_1300, g4793, n_1299);
  not g182933 (n_1298, n_1297);
  nand g182304 (n_1296, g5252, n_9257);
  nand g183253 (n_1295, g2429, n_9257);
  nand g183249 (n_1294, g3841, n_9257);
  nand g183133 (n_1293, g3263, n_9257);
  nand g182697 (n_1292, g2815, n_9257);
  nand g183237 (n_1291, g5268, n_9257);
  nand g183225 (n_1290, g324, n_9257);
  nand g183231 (n_1289, g2357, n_9257);
  nand g182319 (n_1288, g1178, n_130);
  nand g183217 (n_1287, g2848, n_9257);
  nand g182312 (n_1286, g3562, n_9257);
  nand g182314 (n_1285, g3554, n_9257);
  wire w235, w236, w237, w238;
  nand g182069 (n_1284, w236, w238);
  nand g266 (w238, w237, g232);
  not g265 (w237, g225);
  nand g264 (w236, w235, g225);
  not g263 (w235, g232);
  nand g183201 (n_1283, g2193, n_9257);
  nand g183197 (n_1282, g962, n_9257);
  nand g183195 (n_1281, g2223, n_9257);
  nand g183185 (n_1280, g3917, n_9257);
  nand g183175 (n_1279, g5897, n_9257);
  nand g183173 (n_1278, g5595, n_9257);
  nand g183169 (n_1277, g5037, n_9257);
  nand g182545 (n_1276, g2070, n_9257);
  nand g182404 (n_1275, g2384, n_85);
  nand g183159 (n_1274, g2579, n_9257);
  nand g183161 (n_1273, g1141, n_9257);
  nand g182296 (n_1272, g6625, n_9257);
  nand g183147 (n_1271, g4515, n_9257);
  nand g183152 (n_1270, g6573, n_9257);
  nand g183151 (n_1269, g2227, n_9257);
  nand g183143 (n_1268, g3171, n_9257);
  nand g183144 (n_1267, g832, n_9257);
  nand g183141 (n_1266, g1798, n_9257);
  nand g182695 (n_1265, g1542, n_9257);
  nand g183137 (n_1264, g3578, n_9257);
  nand g182283 (n_1263, g1974, n_9257);
  nand g182693 (n_1262, g3558, n_9257);
  nand g182516 (n_1261, g4983, n_1260);
  nand g182570 (n_1259, g5909, n_9257);
  nand g182723 (n_1258, g3925, n_9257);
  nand g183128 (n_1257, g4593, n_9257);
  nand g182272 (n_1256, g446, n_9257);
  nand g183127 (n_1255, g2791, n_9257);
  nand g183125 (n_1254, g3231, n_9257);
  nand g183123 (n_1253, new_g7051_, n_9257);
  nand g183116 (n_1252, g3347, n_9257);
  nor g183118 (n_1251, g35, n_3986);
  nand g183114 (n_1250, g1124, n_9257);
  nand g182268 (n_1249, g5957, n_9257);
  nand g182571 (n_1248, g2803, n_9257);
  nand g182726 (n_1247, g2169, n_9257);
  nand g182579 (n_1246, g6509, n_9257);
  nand g183104 (n_1245, g3199, n_9257);
  nand g183105 (n_1244, g5913, n_9257);
  nand g183050 (n_1243, g5579, n_9257);
  nand g183092 (n_1242, g1521, n_9257);
  nand g183096 (n_1241, g5933, n_9257);
  nand g183094 (n_1240, g2779, n_9257);
  nand g183086 (n_1239, g1830, n_9257);
  nand g183078 (n_1238, g6271, n_9257);
  nand g183079 (n_1237, g4172, n_9257);
  not g182899 (n_1236, n_285);
  nand g183068 (n_1235, g1844, n_9257);
  nand g182691 (n_1234, g2537, n_9257);
  nand g183058 (n_1233, g3606, n_9257);
  nand g183062 (n_1232, g5535, n_9257);
  nand g183056 (n_1231, g3582, n_9257);
  nand g183048 (n_1230, g1955, n_9257);
  nand g183038 (n_1229, g2380, n_9257);
  nand g183031 (n_1228, g6239, n_9257);
  nand g183032 (n_1227, g6311, n_9257);
  nand g183022 (n_1226, g1691, n_9257);
  nand g183018 (n_1225, g3129, n_9257);
  nand g182690 (n_1224, g2907, n_9257);
  nand g182689 (n_1223, g1792, n_9257);
  nand g183010 (n_1222, g1748, n_9257);
  nand g182684 (n_1221, g1840, n_9257);
  nand g182678 (n_1220, g1189, n_9257);
  not g182970 (n_1219, n_1596);
  nor g182397 (n_1218, g5097, n_27);
  nand g182676 (n_1215, g1592, n_9257);
  nand g182674 (n_1214, g5563, n_9257);
  nand g182494 (n_1213, new_g8038_, n_9257);
  nand g182518 (n_1212, n_906, n_2866);
  not g182910 (n_1211, n_327);
  not g182913 (n_1210, n_324);
  not g182952 (n_1208, n_1548);
  nand g183042 (n_1207, g2024, n_9257);
  nand g182670 (n_1206, g2563, n_9257);
  nand g182668 (n_1205, g2093, n_9257);
  nand g182667 (n_1204, g542, n_9257);
  nand g182664 (n_1202, g1211, n_9257);
  nand g182662 (n_1201, g5587, n_9257);
  nand g183149 (n_1200, g4358, n_9257);
  nand g182658 (n_1199, g6657, n_9257);
  nand g182656 (n_1198, g1437, n_9257);
  nand g182565 (n_1197, g1454, n_9257);
  nand g182655 (n_1196, g6390, n_9257);
  nand g182568 (n_1195, g1351, n_9257);
  nand g183297 (n_1194, n_470, n_905);
  nand g182654 (n_1193, g1094, n_9257);
  nand g182650 (n_1192, g2671, n_9257);
  nand g182687 (n_1191, g4264, n_9257);
  nand g182375 (n_1190, g1536, n_9257);
  nand g182648 (n_1189, g2441, n_9257);
  nor g182646 (n_1188, g35, n_6814);
  nand g182644 (n_1187, g3480, n_9257);
  not g182971 (n_1186, n_1421);
  not g182934 (n_1185, n_436);
  nand g182722 (n_1184, g3191, n_9257);
  nand g183292 (n_1183, g6275, n_9257);
  not g182902 (n_1182, n_284);
  nand g182719 (n_1181, g5841, n_9257);
  nand g182718 (n_1180, g2303, n_9257);
  nand g182716 (n_1179, g3512, n_9257);
  nand g182714 (n_1178, g6243, n_9257);
  nand g182694 (n_1177, g2912, n_9257);
  nand g182707 (n_1176, g2384, n_9257);
  nand g182708 (n_1175, g2311, n_9257);
  nor g182383 (n_1174, g411, n_1173);
  wire w239, w240, w241, w242;
  nand g181879 (n_1172, w240, w242);
  nand g271 (w242, w241, g182);
  not g270 (w241, g452);
  nand g268 (w240, w239, g452);
  not g267 (w239, g182);
  nand g182657 (n_1171, g5921, n_9257);
  nand g182704 (n_1170, g4273, n_9257);
  nand g182700 (n_1169, g2941, n_9257);
  nand g182555 (n_1168, g3941, n_9257);
  not g182923 (n_1167, n_1166);
  nand g183337 (n_1165, g35, n_617);
  wire w243, w244, w245, w246;
  nand g181874 (n_1164, w244, w246);
  nand g275 (w246, w245, g661);
  not g274 (w245, g728);
  nand g273 (w244, w243, g728);
  not g272 (w243, g661);
  nand g183054 (n_1163, g2827, n_9257);
  wire w247, w248, w249, w250;
  nand g181880 (n_1162, w248, w250);
  nand g280 (w250, w249, g358);
  not g279 (w249, g376);
  nand g277 (w248, w247, g376);
  not g276 (w247, g358);
  wire w251, w252, w253, w254;
  nand g181881 (n_1161, w252, w254);
  nand g285 (w254, w253, g392);
  not g284 (w253, g405);
  nand g282 (w252, w251, g405);
  not g281 (w251, g392);
  nand g182550 (n_1160, g2606, n_9257);
  not g182927 (n_1159, n_1158);
  wire w255, w256, w257, w258;
  nand g181891 (n_1157, w256, w258);
  nand g290 (w258, w257, g718);
  not g289 (w257, g655);
  nand g288 (w256, w255, g655);
  not g286 (w255, g718);
  not g182929 (n_1156, n_1155);
  nand g182660 (n_1154, g1913, n_9257);
  nand g182641 (n_1153, g2771, n_9257);
  nand g182698 (n_1152, g3155, n_9257);
  nand g183012 (n_1151, g2652, n_9257);
  nand g182558 (n_1150, g5599, n_9257);
  not g182921 (n_1149, n_1148);
  nand g182612 (n_1147, g2389, n_9257);
  nand g182703 (n_1146, g2960, n_9257);
  nand g182643 (n_1145, g3913, n_9257);
  nand g182640 (n_1144, g996, n_9257);
  nand g182692 (n_1143, g2902, n_9257);
  nand g182639 (n_1142, g5248, n_9257);
  nand g182688 (n_1141, g142, n_9257);
  nand g182369 (n_1140, g2250, n_23);
  not g182917 (n_1139, n_306);
  not g182192 (n_1138, g4452);
  nand g182269 (n_1137, g2338, n_9257);
  nand g182270 (n_1136, g3752, n_9257);
  nand g182271 (n_1135, g1339, n_9257);
  nand g183238 (n_1134, g5138, n_9257);
  nand g182277 (n_1133, g1135, n_9257);
  nor g182526 (n_1132, g4035, n_1994);
  nand g182279 (n_1131, g1720, n_9257);
  nand g182280 (n_1130, g794, n_9257);
  nand g182281 (n_1129, g5511, n_9257);
  nand g182282 (n_1128, g1886, n_9257);
  nand g182573 (n_1127, g5567, n_9257);
  nand g182286 (n_1126, g262, n_9257);
  nand g182287 (n_1125, g3546, n_9257);
  nand g182288 (n_1124, g2060, n_9257);
  nand g182681 (n_1123, g2856, n_9257);
  nand g182292 (n_1122, g2844, n_9257);
  nand g182293 (n_1121, g6609, n_9257);
  nand g182294 (n_1120, g291, n_9257);
  nand g182295 (n_1119, g3574, n_9257);
  nand g182297 (n_1118, g6291, n_9257);
  nand g182298 (n_1117, g5551, n_9257);
  nand g182301 (n_1116, new_g7074_, n_9257);
  nand g182302 (n_1115, g1199, n_9257);
  nand g182535 (n_1114, g2823, n_9257);
  nand g182308 (n_1113, g6235, n_9257);
  nand g182309 (n_1112, g5615, n_9257);
  nand g182310 (n_1111, g298, n_9257);
  nand g182311 (n_1110, g6251, n_9257);
  nand g182313 (n_1109, g2299, n_9257);
  nand g182323 (n_1106, g1668, n_9257);
  nand g182324 (n_1105, g6549, n_9257);
  nand g182327 (n_1103, g1521, n_232);
  nand g182331 (n_1101, g4849, n_20);
  nand g182334 (n_1100, g4382, n_1099);
  nand g182337 (n_1097, g6641, n_9257);
  nand g182339 (n_1095, g4076, n_626);
  nand g182680 (n_1094, g278, n_9257);
  nor g182341 (n_1093, g4269, n_242);
  nand g182342 (n_1092, g4659, n_190);
  nand g182679 (n_1091, g1472, n_9257);
  not g182901 (n_1090, n_322);
  nand g182355 (n_1086, g2514, n_1085);
  nand g182356 (n_1084, g2648, n_1083);
  nand g182357 (n_1082, g1821, n_1081);
  nand g182358 (n_1080, g1955, n_1079);
  nand g182362 (n_1076, new_g10354_, n_230);
  nand g182367 (n_1075, g1959, n_235);
  nand g182368 (n_1074, g20899, n_223);
  nand g182371 (n_1073, g2518, n_196);
  nand g182372 (n_1072, g2652, n_200);
  nand g182374 (n_1071, g1825, n_34);
  nand g182677 (n_1070, g1379, n_9257);
  nand g182378 (n_1069, g691, n_9257);
  nand g182380 (n_1068, g1691, n_192);
  nand g182386 (n_1067, g4264, n_139);
  nand g182387 (n_1066, g2421, n_9257);
  nand g182389 (n_1065, g1564, n_215);
  not g182911 (n_1064, n_263);
  nand g182396 (n_1063, g2173, n_9257);
  nand g182673 (n_1062, g2864, n_9257);
  nand g182406 (n_1061, g1988, n_9257);
  nor g182409 (n_1060, g405, n_1059);
  nand g182671 (n_1058, g1367, n_9257);
  nand g182410 (n_1057, g1862, n_9257);
  nor g182411 (n_1056, g1030, n_1055);
  nand g182412 (n_1054, g667, n_9257);
  nand g182414 (n_1053, g1748, n_7);
  nand g182415 (n_1052, g2575, n_211);
  nand g182416 (n_1051, g10500, n_1050);
  nand g182418 (n_1049, g546, n_9257);
  nand g182419 (n_1048, g2089, n_1047);
  nand g182420 (n_1046, g1644, n_9257);
  nand g182422 (n_1045, g2413, n_9257);
  nor g182359 (n_1044, g827, n_1043);
  nand g182424 (n_1042, g2047, n_9257);
  nor g182425 (n_1041, g5029, n_1040);
  nand g182426 (n_1039, g744, n_9257);
  nand g182428 (n_1038, g6247, n_9257);
  nand g182429 (n_1037, g5467, n_9257);
  nand g182430 (n_1036, g4643, n_9257);
  nand g182431 (n_1035, g3050, n_9257);
  nand g182433 (n_1034, g5965, n_9257);
  nand g182434 (n_1033, g5961, n_9257);
  nand g182435 (n_1032, g518, n_9257);
  nor g182438 (n_1031, g1906, n_1030);
  nand g182440 (n_1029, g6505, n_9257);
  nand g182441 (n_1028, g2093, n_179);
  nand g182442 (n_1027, g5092, n_1026);
  nand g182443 (n_1025, g6381, n_9257);
  nand g182696 (n_1024, g6613, n_9257);
  nand g182446 (n_1023, g2975, n_9257);
  nand g182450 (n_1022, g1600, n_9257);
  nand g182451 (n_1021, g37, n_9257);
  nand g182408 (n_1020, g10527, n_1019);
  nand g182453 (n_1018, g1882, n_903);
  nand g182455 (n_1017, g2173, n_451);
  nand g182457 (n_1016, g6555, n_9257);
  nand g182458 (n_1015, g1612, n_453);
  nand g182459 (n_1014, g2016, n_480);
  nand g182462 (n_1013, g3937, n_9257);
  nand g182464 (n_1012, g2331, n_1011);
  nand g182465 (n_1010, g1608, n_1009);
  nand g182466 (n_1008, g5689, n_9257);
  nand g182467 (n_1007, g837, n_3916);
  nor g182469 (n_1006, g2599, n_1005);
  nand g182470 (n_1004, g5471, n_9257);
  not g182960 (n_1003, n_2290);
  nand g182473 (n_1002, g5905, n_9257);
  nand g182476 (n_1001, g5120, n_9257);
  nand g182477 (n_1000, g3338, n_9257);
  nor g182479 (n_999, g4991, n_998);
  nand g182482 (n_997, g3207, n_9257);
  nand g182483 (n_996, g847, n_9);
  nand g182485 (n_995, g6219, n_9257);
  nor g182486 (n_994, g5016, n_1916);
  nor g182487 (n_993, g4515, n_3509);
  nand g182489 (n_992, g12923, n_37);
  nand g182490 (n_991, g2361, n_9257);
  nor g182491 (n_990, g4801, n_136);
  nand g182638 (n_989, g2437, n_9257);
  nand g183233 (n_988, g3550, n_9257);
  nand g182497 (n_987, g534, n_9257);
  nand g182501 (n_986, g4483, n_9257);
  nand g182503 (n_985, g890, n_9257);
  nand g182505 (n_984, g5889, n_9257);
  nor g182506 (n_983, g2040, n_982);
  nand g182507 (n_981, g5857, n_9257);
  nand g182509 (n_980, g2579, n_978);
  nand g182512 (n_979, g2571, n_978);
  nand g182513 (n_977, g781, n_9257);
  nand g182514 (n_976, g2437, n_975);
  nand g182517 (n_974, g209, n_9257);
  nand g182521 (n_973, g2950, n_9257);
  nand g182522 (n_972, g4443, n_9257);
  not g182907 (n_971, n_331);
  nand g182524 (n_970, g3259, n_9257);
  nand g182525 (n_969, g3530, n_968);
  nand g182527 (n_967, g283, n_9257);
  nand g182528 (n_966, g1008, n_103);
  nand g182529 (n_965, g3179, n_9257);
  nand g182530 (n_964, g4776, n_9257);
  nand g182532 (n_963, g4584, n_962);
  nand g182533 (n_961, g1932, n_9257);
  nand g182665 (n_960, g4340, n_9257);
  nand g182536 (n_959, g2795, n_9257);
  nand g182539 (n_958, g358, n_957);
  nor g182543 (n_956, new_g10354_, n_4542);
  nand g182637 (n_955, g437, n_9257);
  not g182218 (n_954, n_1955);
  nand g182546 (n_953, g3161, n_9257);
  nand g182549 (n_952, g5945, n_9257);
  nand g182551 (n_951, g5543, n_9257);
  nand g182552 (n_950, g3227, n_9257);
  nand g182554 (n_949, g5485, n_9257);
  nand g182557 (n_948, g2783, n_9257);
  nand g182561 (n_947, g3929, n_9257);
  nand g182562 (n_946, g1105, n_9257);
  nand g182564 (n_945, g168, n_9257);
  nand g182567 (n_944, g3901, n_9257);
  nand g182569 (n_943, g3957, n_9257);
  nand g182572 (n_942, g5124, n_9257);
  nand g182574 (n_941, g4633, n_9257);
  nand g182575 (n_940, g5603, n_9257);
  nand g182578 (n_939, g6617, n_9257);
  nand g182580 (n_938, g822, n_9257);
  nand g182581 (n_937, g6585, n_9257);
  nand g182583 (n_936, g385, n_9257);
  not g182906 (n_935, n_339);
  nand g182586 (n_934, g4040, n_9257);
  nand g182590 (n_933, g5495, n_9257);
  nand g182593 (n_932, g2485, n_9257);
  nand g182595 (n_931, g4388, n_9257);
  nand g182598 (n_930, g4621, n_9257);
  nand g182599 (n_929, g2999, n_9257);
  nand g182600 (n_928, g5925, n_9257);
  nand g182603 (n_927, g5619, n_9257);
  nand g182604 (n_926, g20652, n_9257);
  nand g182610 (n_925, new_g7004_, n_9257);
  nand g182611 (n_924, g5698, n_9257);
  nand g182616 (n_923, g3893, n_9257);
  nand g182617 (n_922, g2449, n_9257);
  nand g182618 (n_921, g5607, n_9257);
  nand g182620 (n_920, g2403, n_9257);
  nand g182626 (n_919, g6177, n_9257);
  nand g182627 (n_918, g5813, n_9257);
  nand g182629 (n_917, g3590, n_9257);
  nand g182630 (n_916, g1706, n_9257);
  nand g182633 (n_915, g3889, n_9257);
  nand g182859 (n_1545, new_g6928_, n_907);
  not g182950 (n_1966, n_914);
  wire w259, w260, w261, w262;
  nand g182084 (n_1563, w260, w262);
  nand g296 (w262, w261, g4040);
  not g295 (w261, g11418);
  nand g293 (w260, w259, g11418);
  not g292 (w259, g4040);
  wire w263, w264, w265, w266;
  nand g182081 (n_1444, w264, w266);
  nand g302 (w266, w265, g5689);
  not g300 (w265, g12300);
  nand g299 (w264, w263, g12300);
  not g297 (w263, g5689);
  wire w267, w268, w269, w270;
  nand g182064 (n_3758, w268, w270);
  nand g307 (w270, w269, g8358);
  not g306 (w269, g191);
  nand g304 (w268, w267, g191);
  not g303 (w267, g8358);
  wire w271, w272, w273, w274;
  nand g182073 (n_1566, w272, w274);
  nand g312 (w274, w273, g3689);
  not g310 (w273, g11388);
  nand g309 (w272, w271, g11388);
  not g308 (w271, g3689);
  nand g183583 (n_1435, n_912, n_913);
  nand g182796 (n_1552, g2599, n_134);
  nor g183566 (n_1984, g890, n_9257);
  nand g183565 (n_1439, g35, n_2866);
  nand g183530 (n_1588, g35, n_49);
  not g182938 (n_1948, n_398);
  nand g182743 (n_1519, g2465, n_911);
  nand g183538 (n_1591, g35, n_2376);
  not g182968 (n_1890, n_910);
  not g182961 (n_4143, n_909);
  not g182974 (n_1732, n_2227);
  nand g183613 (n_1413, n_907, n_908);
  not g182232 (n_3197, new_g7717_);
  nand g182773 (n_1707, g3873, n_599);
  nand g183587 (n_2032, g35, n_135);
  nor g182804 (n_1894, new_g10795_, n_906);
  nand g182774 (n_2761, g5881, n_905);
  nand g182835 (n_1709, g5511, n_47);
  nand g182841 (n_1726, g6549, n_16);
  nand g182839 (n_1716, g3857, n_17);
  nand g182843 (n_1713, g5164, n_212);
  nand g183608 (n_2325, n_475, n_904);
  nor g183571 (n_1920, g4349, n_9257);
  nand g182817 (n_8549, g1917, n_903);
  nand g182761 (n_1724, g3171, n_816);
  nand g183599 (n_2475, g35, n_1551);
  not g182978 (n_2856, n_412);
  not g182991 (n_3272, n_3789);
  nand g183601 (n_2631, g35, n_1556);
  nand g182871 (n_5464, g5297, n_902);
  nand g182879 (n_5466, new_g10366_, n_901);
  nor g183588 (n_4343, n_479, n_450);
  not g182993 (n_5150, n_900);
  not g183000 (n_3627, n_899);
  not g183006 (n_5197, n_898);
  not g182989 (n_5170, n_897);
  not g183007 (n_5154, n_896);
  not g183003 (n_5160, n_895);
  not g183002 (n_5220, n_894);
  not g182990 (n_5193, n_893);
  not g182999 (n_5152, n_892);
  nand g182844 (n_6011, n_59, n_3496);
  nand g183263 (n_891, g1902, n_9257);
  nand g182740 (n_890, g2165, n_9257);
  nand g182741 (n_889, g1448, n_9257);
  nand g182738 (n_888, g5917, n_9257);
  nand g182468 (n_887, g336, n_9257);
  nand g182587 (n_886, g2648, n_9257);
  nand g182448 (n_885, g2307, n_452);
  not g182904 (n_884, n_292);
  nand g183207 (n_883, g3961, n_9257);
  nand g183203 (n_882, g4785, n_9257);
  not g182936 (n_881, n_880);
  nand g183264 (n_879, g2246, n_9257);
  nand g183266 (n_878, g4064, n_9257);
  nand g183046 (n_877, g3111, n_9257);
  nand g183308 (n_876, n_3691, n_3509);
  not g182955 (n_875, n_1418);
  nand g182474 (n_874, g3235, n_9257);
  nand g182267 (n_872, g2204, n_9257);
  nand g183208 (n_871, g2476, n_9257);
  nand g182720 (n_870, g6581, n_9257);
  nand g183030 (n_869, g4849, n_9257);
  nand g182606 (n_868, g3945, n_9257);
  nand g182452 (n_867, g2327, n_9257);
  nand g182605 (n_866, g3817, n_9257);
  not g182957 (n_865, n_1699);
  nand g182449 (n_864, g2441, n_463);
  nand g182480 (n_863, g2351, n_9257);
  nand g182423 (n_862, g1087, n_99);
  nand g183199 (n_861, g5256, n_9257);
  nand g182601 (n_860, g5170, n_9257);
  nor g182608 (n_859, g35, n_858);
  nand g182454 (n_857, g3251, n_9257);
  not g182918 (n_856, n_855);
  nand g182275 (n_854, g3211, n_9257);
  nand g182607 (n_853, g4975, n_9257);
  nand g182278 (n_852, g3614, n_9257);
  nand g182437 (n_851, g4116, n_9257);
  not g182193 (n_850, n_849);
  nand g182445 (n_848, g2599, n_1005);
  nand g182274 (n_847, g699, n_9257);
  nand g183153 (n_846, g1878, n_9257);
  nand g183024 (n_845, g6736, n_9257);
  nand g182602 (n_844, g4311, n_9257);
  nand g183211 (n_843, g2036, n_9257);
  nand g183267 (n_842, g812, n_9257);
  nand g183209 (n_841, g2051, n_9257);
  not g182191 (n_840, g347);
  nand g182344 (n_839, g4674, n_177);
  nand g183317 (n_838, n_460, n_474);
  nand g183214 (n_837, g4239, n_9257);
  nand g183272 (n_836, g4489, n_9257);
  nand g183246 (n_835, g3566, n_9257);
  not g182217 (n_834, n_1573);
  nand g182488 (n_833, g6255, n_9257);
  nand g183275 (n_832, g5583, n_9257);
  nand g183271 (n_831, new_g7097_, n_9257);
  nand g182710 (n_830, g2994, n_9257);
  nand g182553 (n_829, g3594, n_9257);
  nand g183321 (n_828, g35, n_6582);
  nand g183213 (n_827, g20763, n_9257);
  nand g183129 (n_826, g1874, n_9257);
  nand g183196 (n_825, g2799, n_9257);
  nand g182669 (n_824, g2610, n_9257);
  nand g182869 (n_823, new_g10409_, n_822);
  nand g183326 (n_821, g35, n_155);
  not g182224 (n_820, g4681);
  nand g183245 (n_819, g1111, n_9257);
  nand g182498 (n_818, g3203, n_9257);
  nor g183376 (n_817, n_9257, n_816);
  nand g182495 (n_815, g3255, n_9257);
  nand g182456 (n_814, g3401, n_9257);
  not g182932 (n_813, n_433);
  not g182900 (n_812, n_314);
  not g182903 (n_811, n_265);
  not g182905 (n_810, n_397);
  not g182909 (n_809, n_355);
  not g182912 (n_808, n_257);
  not g182916 (n_807, n_419);
  not g182922 (n_806, n_264);
  not g182925 (n_805, n_804);
  not g182935 (n_803, n_802);
  not g182951 (n_801, n_1425);
  not g182959 (n_800, n_1422);
  nand g183066 (n_799, g5929, n_9257);
  nand g183254 (n_798, g5216, n_9257);
  nand g183279 (n_797, g3813, n_9257);
  nand g183110 (n_796, g225, n_9257);
  nand g182588 (n_795, g4462, n_9257);
  nand g183212 (n_794, g3506, n_9257);
  nand g183011 (n_793, g3857, n_9257);
  nand g183013 (n_792, g3466, n_9257);
  nand g183015 (n_791, g2177, n_9257);
  nand g183016 (n_790, g6653, n_9257);
  nand g183017 (n_789, g2819, n_9257);
  nand g183019 (n_788, g776, n_9257);
  nand g183020 (n_787, g2523, n_9257);
  nand g183021 (n_786, g1554, n_9257);
  nand g183023 (n_785, g4076, n_9257);
  nand g183025 (n_784, g5591, n_9257);
  nand g183027 (n_783, g5559, n_9257);
  nand g183028 (n_782, g2775, n_9257);
  nand g183029 (n_781, g3831, n_9257);
  nand g183033 (n_780, g6637, n_9257);
  nand g183035 (n_779, g6163, n_9257);
  nand g183036 (n_778, g2533, n_9257);
  nand g183037 (n_777, g3949, n_9257);
  nand g183039 (n_776, g146, n_9257);
  nand g183040 (n_775, g1171, n_9257);
  nand g183041 (n_774, g482, n_9257);
  nand g183043 (n_773, g5052, n_9257);
  nand g183044 (n_772, g3602, n_9257);
  nand g183045 (n_771, g5901, n_9257);
  nand g183047 (n_770, g1221, n_9257);
  nand g183049 (n_769, g3921, n_9257);
  nand g183051 (n_768, g5817, n_9257);
  nand g183052 (n_767, g2619, n_9257);
  nand g183053 (n_766, g3933, n_9257);
  nand g182538 (n_765, g3542, n_9257);
  nand g183055 (n_764, g1484, n_9257);
  nand g183057 (n_763, g1099, n_9257);
  nand g183059 (n_762, g2868, n_9257);
  nand g183060 (n_761, g5272, n_9257);
  nand g183061 (n_760, g1768, n_9257);
  nand g183063 (n_759, g5029, n_9257);
  nand g183064 (n_758, g150, n_9257);
  nand g183065 (n_757, g2575, n_9257);
  nand g182432 (n_756, g2922, n_9257);
  nand g183067 (n_755, g5224, n_9257);
  nand g183069 (n_754, g6279, n_9257);
  nand g183098 (n_753, g1041, n_9257);
  nand g183071 (n_752, g4112, n_9257);
  nand g183073 (n_751, g3490, n_9257);
  nand g183075 (n_750, g4176, n_9257);
  nand g183076 (n_749, g4122, n_9257);
  nand g183077 (n_748, g3909, n_9257);
  nand g183081 (n_747, g6605, n_9257);
  not g182919 (n_746, n_745);
  nand g183083 (n_744, g763, n_9257);
  nand g183084 (n_743, g1890, n_9257);
  nand g183085 (n_742, g5260, n_9257);
  nand g183087 (n_741, g6565, n_9257);
  nand g183089 (n_740, g6283, n_9257);
  nand g183091 (n_739, g6621, n_9257);
  nand g183093 (n_738, g2016, n_9257);
  nand g182735 (n_737, g1183, n_9257);
  nand g183095 (n_736, g2153, n_9257);
  nand g183097 (n_735, g1926, n_9257);
  nand g183099 (n_734, g4146, n_9257);
  nand g183100 (n_733, g5208, n_9257);
  nand g183101 (n_732, g4966, n_9257);
  nand g182663 (n_731, g4584, n_9257);
  nand g183103 (n_730, g1882, n_9257);
  nand g183107 (n_729, g1608, n_9257);
  nand g183109 (n_728, g6523, n_9257);
  nand g183111 (n_727, g1710, n_9257);
  nand g183295 (n_726, g35, n_6359);
  nand g183113 (n_725, g5863, n_9257);
  nand g183115 (n_724, g1526, n_9257);
  nand g183117 (n_723, g5164, n_9257);
  nand g183072 (n_722, g2461, n_9257);
  nand g183120 (n_721, g1779, n_9257);
  nand g183122 (n_720, g1740, n_9257);
  nand g183124 (n_719, g2089, n_9257);
  nand g183126 (n_718, g1964, n_9257);
  nand g183130 (n_717, new_g6875_, n_9257);
  nand g183131 (n_716, g2984, n_9257);
  nand g183132 (n_715, g4793, n_9257);
  nand g183134 (n_714, g4659, n_9257);
  nand g183136 (n_713, g6649, n_9257);
  nand g183138 (n_712, g5517, n_9257);
  nand g183140 (n_711, g1008, n_9257);
  nand g183142 (n_710, g6307, n_9257);
  nand g182730 (n_709, g2547, n_9257);
  nand g183146 (n_708, g5220, n_9257);
  nand g183148 (n_707, g1193, n_9257);
  nand g183150 (n_706, g3570, n_9257);
  nand g183261 (n_705, g2625, n_9257);
  nand g183154 (n_704, g2008, n_9257);
  nand g183155 (n_703, g1821, n_9257);
  nand g183156 (n_702, g1030, n_9257);
  nand g183180 (n_701, g1467, n_9257);
  nand g183158 (n_700, g4601, n_9257);
  nand g183160 (n_699, g758, n_9257);
  nand g183162 (n_698, g1870, n_9257);
  nand g183163 (n_697, g5200, n_9257);
  nand g183164 (n_696, g2860, n_9257);
  nand g183166 (n_695, g6044, n_9257);
  nand g183167 (n_694, g1306, n_9257);
  nand g183168 (n_693, g2970, n_9257);
  nand g183170 (n_692, g2315, n_9257);
  nand g183171 (n_691, g2279, n_9257);
  nand g183172 (n_690, g1917, n_9257);
  nand g182609 (n_689, g232, n_9257);
  nand g183174 (n_688, g1756, n_9257);
  nand g182635 (n_687, g2004, n_9257);
  nand g183178 (n_686, g1514, n_9257);
  nand g183179 (n_685, g1564, n_9257);
  nand g182659 (n_684, g5555, n_9257);
  nand g183182 (n_683, g2287, n_9257);
  nand g183184 (n_682, g2567, n_9257);
  nand g183186 (n_681, g2098, n_9257);
  nand g183187 (n_680, g1345, n_9257);
  nand g183188 (n_679, g2491, n_9257);
  nand g183190 (n_678, g2255, n_9257);
  nand g182515 (n_677, g1752, n_580);
  nand g183192 (n_676, g4300, n_9257);
  nand g183194 (n_675, g6263, n_9257);
  nand g183281 (n_674, g6295, n_9257);
  nand g183198 (n_673, g2433, n_9257);
  nand g183200 (n_672, g1616, n_9257);
  nand g183202 (n_671, g6098, n_9257);
  nand g183205 (n_670, g5571, n_9257);
  nand g183206 (n_669, g1664, n_9257);
  nand g183210 (n_668, g6303, n_9257);
  nand g183215 (n_667, g790, n_9257);
  nand g183216 (n_666, g2898, n_9257);
  nand g183218 (n_665, g753, n_9257);
  nand g183121 (n_664, g4411, n_9257);
  nand g183226 (n_663, new_g12440_, n_9257);
  nand g183227 (n_662, g1024, n_9257);
  nand g183228 (n_661, g405, n_9257);
  nand g183230 (n_660, g3195, n_9257);
  nand g183234 (n_659, g5611, n_9257);
  nand g183236 (n_658, g1978, n_9257);
  nand g183239 (n_657, g1129, n_9257);
  nand g183240 (n_656, g3247, n_9257);
  nand g183242 (n_655, g6629, n_9257);
  nand g183244 (n_654, g157, n_9257);
  nand g182559 (n_653, g749, n_9257);
  nand g183283 (n_652, g1728, n_9257);
  nand g183250 (n_651, g4049, n_9257);
  nand g183252 (n_650, g2852, n_9257);
  nand g183258 (n_649, g401, n_9257);
  nand g183262 (n_648, g3698, n_9257);
  nand g183265 (n_647, g2807, n_9257);
  nand g183268 (n_646, g2161, n_9257);
  nand g183270 (n_645, g1478, n_9257);
  nand g183274 (n_644, g1620, n_9257);
  nand g182653 (n_643, g3897, n_9257);
  nand g183276 (n_642, g5212, n_9257);
  nand g183278 (n_641, g1002, n_9257);
  nand g183280 (n_640, g4983, n_9257);
  nand g182563 (n_639, g6299, n_9257);
  nand g182584 (n_638, g2936, n_9257);
  nand g183282 (n_637, g2307, n_9257);
  nand g183284 (n_636, g1442, n_9257);
  nand g183286 (n_635, g1959, n_9257);
  nand g182651 (n_634, g2886, n_9257);
  nand g183290 (n_633, g3953, n_9257);
  nand g183293 (n_632, n_9257, n_631);
  nand g183088 (n_630, g5057, n_9257);
  nand g183298 (n_629, g35, n_169);
  nand g183299 (n_628, n_9257, n_2870);
  nand g183300 (n_627, n_9257, n_626);
  nand g183301 (n_625, g35, n_624);
  nand g183304 (n_623, g35, n_24);
  nand g183305 (n_622, n_9257, n_102);
  nor g182728 (n_621, g35, n_620);
  nand g183310 (n_619, g35, n_6580);
  nand g183313 (n_618, n_617, n_968);
  nand g182652 (n_616, g5062, n_9257);
  nand g183314 (n_615, g6645, n_9257);
  nand g183320 (n_614, g35, n_108);
  nand g183014 (n_613, g767, n_9257);
  nand g183327 (n_612, n_1040, n_1891);
  nand g183329 (n_611, g35, n_80);
  nand g183330 (n_610, n_9257, n_238);
  nand g183336 (n_609, g35, n_4492);
  nand g182647 (n_608, g3530, n_9257);
  nand g183339 (n_607, n_467, n_477);
  not g182251 (n_606, g23683);
  nand g183157 (n_605, g239, n_9257);
  nand g182734 (n_604, g538, n_9257);
  nand g182649 (n_603, g5831, n_9257);
  nand g182484 (n_602, g5046, n_601);
  nand g183389 (n_600, n_599, n_476);
  nand g183251 (n_598, g5953, n_9257);
  nor g183315 (n_597, g4258, n_9257);
  nand g182504 (n_596, g5062, n_491);
  nand g183430 (n_595, n_5340, n_1445);
  nand g183432 (n_594, n_468, n_466);
  nand g182340 (n_593, g8786, n_592);
  nand g183479 (n_591, n_465, n_471);
  nand g183296 (n_590, n_9257, n_182);
  not g182939 (n_589, n_334);
  nand g183285 (n_588, g5188, n_9257);
  nand g182502 (n_587, g424, n_9257);
  nand g182739 (n_586, g1696, n_9257);
  nand g183247 (n_585, g4492, n_9257);
  nand g182682 (n_584, g358, n_9257);
  nand g183434 (n_583, n_455, n_582);
  nand g182510 (n_581, g1744, n_580);
  nand g182500 (n_579, g5547, n_9257);
  nand g182461 (n_578, g2811, n_9257);
  nand g182447 (n_577, g2040, n_982);
  nand g182686 (n_574, g5204, n_9257);
  nand g183243 (n_573, g2295, n_9257);
  nand g182285 (n_572, g2181, n_9257);
  nand g182613 (n_571, g1018, n_9257);
  nand g183235 (n_570, g1783, n_9257);
  nand g183248 (n_569, g5041, n_9257);
  nor g182614 (n_568, g35, n_968);
  nand g182499 (n_567, g6159, n_9257);
  nand g183219 (n_566, g5244, n_9257);
  nor g182496 (n_565, g2331, n_1011);
  nand g182493 (n_564, g3187, n_9257);
  nand g182547 (n_561, g5575, n_9257);
  nand g182636 (n_560, g2595, n_9257);
  nand g182702 (n_559, g3243, n_9257);
  not g182908 (n_558, n_352);
  nand g183080 (n_557, g2122, n_9257);
  nand g182284 (n_556, g2265, n_9257);
  nand g182642 (n_555, g6444, n_9257);
  nand g182492 (n_554, g6035, n_9257);
  nand g182645 (n_553, g5232, n_9257);
  nand g182326 (n_552, g55, n_96);
  nand g183183 (n_551, g246, n_9257);
  nand g182520 (n_550, g1373, n_9257);
  nand g183165 (n_549, g2787, n_9257);
  nand g182724 (n_548, g5196, n_9257);
  nand g182540 (n_547, g1736, n_9257);
  nand g182634 (n_545, g3610, n_9257);
  nand g182472 (n_544, g5873, n_9257);
  nand g183220 (n_543, g3863, n_9257);
  nand g182508 (n_542, g417, n_9257);
  nand g183009 (n_541, g6227, n_9257);
  nand g182537 (n_540, g2681, n_9257);
  nand g182320 (n_539, n_36, n_483);
  nand g182585 (n_538, g20899, n_9257);
  nand g182481 (n_537, g3215, n_9257);
  nand g182478 (n_536, g3873, n_9257);
  nor g182566 (n_535, g35, n_534);
  nand g182534 (n_533, g4253, n_9257);
  nand g182632 (n_532, g6187, n_9257);
  nand g182631 (n_531, g1361, n_9257);
  nand g182548 (n_530, g1036, n_9257);
  nand g182316 (n_529, g3598, n_9257);
  nand g182619 (n_528, g5352, n_9257);
  nand g182307 (n_527, g817, n_9257);
  nand g182475 (n_526, g3223, n_9257);
  nand g183462 (n_525, n_209, n_524);
  nand g182523 (n_523, g370, n_9257);
  nand g182306 (n_522, g2571, n_9257);
  nand g182290 (n_521, g3689, n_9257);
  nand g182289 (n_520, g3586, n_9257);
  nand g183224 (n_519, g294, n_9257);
  nand g182303 (n_518, g6589, n_9257);
  nand g182628 (n_517, g739, n_9257);
  nand g182615 (n_516, g5236, n_9257);
  nand g183291 (n_515, g2112, n_9257);
  nand g183145 (n_514, g6287, n_9257);
  nand g183287 (n_513, g4486, n_9257);
  nand g183306 (n_512, n_147, n_511);
  nand g183221 (n_510, g785, n_9257);
  not g182915 (n_509, n_317);
  nand g183289 (n_508, g2217, n_9257);
  nand g183223 (n_507, g1996, n_9257);
  nand g183288 (n_506, g2583, n_9257);
  wire w275, w276, w277, w278;
  nand g182071 (n_505, w276, w278);
  nand g317 (w278, w277, g262);
  not g315 (w277, g239);
  nand g314 (w276, w275, g239);
  not g313 (w275, g262);
  nand g182299 (n_504, g2767, n_9257);
  nand g183034 (n_503, g3881, n_9257);
  nand g183139 (n_502, g3139, n_9257);
  nand g182377 (n_501, g1221, n_4);
  nand g182471 (n_500, g550, n_9257);
  nand g183135 (n_499, g1604, n_9257);
  nand g182625 (n_498, g5949, n_9257);
  nand g183222 (n_497, g2514, n_9257);
  nand g182621 (n_496, g5148, n_9257);
  nand g182463 (n_495, g1802, n_9257);
  nand g182623 (n_494, g3239, n_9257);
  nand g182624 (n_493, g21176, n_9257);
  nor g183391 (n_492, n_491, n_1891);
  nand g182622 (n_490, g255, n_9257);
  nand g182300 (n_489, g1657, n_9257);
  nand g183507 (n_1452, n_461, n_488);
  not g182953 (n_3320, n_487);
  wire w279, w280, w281, w282;
  nand g182080 (n_1562, w280, w282);
  nand g322 (w282, w281, g12422);
  not g321 (w281, g6381);
  nand g320 (w280, w279, g6381);
  not g318 (w279, g12422);
  nand g183524 (n_1705, n_816, n_464);
  wire w283, w284, w285, w286;
  nand g182083 (n_1443, w284, w286);
  nand g327 (w286, w285, g6727);
  not g326 (w285, g12470);
  nand g325 (w284, w283, g12470);
  not g323 (w283, g6727);
  nand g183575 (n_1436, n_485, n_486);
  wire w287, w288, w289, w290;
  nand g182085 (n_1430, w288, w290);
  nand g332 (w290, w289, g25219);
  not g331 (w289, g12238);
  nand g330 (w288, w287, g12238);
  not g328 (w287, g25219);
  wire w291, w292, w293, w294;
  nand g182086 (n_1553, w292, w294);
  nand g338 (w294, w293, g3338);
  not g337 (w293, g11349);
  nand g335 (w292, w291, g11349);
  not g334 (w291, g3338);
  nand g183529 (n_1456, g35, n_6562);
  nand g182778 (n_1432, g691, n_195);
  nor g183532 (n_3969, g1199, n_9257);
  nand g183612 (n_1547, n_469, n_901);
  nand g182742 (n_1489, g1772, n_488);
  nand g182744 (n_1487, g2197, n_484);
  nand g182745 (n_1875, g5016, n_1916);
  wire w295, w296, w297, w298;
  nand g182082 (n_1446, w296, w298);
  nand g343 (w298, w297, g6035);
  not g342 (w297, g12350);
  nand g340 (w296, w295, g12350);
  not g339 (w295, g6035);
  nor g182747 (n_1926, g4322, n_1805);
  nor g182754 (n_1886, g376, n_957);
  nand g183572 (n_1437, g35, n_191);
  fflopd g34_reg(.CK (clock), .D (n_483), .Q (g55));
  nand g183567 (n_1555, g35, n_183);
  nand g183544 (n_1460, n_457, n_484);
  nor g183543 (n_2331, g1306, n_9257);
  nand g183539 (n_1616, g35, n_6361);
  nand g183535 (n_1458, g35, n_54);
  nor g183533 (n_3903, g1542, n_9257);
  nand g183528 (n_1454, g35, n_6560);
  nand g182875 (n_1411, new_g7004_, n_106);
  nand g183540 (n_1605, n_456, n_911);
  nand g182750 (n_1728, g1906, n_1317);
  nor g183513 (n_1893, n_9257, n_2638);
  not g182977 (n_1889, n_1610);
  nand g182876 (n_1410, new_g7051_, n_462);
  nand g182874 (n_1540, new_g7028_, n_458);
  nand g182866 (n_1409, new_g10371_, n_482);
  nand g182864 (n_1414, g6209, n_0);
  nand g182860 (n_1412, g3161, n_70);
  nand g182858 (n_1543, new_g7074_, n_109);
  nand g182853 (n_1415, g3863, n_43);
  nand g182849 (n_1542, g5517, n_231);
  nand g182846 (n_1541, g5863, n_50);
  nand g183595 (n_1423, n_481, n_482);
  nand g182845 (n_1544, g3512, n_3);
  nand g182834 (n_1416, g6555, n_77);
  nand g182833 (n_1546, g5170, n_10);
  nand g182831 (n_1424, g2051, n_480);
  nand g182830 (n_1426, g1648, n_2109);
  not g182229 (n_4424, g1585);
  nand g182768 (n_1560, g1171, n_479);
  nand g182785 (n_1431, n_150, n_2638);
  nand g182801 (n_1427, g2331, n_208);
  nand g182799 (n_1428, g1636, n_582);
  nand g182792 (n_1557, g2040, n_46);
  nand g182791 (n_1429, n_38, n_2640);
  nand g182877 (n_3614, new_g10405_, n_478);
  nand g182837 (n_1711, g3506, n_137);
  nand g182764 (n_2811, g6227, n_477);
  nand g182772 (n_2766, g3881, n_476);
  nand g182872 (n_2996, new_g7097_, n_475);
  nand g182775 (n_2957, g5535, n_474);
  nand g183551 (n_1853, g35, n_484);
  nand g182756 (n_2506, g4899, n_913);
  nor g183574 (n_1918, n_9257, n_473);
  nand g182755 (n_1892, g4709, n_486);
  nand g183570 (n_1780, g35, n_488);
  nor g182776 (n_1950, g1526, n_472);
  nand g182758 (n_2733, g5188, n_471);
  nand g182759 (n_1722, g5873, n_470);
  nand g183580 (n_1738, g35, n_911);
  nand g182873 (n_4831, new_g6875_, n_469);
  nand g183557 (n_2423, n_90, n_5340);
  nand g182840 (n_1727, g6203, n_91);
  nand g182838 (n_1723, g5857, n_14);
  nand g182836 (n_1708, g3155, n_18);
  nand g182868 (n_4444, new_g10375_, n_908);
  nand g182766 (n_1715, g6565, n_468);
  nand g183560 (n_8116, g35, n_1026);
  nand g182760 (n_1710, g6219, n_467);
  nand g182763 (n_2738, g6573, n_466);
  nand g182827 (n_1850, g1526, n_472);
  nand g182777 (n_1720, g5180, n_465);
  nand g182779 (n_2796, g3179, n_464);
  nand g182816 (n_8546, g2476, n_463);
  nand g183614 (n_2296, n_462, n_478);
  nand g182780 (n_1706, g3522, n_617);
  nand g182783 (n_1803, g1772, n_461);
  not g183004 (n_1945, n_4842);
  nor g182789 (n_2719, g4709, n_486);
  nor g182803 (n_2721, g4899, n_913);
  nand g182767 (n_1721, g5527, n_460);
  nand g183610 (n_2294, n_458, n_459);
  nand g182797 (n_1763, g2197, n_457);
  nand g182795 (n_1867, g2465, n_456);
  nor g182794 (g25259, g1636, n_455);
  not g182976 (n_1972, n_454);
  nand g182878 (n_3616, new_g10401_, n_459);
  nor g182808 (n_8579, g1760, n_580);
  nand g182809 (n_8550, g1648, n_453);
  nand g182811 (n_8548, g2342, n_452);
  nand g182814 (n_8551, g2208, n_451);
  nor g182815 (n_8577, g2587, n_978);
  nand g182824 (n_3378, g1442, n_42);
  nand g182826 (n_7970, g1099, n_86);
  nand g183602 (n_2359, g35, n_1438);
  nand g182870 (n_5462, new_g10413_, n_904);
  nand g183600 (n_2626, g35, n_1441);
  nand g183597 (n_2623, g35, n_1550);
  nand g183594 (n_2457, g35, n_1442);
  nand g182828 (n_2544, g1183, n_450);
  nand g183598 (n_2497, g35, n_1549);
  nand g182881 (n_6159, new_g6905_, n_481);
  nor g183593 (n_1958, g7916, n_9257);
  nor g183590 (n_1980, g7946, n_9257);
  nand g183603 (n_2597, g35, n_1440);
  not g183001 (n_5195, n_449);
  not g182988 (n_5148, n_448);
  not g183005 (n_5044, n_447);
  not g182998 (n_5216, n_446);
  nand g182854 (n_5346, g667, n_237);
  not g183008 (g25114, n_445);
  nor g183348 (n_444, g5863, g5857);
  nand g183443 (n_443, g35, g4157);
  nand g183346 (n_442, g2476, g2449);
  nand g183450 (n_441, g35, g546);
  nor g182365 (n_440, g2547, g2541);
  nand g183452 (n_439, g35, g2491);
  nand g183351 (n_438, g35, g2917);
  nand g183371 (n_437, g2279, g2273);
  nand g183516 (n_436, g35, g4264);
  nor g182388 (n_435, g2413, g2407);
  nand g183403 (n_434, g2319, g2311);
  nand g183509 (n_433, g35, g9019);
  nand g183405 (n_432, g35, g1644);
  nand g183352 (n_431, g5011, g4836);
  nand g183360 (n_430, g35, g21292);
  nand g183506 (n_429, g35, g4653);
  nand g183332 (n_428, g35, g2882);
  nand g183345 (n_427, g370, g8719);
  nand g183342 (n_426, g35, g3689);
  nand g183350 (n_425, g723, g817);
  nor g182400 (n_424, g1489, g1442);
  nand g183341 (n_423, g35, g4411);
  nand g183333 (n_422, g2265, g2259);
  nor g183344 (n_421, g3161, g3155);
  nand g183427 (n_420, g35, g1779);
  nand g183483 (n_419, g12470, g6585);
  nand g183431 (n_418, g35, g4172);
  nand g183404 (n_417, g35, g2860);
  nor g183311 (n_416, new_g10383_, g4608);
  nor g182401 (n_415, g1974, g1968);
  nand g183436 (n_414, g35, g4176);
  nor g182392 (n_413, g1840, g1834);
  nand g183592 (n_412, g1514, g1526);
  nand g183377 (n_411, g1624, g1604);
  nor g182363 (n_410, g490, new_g8038_);
  nand g183484 (n_409, g35, g2047);
  nor g182366 (n_408, g5148, g5142);
  nor g182373 (n_407, g3139, g3133);
  nor g182403 (n_406, g1854, g1848);
  nand g183429 (n_405, g5148, g5142);
  nor g183316 (n_404, g5170, g5164);
  nand g183387 (n_403, g6187, g6181);
  nand g183501 (n_402, g35, g1548);
  nor g182405 (n_401, g3490, g3484);
  nor g182385 (n_400, g1706, g1700);
  nand g183481 (n_399, g35, g1913);
  nand g183522 (n_398, g35, g862);
  nand g183390 (n_397, g1894, g1874);
  nand g183470 (n_396, g35, g2868);
  nand g183469 (n_395, g35, g5092);
  nand g183466 (n_394, g2941, g2936);
  nand g183459 (n_393, g35, g2960);
  nand g183438 (n_392, g35, g1772);
  nand g183475 (n_391, g35, g2852);
  nand g183456 (n_390, g35, g5689);
  nand g183395 (n_389, g4157, g4146);
  nor g182370 (n_388, g2681, g2675);
  nand g183457 (n_387, g35, g2844);
  nor g182333 (n_386, g538, g209);
  nand g183455 (n_385, g35, g2894);
  nand g183451 (n_384, g35, g1484);
  nor g182398 (n_383, g2265, g2259);
  nand g183448 (n_382, g2975, g2970);
  nand g183446 (n_381, g2208, g2181);
  nand g183356 (n_380, g35, g37);
  nor g182395 (n_379, g6187, g6181);
  nand g183447 (n_378, g35, g4443);
  nand g183324 (n_377, g35, g2994);
  nand g183449 (n_376, g35, g2066);
  nand g183440 (n_375, g1706, g1700);
  nand g183435 (n_374, g2533, g2527);
  nor g182382 (n_373, g3841, g3835);
  nand g183428 (n_372, g35, g6035);
  nand g183425 (n_371, g35, g2922);
  nor g182394 (n_370, g5841, g5835);
  nor g182391 (n_369, g2122, g2116);
  nor g182332 (n_368, g4093, g4076);
  nor g182347 (n_367, g4297, g10122);
  nor g182351 (n_366, g2223, g2204);
  nor g182346 (n_365, g11447, g8783);
  nand g183323 (n_364, g753, g655);
  nor g182381 (n_363, g1559, g1548);
  nor g182384 (n_362, g1720, g1714);
  nor g182402 (n_361, g2279, g2273);
  nor g182541 (n_360, g979, g1052);
  nor g182542 (n_359, g1322, g1395);
  nor g182350 (n_358, g4405, g7243);
  nand g183419 (n_357, g1024, g1002);
  nand g183415 (n_356, g2028, g2020);
  nand g183408 (n_355, g11418, g3893);
  nand g183410 (n_354, g35, g2848);
  nor g182364 (n_353, g6533, g6527);
  nand g183407 (n_352, g6745, g35);
  nand g183325 (n_351, g1720, g1714);
  nand g183328 (n_350, g35, g2338);
  nand g183340 (n_349, g35, g2606);
  nor g182343 (n_348, g4864, g4836);
  nand g183357 (n_347, g35, g4249);
  nand g183363 (n_346, g6744, g35);
  nand g183365 (n_345, g2955, g2950);
  nand g183368 (n_344, g35, g6381);
  nand g183374 (n_343, g1379, g1345);
  nand g183378 (n_342, g35, g2950);
  nand g183384 (n_341, g35, g2936);
  nand g183386 (n_340, g35, g2873);
  nand g183393 (n_339, g401, g405);
  nand g183396 (n_338, g35, g1932);
  nand g183406 (n_337, g35, g2856);
  nand g183504 (n_1324, g35, g5817);
  nand g183495 (n_804, g35, g25219);
  nand g183518 (n_2217, g35, g12923);
  nor g183537 (n_4291, g1171, g1183);
  nand g183625 (n_445, new_g7004_, g5297);
  nand g183564 (n_909, g35, g1008);
  nand g183492 (n_1166, g1221, g1205);
  nand g183508 (n_1506, g35, g5180);
  nand g183488 (n_745, g35, g5535);
  nand g183514 (n_1773, g6750, g35);
  nand g183521 (n_575, g35, g1129);
  fflopd g4281_reg(.CK (clock), .D (g8839), .Q (g4281));
  fflopd g4297_reg(.CK (clock), .D (g10122), .Q (g4297));
  nand g183616 (n_892, new_g7028_, new_g10401_);
  nand g183589 (n_454, g35, g7916);
  nand g183618 (n_449, g6555, g6549);
  fflopd g191_reg(.CK (clock), .D (g8358), .Q (g191));
  fflopd g4291_reg(.CK (clock), .D (g9019), .Q (g4291));
  nand g183620 (n_895, g3512, g3506);
  nand g183606 (n_893, g3863, g3857);
  nand g183605 (n_897, g3161, g3155);
  nand g183494 (n_1378, g35, g6573);
  nand g183497 (n_1158, g35, g3881);
  nand g183517 (n_1500, g35, g5527);
  nand g183502 (n_1155, g1564, g1548);
  nand g183578 (n_910, g35, g3530);
  nand g183617 (n_899, new_g6905_, new_g10371_);
  nand g183519 (n_802, g4601, g4593);
  fflopd g4452_reg(.CK (clock), .D (g7245), .Q (g4452));
  nor g183536 (n_1561, g1514, g1526);
  nand g183520 (n_880, g35, g5188);
  fflopd g4411_reg(.CK (clock), .D (g7257), .Q (g4411));
  nor g183577 (n_6016, g2070, g1996);
  fflopd g1333_reg(.CK (clock), .D (g8475), .Q (g1333));
  fflopd g4180_reg(.CK (clock), .D (g8789), .Q (g4180));
  nor g182806 (n_1573, g4141, g4082);
  nand g183582 (n_1421, g3179, g3171);
  fflopd g4188_reg(.CK (clock), .D (g11447), .Q (g8783));
  nand g183555 (n_1417, g5881, g5873);
  nor g183559 (n_5383, g2629, g2555);
  nand g183584 (n_1420, g5535, g5527);
  fflopd g2715_reg(.CK (clock), .D (g35), .Q (new_g7717_));
  nand g183554 (n_1418, g3530, g3522);
  nand g183581 (n_1596, g4849, g4843);
  nand g183579 (n_1577, g35, g3522);
  nand g183568 (n_1694, g35, g4388);
  nand g183591 (n_1610, g385, g376);
  nand g183556 (n_1699, g35, g3466);
  nand g183553 (n_3736, g35, g6163);
  fflopd g4871_reg(.CK (clock), .D (g4864), .Q (g4871));
  fflopd g1079_reg(.CK (clock), .D (g17291), .Q (g17316));
  nor g182823 (n_7848, g1146, g1099);
  fflopd g4674_reg(.CK (clock), .D (g4646), .Q (g4674));
  fflopd g4681_reg(.CK (clock), .D (g4674), .Q (g4681));
  fflopd g1430_reg(.CK (clock), .D (g17423), .Q (g1430));
  fflopd g6329_reg(.CK (clock), .D (g12422), .Q (g14779));
  fflopd g5290_reg(.CK (clock), .D (g12238), .Q (g14662));
  fflopd g6675_reg(.CK (clock), .D (g12470), .Q (g14828));
  fflopd g3281_reg(.CK (clock), .D (g11349), .Q (g13895));
  fflopd g3983_reg(.CK (clock), .D (g11418), .Q (g13966));
  nor g183611 (n_6886, new_g7004_, g5297);
  fflopd g1242_reg(.CK (clock), .D (g12919), .Q (g23683));
  nand g183381 (n_336, g1854, g1848);
  nand g183412 (n_335, g5841, g5835);
  nand g183526 (n_334, g35, g9251);
  nand g183411 (n_333, g35, g2465);
  nand g183355 (n_332, g3490, g3484);
  nand g183400 (n_331, g4765, g4709);
  nand g183413 (n_330, g35, g269);
  nand g183349 (n_329, g832, g827);
  nand g183385 (n_328, g1926, g1878);
  nand g183414 (n_327, g4955, g4899);
  nor g183307 (n_326, g3512, g3506);
  nand g183354 (n_325, g35, g1798);
  nand g183442 (n_324, g896, g890);
  nand g183478 (n_323, g35, new_g6961_);
  nand g183358 (n_322, g1624, g1616);
  nand g183482 (n_321, g2342, g2315);
  nor g182393 (n_320, g1988, g1982);
  nand g183477 (n_319, g2217, g2169);
  nand g183399 (n_318, g2122, g2116);
  nand g183480 (n_317, g4358, g4349);
  nand g183454 (n_316, g35, g3171);
  nand g183418 (n_315, g1988, g1982);
  nand g183353 (n_314, g2185, g2165);
  nor g183362 (n_313, g232, g225);
  nand g183416 (n_312, g1783, g1756);
  nand g183444 (n_311, g35, g2864);
  nand g183417 (n_310, g1974, g1968);
  nand g183445 (n_309, g35, g2223);
  nand g183361 (n_308, g2453, g2433);
  nand g183359 (n_307, g2547, g2541);
  nand g183485 (n_306, g11388, g3542);
  nand g183472 (n_305, g4486, g4483);
  nand g183409 (n_304, g1894, g1886);
  nor g183312 (n_303, g6555, g6549);
  nand g183366 (n_302, g3139, g3133);
  nand g183474 (n_301, g2051, g2024);
  nor g182321 (n_300, g4674, g4646);
  nand g183421 (n_299, g1840, g1834);
  nand g183476 (n_298, g35, g2907);
  nor g182379 (n_297, g2533, g2527);
  nand g183402 (n_296, g6533, g6527);
  nand g183364 (n_295, g35, g2898);
  nand g183471 (n_294, g35, g2197);
  nand g183367 (n_293, g2185, g2177);
  nand g183388 (n_292, g12300, g5547);
  nor g182544 (n_291, g7946, g8475);
  nor g183319 (n_290, g5517, g5511);
  nand g183369 (n_289, g1917, g1890);
  nand g183335 (n_288, g35, g20652);
  nand g183473 (n_287, g5495, g5489);
  nor g183318 (n_286, g3863, g3857);
  fflopd g4474_reg(.CK (clock), .D (g4467), .Q (new_g12875_));
  nand g183322 (n_285, g2319, g2299);
  nand g183372 (n_284, g35, g21176);
  nand g183398 (n_283, g1792, g1740);
  nand g183373 (n_282, g35, g4146);
  nand g183460 (n_281, g35, g2970);
  nand g183439 (n_280, g35, g2357);
  nand g183503 (n_279, g35, g4843);
  nand g183424 (n_278, g35, g6727);
  nand g183437 (n_277, g2351, g2303);
  nand g183397 (n_276, g2060, g2012);
  nand g183441 (n_275, g2907, g2902);
  nand g183394 (n_274, g232, g225);
  nand g183392 (n_273, g35, g2975);
  nand g183347 (n_272, g35, g2625);
  nand g183422 (n_271, g5057, g5022);
  nand g183423 (n_270, g2413, g2407);
  nor g182376 (n_269, g862, g896);
  nand g183370 (n_268, g3841, g3835);
  nand g183420 (n_267, g35, g2204);
  nor g183303 (n_266, g6209, g6203);
  nand g183375 (n_265, g12350, g5893);
  nand g183491 (n_264, g35, g8839);
  nand g183426 (n_263, g2028, g2008);
  nand g183453 (n_262, g3684, g4871);
  nor g182444 (n_261, g753, g655);
  nand g183343 (n_260, g12923, g17423);
  nand g183468 (n_259, g2917, g2912);
  nand g183461 (n_258, g35, g4245);
  nand g183433 (n_257, g2453, g2445);
  nor g182390 (n_256, g5495, g5489);
  nand g183401 (n_255, g2619, g2567);
  nand g183463 (n_254, g554, g807);
  nand g183465 (n_253, g35, g4253);
  nand g183382 (n_252, g35, g2472);
  nand g183458 (n_251, g35, g2912);
  nand g183383 (n_250, g35, g2941);
  nand g183467 (n_249, g2610, g2583);
  nand g183464 (n_248, g2681, g2675);
  nand g183523 (n_247, g35, g1205);
  nand g183379 (n_246, g4467, new_g6961_);
  nand g183331 (n_245, g35, g1664);
  nand g183380 (n_244, g4646, g21245);
  nand g183525 (n_1881, g6748, g35);
  nand g183609 (n_900, new_g7074_, new_g10409_);
  fflopd g1236_reg(.CK (clock), .D (g10500), .Q (g1236));
  nand g183496 (n_1355, g35, g5124);
  nand g183615 (n_446, g5170, g5164);
  nand g183619 (n_894, g5517, g5511);
  nand g183546 (n_914, g35, g3817);
  nand g183549 (n_487, g35, g6509);
  fflopd g4405_reg(.CK (clock), .D (g7243), .Q (g4405));
  nand g183498 (n_1554, g490, g482);
  nand g183489 (n_1367, g35, g4040);
  nand g183534 (n_1530, g35, g5873);
  nor g182753 (n_1512, g19357, g1333);
  nand g183527 (n_1216, g35, g1135);
  nand g183487 (n_855, g35, g6227);
  nand g183493 (n_1584, g35, g6565);
  nor g182752 (n_849, g499, g518);
  fflopd g4308_reg(.CK (clock), .D (g9251), .Q (g4308));
  nand g183550 (n_1481, g5092, g5084);
  nand g183623 (n_898, g5863, g5857);
  nand g183622 (n_447, g6209, g6203);
  nand g183505 (n_1509, g35, g3873);
  nand g183604 (n_448, new_g7051_, new_g10405_);
  fflopd g1579_reg(.CK (clock), .D (g10527), .Q (g1579));
  nand g183499 (n_1309, g35, g5881);
  nand g183490 (n_1148, g35, g246);
  nor g183542 (n_1559, g4983, g4991);
  nand g183624 (n_896, new_g6928_, new_g10375_);
  nand g183510 (n_1297, g35, g3338);
  nand g183515 (n_2505, g35, g5471);
  nand g183531 (n_1352, g174, g182);
  nand g183585 (n_1625, g4264, g4258);
  nand g183511 (n_1698, g35, g3115);
  nand g183500 (n_1569, g35, g6219);
  nor g183541 (n_1558, g4793, g4801);
  nand g183512 (n_1692, g35, g4153);
  nand g183486 (n_1775, g6749, g35);
  fflopd g347_reg(.CK (clock), .D (g7540), .Q (g347));
  nand g183545 (n_1527, new_g10795_, g4621);
  fflopd g4197_reg(.CK (clock), .D (g8784), .Q (g8785));
  nand g183552 (n_1581, g847, g812);
  fflopd g4204_reg(.CK (clock), .D (g8786), .Q (g8787));
  fflopd g4210_reg(.CK (clock), .D (g8788), .Q (g8789));
  nor g183573 (n_5381, g2361, g2287);
  nand g183576 (n_3104, g1030, g1018);
  nand g183558 (n_3122, g1373, g1361);
  fflopd g1582_reg(.CK (clock), .D (g7946), .Q (g8475));
  fflopd g4207_reg(.CK (clock), .D (g8787), .Q (g8788));
  nand g183548 (n_1548, g6227, g6219);
  nand g183586 (n_2227, g35, g12919);
  fflopd g1239_reg(.CK (clock), .D (g7916), .Q (g8416));
  nor g182800 (n_1934, g174, g182);
  fflopd g4194_reg(.CK (clock), .D (g8783), .Q (g8784));
  nand g183547 (n_1425, g5188, g5180);
  nand g183561 (n_1845, g35, g2988);
  nand g183563 (n_2290, g4659, g4653);
  fflopd g4443_reg(.CK (clock), .D (g7260), .Q (g4443));
  nand g183607 (n_3789, new_g7097_, new_g10413_);
  nand g183562 (n_1422, g3881, g3873);
  nand g183569 (n_1419, g6573, g6565);
  nor g182807 (n_1955, g4057, g4064);
  nand g183621 (n_4842, new_g6875_, new_g10366_);
  fflopd g1422_reg(.CK (clock), .D (g17320), .Q (g17404));
  fflopd g4200_reg(.CK (clock), .D (g8785), .Q (g8786));
  fflopd g1322_reg(.CK (clock), .D (g13272), .Q (g1322));
  fflopd g4864_reg(.CK (clock), .D (g4836), .Q (g4864));
  fflopd g1585_reg(.CK (clock), .D (g12923), .Q (g1585));
  fflopd g1083_reg(.CK (clock), .D (g17316), .Q (g17400));
  nor g183596 (n_6881, new_g7074_, new_g10409_);
  fflopd g1087_reg(.CK (clock), .D (g17400), .Q (g1087));
  fflopd g1426_reg(.CK (clock), .D (g17404), .Q (g17423));
  fflopd g4878_reg(.CK (clock), .D (g4871), .Q (g4878));
  fflopd g5637_reg(.CK (clock), .D (g12300), .Q (g14694));
  fflopd g3632_reg(.CK (clock), .D (g11388), .Q (g13926));
  fflopd g5983_reg(.CK (clock), .D (g12350), .Q (g14738));
  fflopd g1459_reg(.CK (clock), .D (g19357), .Q (g13272));
  fflopd g358_reg(.CK (clock), .D (g8719), .Q (g358));
  not g183914 (n_242, g4273);
  not g183655 (n_241, g2327);
  not g183688 (n_239, g676);
  not g183860 (n_238, g2882);
  not g183890 (n_237, g686);
  not g183714 (n_235, g1955);
  not g183925 (n_234, g3462);
  not g183893 (n_233, g2595);
  not g183667 (n_232, g1532);
  not g184006 (n_231, g5511);
  not g183978 (n_230, g671);
  not g183875 (n_229, g2403);
  not g183664 (n_227, g1844);
  not g183767 (n_226, new_g6961_);
  not g183810 (n_225, g5046);
  not g183900 (n_224, g8787);
  not g183850 (n_223, g550);
  not g183737 (n_222, g1404);
  not g183682 (n_221, g2643);
  not g183731 (n_220, g2807);
  not g183834 (n_219, g1772);
  not g183884 (n_218, g645);
  not g183923 (n_216, g1094);
  not g183724 (n_215, g1548);
  not g183642 (n_214, g4961);
  not g183765 (n_213, g2675);
  not g183752 (n_212, g5170);
  not g183999 (n_211, g2587);
  not g183730 (n_210, g446);
  not g183940 (n_209, g8719);
  not g183749 (n_208, g2287);
  not g183669 (n_207, g2823);
  not g183653 (n_206, g4704);
  not g183675 (n_205, g324);
  not g183815 (n_203, g2051);
  not g183924 (n_200, g2648);
  not g183912 (n_199, g1111);
  not g183942 (n_198, g2236);
  not g183995 (n_197, g482);
  not g183705 (n_196, g2514);
  not g183920 (n_195, g209);
  not g183943 (n_194, g2815);
  not g183657 (n_193, g2795);
  not g183698 (n_192, g1687);
  not g183658 (n_191, g4462);
  not g183704 (n_190, g4653);
  not g183648 (n_189, g2671);
  not g184023 (n_188, g1917);
  not g184054 (n_187, g7916);
  not g183666 (n_183, g4467);
  not g183629 (n_182, g4082);
  not g183684 (n_181, g4849);
  not g183913 (n_179, g2089);
  not g183680 (n_178, g5120);
  not g183630 (n_177, g4821);
  not g183674 (n_176, g2472);
  not g183673 (n_175, g7257);
  not g183980 (n_174, g1442);
  not g183904 (n_173, g1932);
  not g183683 (n_172, g3813);
  not g183809 (n_171, g2208);
  not g183772 (n_170, g827);
  not g183865 (n_169, g4239);
  not g183722 (n_167, g896);
  not g183766 (n_166, g2775);
  not g183702 (n_165, g2084);
  not g183907 (n_164, g6505);
  not g183903 (n_163, g2606);
  not g183662 (n_162, g2338);
  not g183641 (n_161, g4749);
  not g183696 (n_159, g6159);
  not g183769 (n_156, g2803);
  not g183802 (n_155, g12923);
  not g183899 (n_152, g2779);
  not g183972 (n_151, g5821);
  not g183679 (n_150, g1312);
  not g183646 (n_148, g4760);
  not g183956 (n_147, g4349);
  not g183868 (n_146, g3333);
  not g183872 (n_145, g4939);
  not g183672 (n_144, g4443);
  not g183713 (n_143, g4659);
  not g183962 (n_142, g2787);
  not g183676 (n_141, g5813);
  not g183974 (n_139, g4258);
  not g183745 (n_137, g3512);
  not g184021 (n_136, g4793);
  not g183869 (n_135, g4382);
  not g183761 (n_134, g2555);
  not g183934 (n_132, g2116);
  not g183879 (n_130, g1189);
  not g183895 (n_129, g4894);
  not g183861 (n_128, g4754);
  not g183921 (n_127, g5467);
  not g183896 (n_126, g2193);
  not g183781 (n_123, g376);
  not g183663 (n_122, g1632);
  not g183883 (n_120, g1384);
  not g183803 (n_117, g2342);
  not g183797 (n_471, g5180);
  not g184009 (n_1047, g2093);
  not g183735 (n_1434, g996);
  not g183748 (n_2726, g3119);
  not g183792 (n_902, new_g7004_);
  not g183738 (n_1825, g1345);
  not g184036 (n_1909, g392);
  not g183706 (n_2086, g6736);
  not g183743 (n_3308, new_g10383_);
  not g183941 (n_491, g5029);
  not g183916 (n_1043, g723);
  not g183708 (n_2800, g4859);
  not g183768 (g23612, g21292);
  not g183762 (n_1618, g1367);
  not g183947 (n_462, new_g10405_);
  not g184022 (n_1009, g1648);
  not g183687 (n_1099, g4375);
  not g183747 (n_1347, g513);
  not g183919 (n_4138, g336);
  not g183986 (n_2750, g5475);
  not g183677 (n_2079, g3347);
  not g183989 (n_1050, g17400);
  not g183991 (n_1019, g17423);
  not g183758 (n_2455, g1211);
  not g183932 (n_1083, g2652);
  not g183817 (n_998, g4983);
  not g183793 (n_858, g847);
  not g183757 (n_7263, g2661);
  not g183939 (n_3256, g956);
  not g183661 (n_483, g55);
  not g183697 (n_2103, g4049);
  not g183964 (n_2753, g5037);
  not g184062 (n_473, g7946);
  not g184031 (n_468, g6573);
  not g183703 (n_2073, g6044);
  not g183981 (n_907, new_g10375_);
  not g183958 (n_624, g4628);
  not g184017 (n_599, g3881);
  not g183795 (n_5368, g1129);
  not g183994 (n_485, g4709);
  not g183685 (n_4592, g17291);
  not g184010 (n_1030, g1936);
  not g183711 (n_2081, g5352);
  not g183707 (g23002, g37);
  not g184001 (n_2210, g255);
  not g184019 (n_470, g5881);
  not g183979 (n_2816, g3470);
  not g184018 (n_2534, g2485);
  not g183759 (n_457, g2153);
  not g183888 (n_631, g2955);
  not g183977 (n_456, g2421);
  not g183806 (n_903, g1894);
  not g183719 (n_1059, g424);
  not g183835 (n_1260, g4966);
  not g183779 (n_455, g1668);
  not g183811 (n_476, g3873);
  not g183785 (n_1608, g239);
  not g183725 (n_3237, g1002);
  not g183742 (n_458, new_g10401_);
  not g183837 (n_1556, new_g10323_);
  not g183790 (n_2109, g1657);
  not g183786 (n_8069, g1105);
  not g183845 (n_4542, g703);
  not g184011 (n_901, new_g6875_);
  not g184038 (n_8824, g2217);
  not g183831 (n_580, g1783);
  not g183791 (n_472, g1514);
  not g183832 (n_8826, g1792);
  not g183838 (n_2609, g11388);
  not g183775 (n_1040, g5022);
  not g183968 (n_7535, g1024);
  not g184042 (n_1438, new_g7766_);
  not g184008 (n_1805, new_g12440_);
  not g183773 (n_481, new_g10371_);
  not g183778 (n_582, g1592);
  not g184049 (n_2612, g12470);
  not g183935 (n_6890, g1018);
  not g184002 (n_1026, g5084);
  not g183949 (n_4457, g5041);
  not g183840 (n_8825, g2060);
  not g183827 (n_1549, new_g7704_);
  not g183783 (n_1317, g1862);
  not g184055 (n_2621, g11418);
  not g183828 (n_1994, g4878);
  not g184046 (n_4013, g1478);
  not g183823 (n_484, g2227);
  not g184057 (n_5549, g5052);
  not g184064 (n_6361, g4040);
  not g184052 (n_4225, g1448);
  not g184045 (n_2638, g1351);
  not g184013 (n_1891, g5016);
  not g183822 (n_2866, g4643);
  not g183873 (n_113, g441);
  not g183936 (n_111, g2407);
  not g183651 (n_110, g8784);
  not g183756 (n_109, new_g10409_);
  not g183866 (n_108, g218);
  not g183910 (n_107, g17320);
  not g183965 (n_106, g5297);
  not g183690 (n_104, g1124);
  not g183922 (n_103, g1041);
  not g183864 (n_102, g4141);
  not g183931 (n_99, g1221);
  not g183858 (n_96, g2984);
  not g183732 (n_91, g6209);
  not g184029 (n_90, g4601);
  not g183770 (n_88, g1099);
  not g183985 (n_87, g1373);
  not g183918 (n_86, g1152);
  not g183928 (n_85, g2380);
  not g183751 (n_83, g2783);
  not g183709 (n_81, g2079);
  not g184007 (n_80, g5092);
  not g183993 (n_77, g6549);
  not g183905 (n_74, g2375);
  not g183901 (n_72, g2917);
  not g183668 (n_71, g2036);
  not g184005 (n_70, g3155);
  not g183871 (n_68, g2461);
  not g183906 (n_67, g3111);
  not g183634 (n_66, g4119);
  not g183926 (n_63, g142);
  not g183660 (n_62, g2112);
  not g183887 (n_61, g2827);
  not g183892 (n_60, g8789);
  not g183720 (n_59, g1333);
  not g183670 (n_58, g7245);
  not g183780 (n_56, g1087);
  not g183938 (n_54, g12919);
  not g183659 (n_53, g1902);
  not g183852 (n_52, g2873);
  not g183784 (n_50, g5857);
  not g183897 (n_49, g962);
  not g183763 (n_47, g5517);
  not g183987 (n_46, g1996);
  not g183874 (n_44, g4771);
  not g183996 (n_43, g3857);
  not g183908 (n_42, g1495);
  not g183656 (n_41, g2791);
  not g183898 (n_39, g283);
  not g183701 (n_38, g969);
  not g183915 (n_37, g1395);
  not g183627 (n_36, g2980);
  not g183736 (n_35, g2819);
  not g183700 (n_34, g1821);
  not g183911 (n_33, g8786);
  not g183712 (n_32, g4871);
  not g183740 (n_31, new_g8038_);
  not g183633 (n_30, g4492);
  not g183755 (n_29, g822);
  not g183954 (n_27, g20557);
  not g183878 (n_26, g2799);
  not g183961 (n_24, g4264);
  not g183699 (n_23, g2246);
  not g183856 (n_22, g4944);
  not g183643 (n_21, g2066);
  not g183689 (n_20, g4843);
  not g183973 (n_18, g3161);
  not g183753 (n_17, g3863);
  not g183963 (n_16, g6555);
  not g183733 (n_15, g2771);
  not g183750 (n_14, g5863);
  not g183715 (n_13, g146);
  not g183654 (n_12, g2811);
  not g183944 (n_11, g1361);
  not g183776 (n_10, g5164);
  not g184016 (n_9, g837);
  not g183997 (n_7, g1760);
  not g183857 (n_6, g4405);
  not g183782 (n_5, g1430);
  not g183771 (n_4, g1205);
  not g184000 (n_3, g3506);
  not g183902 (n_2, g2767);
  not g183894 (n_1, g1768);
  not g183998 (n_0, g6203);
  not g183754 (n_601, g5057);
  not g183739 (n_1173, g417);
  not g184024 (n_465, g5188);
  not g183820 (n_6311, g2465);
  not g184037 (n_975, g2476);
  not g183992 (n_1651, g370);
  not g183816 (n_511, g4358);
  not g184026 (n_8074, g1135);
  not g183937 (n_2741, g6167);
  not g183960 (n_2862, g6513);
  not g183693 (n_906, g4621);
  not g183789 (n_453, g1624);
  not g183807 (n_452, g2319);
  not g183760 (n_2736, g5128);
  not g184004 (n_912, g4899);
  not g183966 (n_2758, g3821);
  not g183917 (n_534, g164);
  not g183649 (n_626, g4093);
  not g183692 (n_592, g4180);
  not g183801 (n_477, g6219);
  not g183678 (n_2107, g6390);
  not g183764 (n_1433, g1339);
  not g183842 (n_2503, g979);
  not g183734 (n_7571, g2102);
  not g184053 (n_1516, g11349);
  not g183681 (n_1350, g1216);
  not g183774 (n_479, g1183);
  not g183976 (n_461, g1728);
  not g183800 (n_451, g2185);
  not g183982 (n_3739, g832);
  not g183970 (n_469, new_g10366_);
  not g183787 (n_460, g5535);
  not g183841 (n_524, g358);
  not g183716 (n_2088, g3698);
  not g183819 (n_450, g1171);
  not g183741 (n_1085, g2518);
  not g183988 (n_1613, g718);
  not g183844 (n_1593, g12238);
  not g183945 (n_475, new_g10413_);
  not g183813 (n_464, g3171);
  not g183728 (n_7260, g2393);
  not g183818 (n_480, g2028);
  not g183777 (n_962, g4608);
  not g183695 (n_2075, g5698);
  not g183830 (n_1601, g12350);
  not g184048 (n_6309, g2197);
  not g183694 (n_620, g4087);
  not g183808 (n_822, new_g7074_);
  not g184012 (n_467, g6227);
  not g184025 (n_463, g2453);
  not g183836 (n_1299, g4776);
  not g183727 (n_1081, g1825);
  not g183975 (n_1381, g1564);
  not g184020 (n_905, g5873);
  not g183788 (n_474, g5527);
  not g183950 (n_1055, g1036);
  not g183967 (n_1079, g1959);
  not g184027 (n_466, g6565);
  not g184032 (n_1599, g12300);
  not g183812 (n_982, g2070);
  not g183721 (n_6814, g287);
  not g183814 (n_459, new_g7028_);
  not g183846 (n_6560, g3338);
  not g184043 (n_617, g3530);
  not g183796 (n_904, new_g7097_);
  not g184058 (n_1440, new_g7812_);
  not g183804 (n_1005, g2629);
  not g183927 (n_3916, g843);
  not g183843 (n_1442, new_g7791_);
  not g183990 (n_3691, g4311);
  not g183953 (n_957, g385);
  not g183691 (n_2870, g4098);
  not g184044 (n_8829, g2619);
  not g184030 (n_482, new_g6905_);
  not g183798 (n_1011, g2361);
  not g184061 (n_2376, g691);
  not g184051 (n_1551, new_g10295_);
  not g184040 (n_2614, g12422);
  not g184039 (n_1441, new_g7121_);
  not g184034 (n_1550, new_g7738_);
  not g184015 (n_478, new_g7051_);
  not g184060 (n_3512, g4340);
  not g183821 (n_8823, g1926);
  not g184028 (n_908, new_g6928_);
  not g183826 (n_2640, g1008);
  not g184014 (n_816, g3179);
  not g184050 (n_978, g2610);
  not g184033 (n_1445, g4584);
  not g184035 (n_8822, g2351);
  not g183824 (n_913, g4975);
  not g183833 (n_968, g3522);
  not g183825 (n_488, g1802);
  not g183848 (n_6357, g6035);
  not g183794 (n_1916, g5062);
  not g183805 (n_3509, g4322);
  not g183847 (n_6562, g25219);
  not g183829 (n_486, g4785);
  not g184066 (n_6359, g5689);
  not g184047 (n_911, g2495);
  not g183839 (n_4008, g1472);
  not g184067 (n_4492, g6381);
  not g184056 (n_3496, g1322);
  not g184063 (n_6580, g6727);
  not g184059 (n_3986, g4392);
  not g184065 (n_6582, g3689);
  not g184041 (n_5340, g4593);
  not hi_fo_buf185313 (n_9257, g35);
  not g3 (n_10110, n_10109);
  nor g2 (n_10109, g4420, g4427);
  not g185332 (n_10112, n_10111);
  nor g185333 (n_10111, g4242, g4300);
  not g185334 (n_10114, n_10113);
  nor g185335 (n_10113, n_5886, n_8515);
  not g185336 (n_10116, n_10115);
  nor g185337 (n_10115, n_6073, n_8513);
  not g185338 (n_10118, n_10117);
  nor g185339 (n_10117, n_5901, n_8476);
  not g185340 (n_10120, n_10119);
  nor g185341 (n_10119, n_5909, n_8475);
  not g185342 (n_10122, n_10121);
  nor g185343 (n_10121, n_5890, n_8474);
  not g185344 (n_10124, n_10123);
  nor g185345 (n_10123, g355, g333);
  not g185346 (n_10126, n_10125);
  nor g185347 (n_10125, g534, g301);
  not g185348 (n_10128, n_10127);
  nor g185349 (n_10127, n_5900, n_8129);
  nor g185351 (n_10129, n_1216, n_8046);
  nor g185353 (n_10131, n_575, n_8044);
  not g185354 (n_10134, n_10133);
  nor g185355 (n_10133, n_1998, n_7922);
  nor g185357 (n_10135, g8915, g11770);
  not g185358 (n_10138, n_10137);
  nor g185359 (n_10137, n_7537, n_7682);
  not g185362 (n_10142, n_10141);
  nor g185363 (n_10141, n_7193, n_7449);
  not g185364 (n_10144, n_10143);
  nor g185365 (n_10143, n_7170, n_7431);
  not g185366 (n_10146, n_10145);
  nor g185367 (n_10145, n_2382, n_6733);
  not g185368 (n_10148, n_10147);
  nor g185369 (n_10147, n_5872, n_6470);
  not g185370 (n_10150, n_10149);
  nor g185371 (n_10149, n_5813, n_6072);
  not g185372 (n_10152, n_10151);
  nor g185373 (n_10151, n_5707, n_6008);
  not g185374 (n_10154, n_10153);
  nor g185375 (n_10153, n_5687, n_5912);
  not g185376 (n_10156, n_10155);
  nor g185377 (n_10155, n_5654, n_5906);
  not g185378 (n_10158, n_10157);
  nor g185379 (n_10157, n_5630, n_5902);
  not g185380 (n_10160, n_10159);
  nor g185381 (n_10159, n_5604, n_5898);
  not g185382 (n_10162, n_10161);
  nor g185383 (n_10161, n_5668, n_5894);
  not g185384 (n_10164, n_10163);
  nor g185385 (n_10163, n_5572, n_5887);
  nor g185387 (n_10165, g5142, n_6268);
  nor g185389 (n_10167, g6181, n_6271);
  nor g185391 (n_10169, g3484, n_6274);
  not g185392 (g26876, n_10171);
  nor g185393 (n_10171, n_5329, n_5324);
  nor g185395 (n_10173, g3133, n_5776);
  nor g185397 (n_10175, g6527, n_5770);
  nor g185399 (n_10177, g5489, n_5767);
  nor g185401 (n_10179, g5835, n_5783);
  nor g185403 (n_10181, g3835, n_5773);
  nor g185405 (n_10183, g490, n_4696);
  not g185406 (n_10186, n_10185);
  nor g185407 (n_10185, new_g6946_, g4253);
  not g185408 (n_10188, n_10187);
  nor g185409 (n_10187, new_g10354_, n_4373);
  not g185410 (n_10190, n_10189);
  nor g185411 (n_10189, g278, n_4181);
  not g185412 (n_10192, n_10191);
  nor g185413 (n_10191, g4417, n_4106);
  not g185414 (n_10194, n_10193);
  nor g185415 (n_10193, n_1797, n_4079);
  not g185416 (n_10196, n_10195);
  nor g185417 (n_10195, n_3183, n_3265);
  not g185418 (n_10198, n_10197);
  nor g185419 (n_10197, n_2806, n_3202);
  not g185420 (n_10200, n_10199);
  nor g185421 (n_10199, n_2802, n_3147);
  not g185422 (n_10202, n_10201);
  nor g185423 (n_10201, n_2763, n_3137);
  not g185424 (n_10204, n_10203);
  nor g185425 (n_10203, n_2837, n_3132);
  not g185426 (n_10206, n_10205);
  nor g185427 (n_10205, n_2732, n_3116);
  not g185428 (n_10208, n_10207);
  nor g185429 (n_10207, n_2842, n_3094);
  not g185430 (g26875, n_10209);
  nor g185431 (n_10209, n_3408, n_3410);
  not g185432 (n_10212, n_10211);
  nor g185433 (n_10211, g2886, g2946);
  nor g185435 (n_10213, g1559, n_10220);
  not g185436 (n_10216, n_10215);
  nor g185437 (n_10215, n_2002, n_2840);
  not g185438 (n_10218, n_10217);
  nor g185439 (n_10217, n_4193, n_3387);
  not g185440 (n_10220, n_10219);
  nor g185441 (n_10219, g1554, n_2317);
  not g185442 (n_10222, n_10221);
  nor g185443 (n_10221, n_2047, n_2193);
  nor g185445 (n_10223, n_2191, n_2189);
  not g185448 (n_10228, n_10227);
  nor g185449 (n_10227, n_1324, n_1355);
  nor g185451 (n_10229, g1858, g1724);
  not g185452 (n_10232, n_10231);
  nor g185453 (n_10231, g5152, g5138);
  nor g185455 (n_10233, g1664, g1644);
  nor g185457 (n_10235, g1830, g1696);
  not g185458 (n_10238, n_10237);
  nor g185459 (n_10237, g3845, g3831);
  not g185460 (n_10240, n_10239);
  nor g185461 (n_10239, g3143, g3129);
  not g185462 (n_10242, n_10241);
  nor g185463 (n_10241, g3494, g3480);
  not g185464 (n_10244, n_10243);
  nor g185465 (n_10243, g5845, g5831);
  nor g185467 (n_10245, g2389, g2255);
  nor g185469 (n_10247, g2417, g2283);
  not g185470 (n_10250, n_10249);
  nor g185471 (n_10249, g5499, g5485);
  not g185472 (n_10252, n_10251);
  nor g185473 (n_10251, g6191, g6177);
  not g185474 (n_10254, n_10253);
  nor g185475 (n_10253, g6537, g6523);
  not g185476 (n_10256, n_10255);
  nor g185477 (n_10255, n_10129, n_8157);
  not g185478 (n_10258, n_10257);
  nor g185479 (n_10257, n_10131, n_8158);
  nand g185480 (n_10260, n_1733, n_10412);
  nor g185482 (n_10262, g2527, n_10261);
  nand g185483 (n_10261, n_8986, g35);
  nor g185485 (n_10265, g1700, n_10264);
  nand g185486 (n_10264, n_8993, g35);
  nor g185488 (n_10268, g1834, n_10267);
  nand g185489 (n_10267, n_8995, g35);
  nor g185491 (n_10271, g1968, n_10270);
  nand g185492 (n_10270, n_8997, g35);
  nor g185494 (n_10274, g2259, n_10273);
  nand g185495 (n_10273, n_9002, g35);
  nor g185497 (n_10277, n_8610, n_10276);
  nand g185498 (n_10276, g35, g2389);
  nor g185500 (n_10280, n_8614, n_10279);
  nand g185501 (n_10279, g35, g2255);
  nor g185503 (n_10283, n_8612, n_10282);
  nand g185504 (n_10282, g35, g1696);
  nand g185505 (n_10286, n_8219, n_10285);
  wire w299, w300, w301, w302;
  nand g185506 (n_10285, w300, w302);
  nand g348 (w302, w301, g4430);
  not g346 (w301, n_1694);
  nand g345 (w300, w299, n_1694);
  not g344 (w299, g4430);
  nand g185507 (n_10288, n_4812, n_10287);
  nor g185508 (n_10287, n_8126, n_5416);
  nand g185509 (n_10290, n_4801, n_10289);
  nor g185510 (n_10289, n_8115, n_5410);
  nor g185512 (n_10292, n_10327, n_10291);
  nand g185513 (n_10291, n_4880, g35);
  nor g185514 (n_10295, n_7933, n_10294);
  nand g185515 (n_10294, n_7507, n_7645);
  nand g185516 (n_10297, n_4435, n_10296);
  nor g185517 (n_10296, n_7989, n_7869);
  nor g185518 (n_10299, n_7939, n_10298);
  nand g185519 (n_10298, n_7866, n_7634);
  nand g185520 (n_10301, n_10135, n_10300);
  nor g185521 (n_10300, g8917, g8916);
  not g185522 (n_10304, n_10303);
  nor g185523 (n_10303, n_3519, n_10302);
  nand g185524 (n_10302, n_5243, n_7927);
  not g185525 (n_10307, n_10306);
  nor g185526 (n_10306, n_3024, n_10305);
  nand g185527 (n_10305, n_5011, n_7926);
  nand g185528 (n_10309, n_7643, n_10308);
  nor g185529 (n_10308, n_7115, n_5296);
  not g185530 (n_10312, n_10311);
  nor g185531 (n_10311, n_3027, n_10310);
  nand g185532 (n_10310, n_5270, n_7876);
  nor g185534 (n_10314, n_7487, n_10313);
  nand g185535 (n_10313, g35, g1870);
  not g185536 (n_10318, n_10317);
  nor g185537 (n_10317, n_3517, n_10316);
  nand g185538 (n_10316, n_5240, n_7874);
  not g185539 (n_10321, n_10320);
  nor g185540 (n_10320, n_3077, n_10319);
  nand g185541 (n_10319, n_5023, n_7875);
  nor g185543 (n_10323, n_7418, n_10322);
  nand g185544 (n_10322, n_8214, g164);
  not g185545 (n_10327, n_10326);
  nor g185546 (n_10326, g13259, n_10325);
  nand g185547 (n_10325, n_7530, n_1598);
  nor g185549 (n_10329, n_7151, n_10328);
  nand g185550 (n_10328, g35, g1600);
  nor g185552 (n_10332, n_6933, n_10331);
  nand g185553 (n_10331, g35, g2004);
  not g185554 (n_10336, n_10335);
  nor g185555 (n_10335, n_10167, n_10334);
  nand g185556 (n_10334, n_6254, n_919);
  not g185557 (n_10339, n_10338);
  nor g185558 (n_10338, n_10169, n_10337);
  nand g185559 (n_10337, n_6253, n_1187);
  not g185560 (n_10342, n_10341);
  nor g185561 (n_10341, n_10165, n_10340);
  nand g185562 (n_10340, n_6252, n_1134);
  nor g185564 (n_10344, n_6394, n_10343);
  nand g185565 (n_10343, g35, g2563);
  nor g185567 (n_10347, n_6392, n_10346);
  nand g185568 (n_10346, g35, g2295);
  not g185569 (n_10351, n_10350);
  nor g185570 (n_10350, n_10181, n_10349);
  nand g185571 (n_10349, n_6231, n_781);
  not g185572 (n_10354, n_10353);
  nor g185573 (n_10353, n_10173, n_10352);
  nand g185574 (n_10352, n_6244, n_1225);
  not g185575 (n_10357, n_10356);
  nor g185576 (n_10356, n_10175, n_10355);
  nand g185577 (n_10355, n_6225, n_728);
  not g185578 (n_10360, n_10359);
  nor g185579 (n_10359, n_10179, n_10358);
  nand g185580 (n_10358, n_6237, n_603);
  not g185581 (n_10363, n_10362);
  nor g185582 (n_10362, n_10177, n_10361);
  nand g185583 (n_10361, n_6242, n_949);
  not g185584 (n_10366, n_10365);
  nor g185585 (n_10365, n_10183, n_10364);
  nand g185586 (n_10364, n_6190, n_774);
  not g185587 (n_10369, n_10368);
  nor g185588 (n_10368, n_4283, n_10367);
  nand g185589 (n_10367, n_4560, g732);
  nor g185591 (n_10371, g311, n_10370);
  nand g185592 (n_10370, g35, g324);
  not g185593 (n_10375, n_10374);
  nor g185594 (n_10374, n_10213, n_10373);
  nand g185595 (n_10373, n_3606, n_685);
  not g185596 (n_10378, n_10377);
  nor g185597 (n_10377, n_10223, n_10376);
  nand g185598 (n_10376, n_4193, n_3387);
  nand g185599 (n_10380, n_382, n_10379);
  nor g185600 (n_10379, n_3112, n_1564);
  nand g185601 (n_10382, n_2448, n_10381);
  nor g185602 (n_10381, n_2846, n_2845);
  nor g185604 (n_10384, g5033, n_10383);
  nand g185605 (n_10383, n_2650, g35);
  nand g185606 (n_10387, n_10247, n_10386);
  nor g185607 (n_10386, g2685, g2551);
  nand g185608 (n_10389, n_10233, n_10388);
  nor g185609 (n_10388, g1798, g1779);
  nand g185610 (n_10391, n_10235, n_10390);
  nor g185611 (n_10390, g2098, g1964);
  nand g185612 (n_10393, n_1352, n_10392);
  nor g185613 (n_10392, g411, n_1934);
  nand g185614 (n_10395, n_10245, n_10394);
  nor g185615 (n_10394, g2657, g2523);
  nand g185616 (n_10397, n_10229, n_10396);
  nor g185617 (n_10396, g2126, g1992);
  not g185618 (n_10400, n_10399);
  nor g185619 (n_10399, g13272, n_10398);
  nand g185620 (n_10398, n_1512, n_291);
  not g185621 (n_10403, n_10402);
  nor g185622 (n_10402, g1691, n_10401);
  nand g185623 (n_10401, g35, g1687);
  not g185624 (n_10406, n_10405);
  nor g185625 (n_10405, g2384, n_10404);
  nand g185626 (n_10404, g35, g2380);
  not g185627 (n_10409, n_10408);
  nor g185628 (n_10408, g2250, n_10407);
  nand g185629 (n_10407, g35, g2246);
  not g185630 (n_10412, n_10411);
  nand g185631 (n_10411, n_7387, n_10410);
  wire w303, w304, w305, w306;
  nand g185632 (n_10410, w304, w306);
  nand g353 (w306, w305, g1061);
  not g352 (w305, n_1458);
  nand g350 (w304, w303, n_1458);
  not g349 (w303, g1061);
  not g185633 (n_10414, n_10413);
  nor g185634 (n_10413, n_8789, n_10283);
  not g185635 (n_10416, n_10415);
  nor g185636 (n_10415, n_8784, n_10280);
  not g185637 (n_10418, n_10417);
  nor g185638 (n_10417, n_8805, n_10277);
  not g185639 (n_10420, n_10419);
  nor g185640 (n_10419, n_7814, n_10314);
  not g185641 (n_10422, n_10421);
  nor g185642 (n_10421, n_7676, n_10323);
  not g185643 (n_10424, n_10423);
  nor g185644 (n_10423, n_7644, n_10329);
  not g185645 (n_10426, n_10425);
  nor g185646 (n_10425, n_10332, n_7435);
  not g185647 (n_10428, n_10427);
  nor g185648 (n_10427, n_10344, n_7116);
  not g185649 (n_10430, n_10429);
  nor g185650 (n_10429, n_10347, n_7106);
  not g185651 (n_10432, n_10431);
  nor g185652 (n_10431, n_10384, n_5918);
  not g185653 (n_10435, n_10434);
  nor g185654 (n_10434, n_10265, n_10433);
  nand g185655 (n_10433, n_9105, n_586);
  not g185656 (n_10438, n_10437);
  nor g185657 (n_10437, n_10268, n_10436);
  nand g185658 (n_10436, n_9091, n_1239);
  not g185659 (n_10441, n_10440);
  nor g185660 (n_10440, n_10271, n_10439);
  nand g185661 (n_10439, n_9103, n_718);
  not g185662 (n_10444, n_10443);
  nor g185663 (n_10443, n_10262, n_10442);
  nand g185664 (n_10442, n_9107, n_787);
  not g4 (n_10447, n_10446);
  nor g185665 (n_10446, n_10274, n_10445);
  nand g185666 (n_10445, n_9101, n_678);
  not g185667 (n_10450, n_10449);
  nor g185668 (n_10449, n_10292, n_10448);
  nand g185669 (n_10448, n_8043, n_1144);
  not g185670 (n_10453, n_10452);
  nor g185671 (n_10452, n_10371, n_10451);
  nand g185672 (n_10451, n_6494, n_887);
endmodule


module fflopd(CK, D, Q);
  input CK, D;
  output Q;
  wire CK, D;
  wire Q;
  wire next_state;
  reg  qi;
  assign #1 Q = qi;
  assign next_state = D;
  always 
    @(posedge CK) 
      qi <= next_state;
  initial 
    qi <= 1'b0;
endmodule