module multiplier(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6]
     , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] ,
     \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] ,
     \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] ,
     \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] ,
     \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] ,
     \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
     \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
     \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] ,
     \a[63] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] ,
     \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14]
     , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] , \b[21] ,
     \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
     \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
     \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] ,
     \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
     \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
     \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
     \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
     \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] ,
     \f[15] , \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] ,
     \f[22] , \f[23] , \f[24] , \f[25] , \f[26] , \f[27] , \f[28] ,
     \f[29] , \f[30] , \f[31] , \f[32] , \f[33] , \f[34] , \f[35] ,
     \f[36] , \f[37] , \f[38] , \f[39] , \f[40] , \f[41] , \f[42] ,
     \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] , \f[49] ,
     \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
     \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
     \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] ,
     \f[71] , \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] ,
     \f[78] , \f[79] , \f[80] , \f[81] , \f[82] , \f[83] , \f[84] ,
     \f[85] , \f[86] , \f[87] , \f[88] , \f[89] , \f[90] , \f[91] ,
     \f[92] , \f[93] , \f[94] , \f[95] , \f[96] , \f[97] , \f[98] ,
     \f[99] , \f[100] , \f[101] , \f[102] , \f[103] , \f[104] , \f[105]
     , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] , \f[111] ,
     \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
     \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
     \f[124] , \f[125] , \f[126] , \f[127] );
  input \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
       \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] ,
       \b[8] , \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] ,
       \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] , \b[21] ,
       \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
       \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
       \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] ,
       \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
       \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
       \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7]
       , \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] ,
       \f[15] , \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] ,
       \f[22] , \f[23] , \f[24] , \f[25] , \f[26] , \f[27] , \f[28] ,
       \f[29] , \f[30] , \f[31] , \f[32] , \f[33] , \f[34] , \f[35] ,
       \f[36] , \f[37] , \f[38] , \f[39] , \f[40] , \f[41] , \f[42] ,
       \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] , \f[49] ,
       \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
       \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
       \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] ,
       \f[71] , \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] ,
       \f[78] , \f[79] , \f[80] , \f[81] , \f[82] , \f[83] , \f[84] ,
       \f[85] , \f[86] , \f[87] , \f[88] , \f[89] , \f[90] , \f[91] ,
       \f[92] , \f[93] , \f[94] , \f[95] , \f[96] , \f[97] , \f[98] ,
       \f[99] , \f[100] , \f[101] , \f[102] , \f[103] , \f[104] ,
       \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
       \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
       \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] ,
       \f[123] , \f[124] , \f[125] , \f[126] , \f[127] ;
  wire \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
       \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] ,
       \b[8] , \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] ,
       \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] , \b[21] ,
       \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
       \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
       \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] ,
       \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
       \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
       \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  wire \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
       \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] ,
       \f[15] , \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] ,
       \f[22] , \f[23] , \f[24] , \f[25] , \f[26] , \f[27] , \f[28] ,
       \f[29] , \f[30] , \f[31] , \f[32] , \f[33] , \f[34] , \f[35] ,
       \f[36] , \f[37] , \f[38] , \f[39] , \f[40] , \f[41] , \f[42] ,
       \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] , \f[49] ,
       \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
       \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
       \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] ,
       \f[71] , \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] ,
       \f[78] , \f[79] , \f[80] , \f[81] , \f[82] , \f[83] , \f[84] ,
       \f[85] , \f[86] , \f[87] , \f[88] , \f[89] , \f[90] , \f[91] ,
       \f[92] , \f[93] , \f[94] , \f[95] , \f[96] , \f[97] , \f[98] ,
       \f[99] , \f[100] , \f[101] , \f[102] , \f[103] , \f[104] ,
       \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
       \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
       \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] ,
       \f[123] , \f[124] , \f[125] , \f[126] , \f[127] ;
  wire n257, n258, n259, n261, n262, n263, n264, n265;
  wire n266, n267, n268, n269, n270, n271, n272, n273;
  wire n274, n275, n276, n277, n278, n279, n280, n282;
  wire n283, n284, n285, n286, n289, n290, n291, n292;
  wire n293, n294, n295, n296, n297, n298, n299, n300;
  wire n301, n302, n303, n304, n306, n307, n308, n311;
  wire n312, n313, n314, n315, n316, n317, n318, n319;
  wire n320, n321, n322, n323, n324, n325, n326, n327;
  wire n328, n329, n330, n331, n332, n333, n335, n336;
  wire n337, n340, n341, n342, n343, n344, n345, n346;
  wire n347, n348, n349, n350, n351, n352, n353, n354;
  wire n355, n356, n357, n358, n359, n360, n361, n362;
  wire n363, n364, n365, n366, n367, n368, n369, n370;
  wire n371, n372, n373, n374, n375, n376, n377, n378;
  wire n379, n380, n381, n383, n384, n385, n388, n389;
  wire n390, n391, n392, n393, n394, n395, n396, n397;
  wire n398, n399, n400, n401, n402, n403, n404, n405;
  wire n406, n407, n408, n409, n410, n411, n412, n413;
  wire n414, n415, n416, n417, n418, n419, n420, n421;
  wire n422, n423, n425, n426, n427, n428, n429, n430;
  wire n431, n432, n433, n434, n435, n436, n439, n440;
  wire n441, n442, n443, n444, n445, n446, n447, n448;
  wire n449, n450, n453, n454, n455, n456, n457, n458;
  wire n459, n460, n461, n462, n463, n464, n465, n466;
  wire n467, n468, n469, n470, n472, n473, n474, n475;
  wire n478, n479, n480, n481, n482, n483, n484, n485;
  wire n486, n487, n488, n489, n490, n491, n492, n493;
  wire n496, n497, n498, n499, n500, n501, n502, n503;
  wire n504, n505, n506, n507, n508, n509, n510, n511;
  wire n512, n513, n514, n515, n516, n517, n518, n519;
  wire n520, n521, n522, n523, n524, n525, n526, n527;
  wire n528, n529, n530, n531, n532, n533, n534, n535;
  wire n536, n537, n539, n540, n541, n542, n543, n546;
  wire n547, n548, n549, n550, n551, n552, n553, n554;
  wire n555, n556, n557, n560, n561, n562, n563, n564;
  wire n565, n566, n567, n568, n569, n570, n571, n572;
  wire n573, n574, n575, n576, n579, n580, n581, n582;
  wire n583, n584, n585, n586, n587, n588, n589, n590;
  wire n591, n592, n593, n594, n595, n596, n597, n598;
  wire n600, n601, n602, n605, n606, n607, n608, n609;
  wire n610, n611, n612, n613, n614, n615, n616, n617;
  wire n618, n619, n620, n623, n624, n625, n626, n627;
  wire n628, n629, n630, n631, n632, n633, n634, n635;
  wire n636, n637, n638, n639, n640, n641, n642, n645;
  wire n646, n647, n648, n649, n650, n651, n652, n653;
  wire n654, n655, n656, n657, n658, n659, n660, n661;
  wire n662, n663, n664, n666, n667, n668, n669, n672;
  wire n673, n674, n675, n676, n677, n678, n679, n680;
  wire n681, n682, n685, n686, n687, n688, n689, n690;
  wire n691, n692, n693, n694, n695, n696, n697, n698;
  wire n699, n700, n701, n702, n703, n704, n705, n706;
  wire n707, n708, n709, n710, n711, n712, n713, n714;
  wire n715, n716, n717, n718, n719, n720, n721, n722;
  wire n723, n724, n725, n726, n727, n728, n729, n732;
  wire n733, n734, n735, n736, n737, n738, n739, n740;
  wire n741, n742, n743, n744, n745, n746, n747, n748;
  wire n749, n751, n752, n753, n754, n755, n758, n759;
  wire n760, n761, n762, n763, n764, n765, n766, n767;
  wire n768, n769, n772, n773, n774, n775, n776, n777;
  wire n778, n779, n780, n781, n782, n783, n786, n787;
  wire n788, n789, n790, n791, n792, n793, n794, n795;
  wire n796, n797, n798, n799, n800, n801, n802, n803;
  wire n804, n805, n806, n807, n808, n809, n812, n813;
  wire n814, n815, n816, n817, n818, n819, n820, n821;
  wire n822, n823, n824, n825, n826, n827, n828, n829;
  wire n831, n832, n833, n836, n837, n838, n839, n840;
  wire n841, n842, n843, n844, n845, n846, n847, n848;
  wire n849, n850, n851, n854, n855, n856, n857, n858;
  wire n859, n860, n861, n862, n863, n864, n865, n866;
  wire n867, n868, n869, n872, n873, n874, n875, n876;
  wire n877, n878, n879, n880, n881, n882, n883, n884;
  wire n885, n886, n887, n888, n889, n890, n891, n894;
  wire n895, n896, n897, n898, n899, n900, n901, n902;
  wire n903, n904, n905, n906, n907, n908, n909, n910;
  wire n911, n912, n913, n914, n916, n917, n918, n919;
  wire n920, n923, n924, n925, n926, n927, n928, n929;
  wire n930, n931, n932, n933, n936, n937, n938, n939;
  wire n940, n941, n942, n943, n944, n945, n946, n947;
  wire n948, n949, n950, n951, n952, n953, n954, n955;
  wire n956, n957, n958, n959, n960, n961, n962, n963;
  wire n964, n965, n966, n967, n968, n969, n970, n971;
  wire n972, n973, n974, n975, n976, n977, n978, n979;
  wire n980, n983, n984, n985, n986, n987, n988, n989;
  wire n990, n991, n992, n993, n994, n995, n996, n997;
  wire n998, n999, n1002, n1003, n1004, n1005, n1006, n1007;
  wire n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015;
  wire n1016, n1017, n1018, n1019, n1021, n1022, n1023, n1024;
  wire n1025, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  wire n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
  wire n1043, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
  wire n1053, n1054, n1055, n1056, n1057, n1058, n1061, n1062;
  wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
  wire n1071, n1072, n1075, n1076, n1077, n1078, n1079, n1080;
  wire n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088;
  wire n1089, n1090, n1091, n1094, n1095, n1096, n1097, n1098;
  wire n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106;
  wire n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114;
  wire n1115, n1116, n1118, n1119, n1120, n1121, n1122, n1125;
  wire n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133;
  wire n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141;
  wire n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151;
  wire n1152, n1153, n1156, n1157, n1158, n1159, n1160, n1161;
  wire n1162, n1163, n1164, n1167, n1168, n1169, n1170, n1171;
  wire n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179;
  wire n1180, n1181, n1182, n1185, n1186, n1187, n1188, n1189;
  wire n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
  wire n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205;
  wire n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
  wire n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221;
  wire n1222, n1223, n1225, n1226, n1227, n1228, n1231, n1232;
  wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240;
  wire n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1250;
  wire n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258;
  wire n1259, n1262, n1263, n1264, n1265, n1266, n1267, n1268;
  wire n1269, n1270, n1271, n1274, n1275, n1276, n1277, n1278;
  wire n1279, n1280, n1281, n1282, n1283, n1284, n1287, n1288;
  wire n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296;
  wire n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304;
  wire n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312;
  wire n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;
  wire n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;
  wire n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;
  wire n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1345;
  wire n1346, n1347, n1350, n1351, n1352, n1353, n1354, n1355;
  wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
  wire n1364, n1365, n1366, n1369, n1370, n1371, n1372, n1373;
  wire n1374, n1375, n1376, n1377, n1378, n1381, n1382, n1383;
  wire n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391;
  wire n1392, n1393, n1396, n1397, n1398, n1399, n1400, n1401;
  wire n1402, n1403, n1404, n1405, n1406, n1407, n1410, n1411;
  wire n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419;
  wire n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1429;
  wire n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;
  wire n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445;
  wire n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453;
  wire n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1462;
  wire n1463, n1464, n1465, n1468, n1469, n1470, n1471, n1472;
  wire n1473, n1474, n1475, n1476, n1477, n1480, n1481, n1482;
  wire n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1492;
  wire n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500;
  wire n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1510;
  wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
  wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
  wire n1527, n1528, n1531, n1532, n1533, n1534, n1535, n1536;
  wire n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544;
  wire n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552;
  wire n1553, n1554, n1555, n1556, n1557, n1560, n1561, n1562;
  wire n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570;
  wire n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578;
  wire n1579, n1581, n1582, n1583, n1586, n1587, n1588, n1589;
  wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1599;
  wire n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607;
  wire n1608, n1609, n1612, n1613, n1614, n1615, n1616, n1617;
  wire n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625;
  wire n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633;
  wire n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641;
  wire n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649;
  wire n1650, n1651, n1652, n1653, n1654, n1657, n1658, n1659;
  wire n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667;
  wire n1668, n1669, n1670, n1671, n1672, n1673, n1676, n1677;
  wire n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685;
  wire n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693;
  wire n1694, n1695, n1696, n1697, n1698, n1699, n1702, n1703;
  wire n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711;
  wire n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719;
  wire n1720, n1721, n1723, n1724, n1725, n1726, n1729, n1730;
  wire n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1740;
  wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
  wire n1749, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
  wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1768;
  wire n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776;
  wire n1777, n1778, n1779, n1782, n1783, n1784, n1785, n1786;
  wire n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794;
  wire n1795, n1796, n1797, n1798, n1801, n1802, n1803, n1804;
  wire n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812;
  wire n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820;
  wire n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828;
  wire n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836;
  wire n1837, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
  wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
  wire n1855, n1856, n1857, n1858, n1859, n1861, n1862, n1863;
  wire n1864, n1867, n1868, n1869, n1870, n1871, n1872, n1873;
  wire n1874, n1875, n1876, n1879, n1880, n1881, n1882, n1883;
  wire n1884, n1885, n1886, n1887, n1888, n1891, n1892, n1893;
  wire n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901;
  wire n1902, n1903, n1904, n1905, n1906, n1909, n1910, n1911;
  wire n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919;
  wire n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927;
  wire n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937;
  wire n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945;
  wire n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953;
  wire n1954, n1955, n1956, n1959, n1960, n1961, n1962, n1963;
  wire n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971;
  wire n1972, n1973, n1974, n1975, n1978, n1979, n1980, n1981;
  wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
  wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997;
  wire n1999, n2000, n2001, n2002, n2003, n2006, n2007, n2008;
  wire n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016;
  wire n2017, n2020, n2021, n2022, n2023, n2024, n2025, n2026;
  wire n2027, n2028, n2029, n2030, n2033, n2034, n2035, n2036;
  wire n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044;
  wire n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052;
  wire n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060;
  wire n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068;
  wire n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2078;
  wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
  wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
  wire n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104;
  wire n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112;
  wire n2113, n2114, n2115, n2116, n2117, n2120, n2121, n2122;
  wire n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130;
  wire n2131, n2132, n2133, n2134, n2135, n2136, n2139, n2140;
  wire n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148;
  wire n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156;
  wire n2158, n2159, n2160, n2161, n2164, n2165, n2166, n2167;
  wire n2168, n2169, n2170, n2171, n2172, n2175, n2176, n2177;
  wire n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2187;
  wire n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195;
  wire n2196, n2197, n2198, n2199, n2200, n2203, n2204, n2205;
  wire n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213;
  wire n2214, n2217, n2218, n2219, n2220, n2221, n2222, n2223;
  wire n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231;
  wire n2232, n2233, n2236, n2237, n2238, n2239, n2240, n2241;
  wire n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249;
  wire n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257;
  wire n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265;
  wire n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2275;
  wire n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283;
  wire n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291;
  wire n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301;
  wire n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;
  wire n2310, n2311, n2312, n2313, n2315, n2316, n2317, n2318;
  wire n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328;
  wire n2329, n2330, n2333, n2334, n2335, n2336, n2337, n2338;
  wire n2339, n2340, n2341, n2342, n2345, n2346, n2347, n2348;
  wire n2349, n2350, n2351, n2352, n2353, n2354, n2357, n2358;
  wire n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366;
  wire n2367, n2368, n2369, n2370, n2371, n2372, n2375, n2376;
  wire n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384;
  wire n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392;
  wire n2393, n2396, n2397, n2398, n2399, n2400, n2401, n2402;
  wire n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410;
  wire n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418;
  wire n2419, n2420, n2421, n2422, n2423, n2424, n2427, n2428;
  wire n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436;
  wire n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444;
  wire n2445, n2446, n2447, n2448, n2449, n2452, n2453, n2454;
  wire n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462;
  wire n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470;
  wire n2471, n2473, n2474, n2475, n2476, n2479, n2480, n2481;
  wire n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489;
  wire n2490, n2491, n2492, n2493, n2494, n2495, n2498, n2499;
  wire n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507;
  wire n2508, n2511, n2512, n2513, n2514, n2515, n2516, n2517;
  wire n2518, n2519, n2520, n2521, n2524, n2525, n2526, n2527;
  wire n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535;
  wire n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543;
  wire n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551;
  wire n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559;
  wire n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2569;
  wire n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577;
  wire n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585;
  wire n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595;
  wire n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603;
  wire n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611;
  wire n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621;
  wire n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629;
  wire n2630, n2631, n2634, n2635, n2636, n2637, n2638, n2639;
  wire n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647;
  wire n2648, n2649, n2650, n2652, n2653, n2654, n2655, n2656;
  wire n2657, n2658, n2659, n2662, n2663, n2664, n2665, n2666;
  wire n2667, n2668, n2669, n2670, n2671, n2674, n2675, n2676;
  wire n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684;
  wire n2685, n2686, n2687, n2690, n2691, n2692, n2693, n2694;
  wire n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2704;
  wire n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712;
  wire n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720;
  wire n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730;
  wire n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738;
  wire n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746;
  wire n2747, n2748, n2749, n2750, n2753, n2754, n2755, n2756;
  wire n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764;
  wire n2765, n2766, n2767, n2770, n2771, n2772, n2773, n2774;
  wire n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782;
  wire n2783, n2784, n2785, n2786, n2789, n2790, n2791, n2792;
  wire n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800;
  wire n2801, n2802, n2803, n2804, n2807, n2808, n2809, n2810;
  wire n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818;
  wire n2819, n2820, n2821, n2822, n2823, n2824, n2826, n2827;
  wire n2828, n2829, n2832, n2833, n2834, n2835, n2836, n2837;
  wire n2838, n2839, n2840, n2843, n2844, n2845, n2846, n2847;
  wire n2848, n2849, n2850, n2851, n2852, n2855, n2856, n2857;
  wire n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2867;
  wire n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875;
  wire n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2885;
  wire n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893;
  wire n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901;
  wire n2902, n2903, n2906, n2907, n2908, n2909, n2910, n2911;
  wire n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919;
  wire n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927;
  wire n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935;
  wire n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945;
  wire n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953;
  wire n2954, n2957, n2958, n2959, n2960, n2961, n2962, n2963;
  wire n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971;
  wire n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979;
  wire n2980, n2981, n2984, n2985, n2986, n2987, n2988, n2989;
  wire n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997;
  wire n2998, n2999, n3000, n3001, n3003, n3004, n3005, n3006;
  wire n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016;
  wire n3017, n3018, n3019, n3022, n3023, n3024, n3025, n3026;
  wire n3027, n3028, n3029, n3030, n3031, n3032, n3035, n3036;
  wire n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044;
  wire n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052;
  wire n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060;
  wire n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068;
  wire n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076;
  wire n3077, n3080, n3081, n3082, n3083, n3084, n3085, n3086;
  wire n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094;
  wire n3095, n3096, n3099, n3100, n3101, n3102, n3103, n3104;
  wire n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112;
  wire n3113, n3114, n3115, n3116, n3119, n3120, n3121, n3122;
  wire n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130;
  wire n3131, n3132, n3133, n3134, n3135, n3138, n3139, n3140;
  wire n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148;
  wire n3149, n3150, n3151, n3152, n3153, n3154, n3157, n3158;
  wire n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166;
  wire n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174;
  wire n3175, n3176, n3177, n3178, n3179, n3180, n3183, n3184;
  wire n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192;
  wire n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200;
  wire n3202, n3203, n3204, n3205, n3208, n3209, n3210, n3211;
  wire n3212, n3213, n3214, n3215, n3216, n3217, n3220, n3221;
  wire n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229;
  wire n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239;
  wire n3240, n3241, n3242, n3243, n3244, n3245, n3248, n3249;
  wire n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257;
  wire n3258, n3259, n3262, n3263, n3264, n3265, n3266, n3267;
  wire n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275;
  wire n3276, n3277, n3278, n3281, n3282, n3283, n3284, n3285;
  wire n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293;
  wire n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301;
  wire n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309;
  wire n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319;
  wire n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327;
  wire n3328, n3331, n3332, n3333, n3334, n3335, n3336, n3337;
  wire n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345;
  wire n3346, n3347, n3350, n3351, n3352, n3353, n3354, n3355;
  wire n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363;
  wire n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371;
  wire n3372, n3373, n3374, n3377, n3378, n3379, n3380, n3381;
  wire n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389;
  wire n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3398;
  wire n3399, n3400, n3401, n3404, n3405, n3406, n3407, n3408;
  wire n3409, n3410, n3411, n3412, n3413, n3416, n3417, n3418;
  wire n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3428;
  wire n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436;
  wire n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3446;
  wire n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454;
  wire n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462;
  wire n3463, n3464, n3467, n3468, n3469, n3470, n3471, n3472;
  wire n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480;
  wire n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488;
  wire n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3498;
  wire n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506;
  wire n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514;
  wire n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524;
  wire n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532;
  wire n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542;
  wire n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3552;
  wire n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560;
  wire n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568;
  wire n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578;
  wire n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586;
  wire n3587, n3588, n3589, n3590, n3592, n3593, n3594, n3597;
  wire n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605;
  wire n3606, n3607, n3610, n3611, n3612, n3613, n3614, n3615;
  wire n3616, n3617, n3618, n3619, n3620, n3623, n3624, n3625;
  wire n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633;
  wire n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641;
  wire n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649;
  wire n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657;
  wire n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665;
  wire n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675;
  wire n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683;
  wire n3684, n3687, n3688, n3689, n3690, n3691, n3692, n3693;
  wire n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701;
  wire n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709;
  wire n3710, n3713, n3714, n3715, n3716, n3717, n3718, n3719;
  wire n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727;
  wire n3728, n3729, n3732, n3733, n3734, n3735, n3736, n3737;
  wire n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745;
  wire n3746, n3747, n3748, n3749, n3752, n3753, n3754, n3755;
  wire n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763;
  wire n3764, n3765, n3766, n3767, n3768, n3771, n3772, n3773;
  wire n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781;
  wire n3782, n3783, n3784, n3785, n3786, n3787, n3790, n3791;
  wire n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799;
  wire n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807;
  wire n3808, n3809, n3811, n3812, n3813, n3814, n3815, n3818;
  wire n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826;
  wire n3827, n3828, n3831, n3832, n3833, n3834, n3835, n3836;
  wire n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844;
  wire n3845, n3848, n3849, n3850, n3851, n3852, n3853, n3854;
  wire n3855, n3856, n3857, n3858, n3859, n3862, n3863, n3864;
  wire n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872;
  wire n3873, n3874, n3875, n3876, n3877, n3878, n3881, n3882;
  wire n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890;
  wire n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3900;
  wire n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908;
  wire n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916;
  wire n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926;
  wire n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934;
  wire n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3944;
  wire n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952;
  wire n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960;
  wire n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970;
  wire n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978;
  wire n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3988;
  wire n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996;
  wire n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004;
  wire n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014;
  wire n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022;
  wire n4023, n4024, n4026, n4027, n4028, n4029, n4030, n4033;
  wire n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041;
  wire n4042, n4043, n4044, n4047, n4048, n4049, n4050, n4051;
  wire n4052, n4053, n4054, n4055, n4056, n4059, n4060, n4061;
  wire n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069;
  wire n4070, n4071, n4072, n4073, n4074, n4077, n4078, n4079;
  wire n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087;
  wire n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095;
  wire n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105;
  wire n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4115;
  wire n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123;
  wire n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131;
  wire n4132, n4133, n4134, n4135, n4136, n4139, n4140, n4141;
  wire n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149;
  wire n4150, n4151, n4152, n4153, n4156, n4157, n4158, n4159;
  wire n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167;
  wire n4168, n4169, n4170, n4171, n4174, n4175, n4176, n4177;
  wire n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185;
  wire n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193;
  wire n4194, n4195, n4196, n4199, n4200, n4201, n4202, n4203;
  wire n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211;
  wire n4212, n4213, n4214, n4217, n4218, n4219, n4220, n4221;
  wire n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229;
  wire n4230, n4231, n4232, n4233, n4234, n4236, n4237, n4238;
  wire n4239, n4240, n4241, n4242, n4243, n4246, n4247, n4248;
  wire n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256;
  wire n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266;
  wire n4267, n4268, n4269, n4272, n4273, n4274, n4275, n4276;
  wire n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284;
  wire n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292;
  wire n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300;
  wire n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308;
  wire n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316;
  wire n4317, n4318, n4319, n4320, n4321, n4322, n4325, n4326;
  wire n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334;
  wire n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4344;
  wire n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352;
  wire n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360;
  wire n4361, n4364, n4365, n4366, n4367, n4368, n4369, n4370;
  wire n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378;
  wire n4379, n4380, n4383, n4384, n4385, n4386, n4387, n4388;
  wire n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396;
  wire n4397, n4398, n4399, n4400, n4403, n4404, n4405, n4406;
  wire n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414;
  wire n4415, n4416, n4417, n4418, n4419, n4422, n4423, n4424;
  wire n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432;
  wire n4433, n4434, n4435, n4436, n4437, n4438, n4441, n4442;
  wire n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450;
  wire n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4460;
  wire n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468;
  wire n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476;
  wire n4477, n4479, n4480, n4481, n4482, n4483, n4486, n4487;
  wire n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4497;
  wire n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505;
  wire n4506, n4507, n4510, n4511, n4512, n4513, n4514, n4515;
  wire n4516, n4517, n4518, n4519, n4522, n4523, n4524, n4525;
  wire n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533;
  wire n4534, n4537, n4538, n4539, n4540, n4541, n4542, n4543;
  wire n4544, n4545, n4546, n4547, n4548, n4551, n4552, n4553;
  wire n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561;
  wire n4562, n4563, n4564, n4565, n4566, n4567, n4570, n4571;
  wire n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579;
  wire n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587;
  wire n4588, n4589, n4590, n4591, n4592, n4593, n4596, n4597;
  wire n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605;
  wire n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613;
  wire n4614, n4615, n4616, n4617, n4618, n4621, n4622, n4623;
  wire n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631;
  wire n4632, n4633, n4634, n4635, n4636, n4637, n4640, n4641;
  wire n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649;
  wire n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657;
  wire n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665;
  wire n4666, n4667, n4668, n4671, n4672, n4673, n4674, n4675;
  wire n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683;
  wire n4684, n4685, n4686, n4687, n4690, n4691, n4692, n4693;
  wire n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701;
  wire n4702, n4703, n4704, n4705, n4706, n4707, n4709, n4710;
  wire n4711, n4714, n4715, n4716, n4717, n4718, n4719, n4720;
  wire n4721, n4722, n4723, n4724, n4727, n4728, n4729, n4730;
  wire n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738;
  wire n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748;
  wire n4749, n4750, n4753, n4754, n4755, n4756, n4757, n4758;
  wire n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766;
  wire n4767, n4768, n4771, n4772, n4773, n4774, n4775, n4776;
  wire n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784;
  wire n4785, n4786, n4787, n4788, n4789, n4792, n4793, n4794;
  wire n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802;
  wire n4803, n4804, n4805, n4806, n4809, n4810, n4811, n4812;
  wire n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820;
  wire n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828;
  wire n4829, n4830, n4831, n4834, n4835, n4836, n4837, n4838;
  wire n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846;
  wire n4847, n4848, n4851, n4852, n4853, n4854, n4855, n4856;
  wire n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864;
  wire n4865, n4866, n4869, n4870, n4871, n4872, n4873, n4874;
  wire n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882;
  wire n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890;
  wire n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900;
  wire n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908;
  wire n4909, n4910, n4911, n4912, n4913, n4916, n4917, n4918;
  wire n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926;
  wire n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934;
  wire n4935, n4936, n4938, n4939, n4940, n4941, n4944, n4945;
  wire n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953;
  wire n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963;
  wire n4964, n4965, n4966, n4967, n4970, n4971, n4972, n4973;
  wire n4974, n4975, n4976, n4977, n4978, n4979, n4982, n4983;
  wire n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991;
  wire n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001;
  wire n5002, n5003, n5004, n5007, n5008, n5009, n5010, n5011;
  wire n5012, n5013, n5014, n5015, n5016, n5017, n5020, n5021;
  wire n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029;
  wire n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037;
  wire n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045;
  wire n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053;
  wire n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061;
  wire n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069;
  wire n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077;
  wire n5078, n5079, n5080, n5081, n5082, n5083, n5086, n5087;
  wire n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095;
  wire n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5105;
  wire n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113;
  wire n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121;
  wire n5122, n5125, n5126, n5127, n5128, n5129, n5130, n5131;
  wire n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139;
  wire n5140, n5141, n5144, n5145, n5146, n5147, n5148, n5149;
  wire n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157;
  wire n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165;
  wire n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5175;
  wire n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183;
  wire n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191;
  wire n5192, n5194, n5195, n5196, n5199, n5200, n5201, n5202;
  wire n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210;
  wire n5211, n5212, n5213, n5214, n5215, n5218, n5219, n5220;
  wire n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5230;
  wire n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238;
  wire n5239, n5242, n5243, n5244, n5245, n5246, n5247, n5248;
  wire n5249, n5250, n5251, n5254, n5255, n5256, n5257, n5258;
  wire n5259, n5260, n5261, n5262, n5263, n5264, n5267, n5268;
  wire n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276;
  wire n5277, n5278, n5279, n5282, n5283, n5284, n5285, n5286;
  wire n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5296;
  wire n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304;
  wire n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5314;
  wire n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322;
  wire n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330;
  wire n5331, n5332, n5333, n5334, n5335, n5336, n5339, n5340;
  wire n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348;
  wire n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356;
  wire n5357, n5358, n5359, n5360, n5361, n5364, n5365, n5366;
  wire n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374;
  wire n5375, n5376, n5377, n5378, n5379, n5380, n5383, n5384;
  wire n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392;
  wire n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5402;
  wire n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410;
  wire n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418;
  wire n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426;
  wire n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434;
  wire n5435, n5436, n5437, n5438, n5440, n5441, n5442, n5445;
  wire n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453;
  wire n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461;
  wire n5462, n5465, n5466, n5467, n5468, n5469, n5470, n5471;
  wire n5472, n5473, n5474, n5475, n5478, n5479, n5480, n5481;
  wire n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5491;
  wire n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499;
  wire n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509;
  wire n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517;
  wire n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527;
  wire n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535;
  wire n5536, n5537, n5538, n5539, n5540, n5543, n5544, n5545;
  wire n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553;
  wire n5554, n5555, n5556, n5557, n5558, n5559, n5562, n5563;
  wire n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571;
  wire n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579;
  wire n5580, n5581, n5582, n5583, n5584, n5587, n5588, n5589;
  wire n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597;
  wire n5598, n5599, n5600, n5601, n5604, n5605, n5606, n5607;
  wire n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615;
  wire n5616, n5617, n5618, n5619, n5620, n5623, n5624, n5625;
  wire n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633;
  wire n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641;
  wire n5642, n5643, n5644, n5647, n5648, n5649, n5650, n5651;
  wire n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659;
  wire n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667;
  wire n5668, n5671, n5672, n5673, n5674, n5675, n5676, n5677;
  wire n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685;
  wire n5686, n5687, n5688, n5689, n5691, n5692, n5693, n5694;
  wire n5695, n5698, n5699, n5700, n5701, n5702, n5703, n5704;
  wire n5705, n5706, n5707, n5708, n5711, n5712, n5713, n5714;
  wire n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722;
  wire n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732;
  wire n5733, n5736, n5737, n5738, n5739, n5740, n5741, n5742;
  wire n5743, n5744, n5745, n5746, n5749, n5750, n5751, n5752;
  wire n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5762;
  wire n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770;
  wire n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778;
  wire n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786;
  wire n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794;
  wire n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802;
  wire n5803, n5804, n5805, n5806, n5809, n5810, n5811, n5812;
  wire n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820;
  wire n5821, n5822, n5823, n5824, n5825, n5828, n5829, n5830;
  wire n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838;
  wire n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846;
  wire n5847, n5848, n5849, n5850, n5851, n5854, n5855, n5856;
  wire n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864;
  wire n5865, n5866, n5867, n5868, n5869, n5870, n5873, n5874;
  wire n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882;
  wire n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5892;
  wire n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900;
  wire n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908;
  wire n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916;
  wire n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926;
  wire n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934;
  wire n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942;
  wire n5943, n5944, n5945, n5946, n5949, n5950, n5951, n5952;
  wire n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960;
  wire n5961, n5962, n5963, n5964, n5965, n5966, n5968, n5969;
  wire n5970, n5971, n5972, n5973, n5974, n5977, n5978, n5979;
  wire n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5989;
  wire n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997;
  wire n5998, n6001, n6002, n6003, n6004, n6005, n6006, n6007;
  wire n6008, n6009, n6010, n6011, n6014, n6015, n6016, n6017;
  wire n6018, n6019, n6020, n6021, n6022, n6023, n6026, n6027;
  wire n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035;
  wire n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045;
  wire n6046, n6047, n6050, n6051, n6052, n6053, n6054, n6055;
  wire n6056, n6057, n6058, n6059, n6060, n6061, n6064, n6065;
  wire n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073;
  wire n6074, n6075, n6078, n6079, n6080, n6081, n6082, n6083;
  wire n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091;
  wire n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099;
  wire n6100, n6101, n6104, n6105, n6106, n6107, n6108, n6109;
  wire n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117;
  wire n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125;
  wire n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133;
  wire n6134, n6135, n6136, n6137, n6138, n6141, n6142, n6143;
  wire n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151;
  wire n6152, n6153, n6154, n6155, n6156, n6157, n6160, n6161;
  wire n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169;
  wire n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177;
  wire n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185;
  wire n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193;
  wire n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203;
  wire n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6213;
  wire n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221;
  wire n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229;
  wire n6230, n6232, n6233, n6234, n6235, n6238, n6239, n6240;
  wire n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248;
  wire n6249, n6252, n6253, n6254, n6255, n6256, n6257, n6258;
  wire n6259, n6260, n6261, n6262, n6265, n6266, n6267, n6268;
  wire n6269, n6270, n6271, n6272, n6273, n6276, n6277, n6278;
  wire n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286;
  wire n6287, n6290, n6291, n6292, n6293, n6294, n6295, n6296;
  wire n6297, n6298, n6299, n6302, n6303, n6304, n6305, n6306;
  wire n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314;
  wire n6315, n6316, n6317, n6320, n6321, n6322, n6323, n6324;
  wire n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332;
  wire n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6342;
  wire n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350;
  wire n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358;
  wire n6359, n6360, n6361, n6362, n6363, n6364, n6367, n6368;
  wire n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376;
  wire n6377, n6378, n6379, n6380, n6381, n6382, n6385, n6386;
  wire n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394;
  wire n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402;
  wire n6403, n6404, n6405, n6406, n6407, n6410, n6411, n6412;
  wire n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420;
  wire n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428;
  wire n6429, n6430, n6431, n6434, n6435, n6436, n6437, n6438;
  wire n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446;
  wire n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454;
  wire n6455, n6458, n6459, n6460, n6461, n6462, n6463, n6464;
  wire n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472;
  wire n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480;
  wire n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490;
  wire n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498;
  wire n6499, n6500, n6501, n6502, n6504, n6505, n6506, n6509;
  wire n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517;
  wire n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525;
  wire n6526, n6529, n6530, n6531, n6532, n6533, n6534, n6535;
  wire n6536, n6537, n6538, n6539, n6540, n6543, n6544, n6545;
  wire n6546, n6547, n6548, n6549, n6550, n6551, n6554, n6555;
  wire n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563;
  wire n6564, n6567, n6568, n6569, n6570, n6571, n6572, n6573;
  wire n6574, n6575, n6576, n6577, n6580, n6581, n6582, n6583;
  wire n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591;
  wire n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599;
  wire n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607;
  wire n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615;
  wire n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623;
  wire n6624, n6627, n6628, n6629, n6630, n6631, n6632, n6633;
  wire n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641;
  wire n6642, n6643, n6646, n6647, n6648, n6649, n6650, n6651;
  wire n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659;
  wire n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667;
  wire n6668, n6669, n6672, n6673, n6674, n6675, n6676, n6677;
  wire n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685;
  wire n6686, n6687, n6688, n6691, n6692, n6693, n6694, n6695;
  wire n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703;
  wire n6704, n6705, n6706, n6707, n6710, n6711, n6712, n6713;
  wire n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721;
  wire n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729;
  wire n6730, n6731, n6732, n6733, n6734, n6737, n6738, n6739;
  wire n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747;
  wire n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755;
  wire n6756, n6757, n6758, n6759, n6760, n6763, n6764, n6765;
  wire n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773;
  wire n6774, n6775, n6776, n6777, n6778, n6779, n6782, n6783;
  wire n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791;
  wire n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799;
  wire n6800, n6802, n6803, n6804, n6805, n6806, n6809, n6810;
  wire n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6820;
  wire n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828;
  wire n6829, n6832, n6833, n6834, n6835, n6836, n6837, n6838;
  wire n6839, n6840, n6841, n6844, n6845, n6846, n6847, n6848;
  wire n6849, n6850, n6851, n6852, n6853, n6854, n6857, n6858;
  wire n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866;
  wire n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876;
  wire n6877, n6878, n6881, n6882, n6883, n6884, n6885, n6886;
  wire n6887, n6888, n6889, n6890, n6893, n6894, n6895, n6896;
  wire n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904;
  wire n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914;
  wire n6915, n6916, n6917, n6918, n6921, n6922, n6923, n6924;
  wire n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932;
  wire n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940;
  wire n6941, n6942, n6943, n6944, n6947, n6948, n6949, n6950;
  wire n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958;
  wire n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966;
  wire n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974;
  wire n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6984;
  wire n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992;
  wire n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000;
  wire n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010;
  wire n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018;
  wire n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026;
  wire n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034;
  wire n7035, n7036, n7037, n7040, n7041, n7042, n7043, n7044;
  wire n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052;
  wire n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060;
  wire n7061, n7062, n7063, n7066, n7067, n7068, n7069, n7070;
  wire n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078;
  wire n7079, n7080, n7081, n7082, n7083, n7085, n7086, n7087;
  wire n7088, n7089, n7090, n7091, n7094, n7095, n7096, n7097;
  wire n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7107;
  wire n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115;
  wire n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125;
  wire n7126, n7127, n7128, n7129, n7132, n7133, n7134, n7135;
  wire n7136, n7137, n7138, n7139, n7140, n7141, n7144, n7145;
  wire n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153;
  wire n7154, n7155, n7156, n7157, n7158, n7159, n7162, n7163;
  wire n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171;
  wire n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179;
  wire n7180, n7181, n7184, n7185, n7186, n7187, n7188, n7189;
  wire n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197;
  wire n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205;
  wire n7206, n7209, n7210, n7211, n7212, n7213, n7214, n7215;
  wire n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223;
  wire n7224, n7227, n7228, n7229, n7230, n7231, n7232, n7233;
  wire n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241;
  wire n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249;
  wire n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259;
  wire n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267;
  wire n7268, n7269, n7270, n7271, n7272, n7273, n7276, n7277;
  wire n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285;
  wire n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293;
  wire n7294, n7295, n7296, n7297, n7300, n7301, n7302, n7303;
  wire n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311;
  wire n7312, n7313, n7314, n7317, n7318, n7319, n7320, n7321;
  wire n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329;
  wire n7330, n7331, n7332, n7333, n7336, n7337, n7338, n7339;
  wire n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347;
  wire n7348, n7349, n7350, n7351, n7352, n7355, n7356, n7357;
  wire n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365;
  wire n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7374;
  wire n7375, n7376, n7377, n7380, n7381, n7382, n7383, n7384;
  wire n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7394;
  wire n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402;
  wire n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412;
  wire n7413, n7414, n7415, n7418, n7419, n7420, n7421, n7422;
  wire n7423, n7424, n7425, n7426, n7427, n7428, n7431, n7432;
  wire n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440;
  wire n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448;
  wire n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456;
  wire n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464;
  wire n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472;
  wire n7473, n7474, n7475, n7478, n7479, n7480, n7481, n7482;
  wire n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490;
  wire n7491, n7492, n7493, n7494, n7497, n7498, n7499, n7500;
  wire n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508;
  wire n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516;
  wire n7517, n7518, n7519, n7520, n7523, n7524, n7525, n7526;
  wire n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534;
  wire n7535, n7536, n7537, n7538, n7539, n7542, n7543, n7544;
  wire n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552;
  wire n7553, n7554, n7555, n7556, n7557, n7558, n7561, n7562;
  wire n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570;
  wire n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578;
  wire n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7588;
  wire n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596;
  wire n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604;
  wire n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7614;
  wire n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622;
  wire n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630;
  wire n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640;
  wire n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648;
  wire n7649, n7652, n7653, n7654, n7655, n7656, n7657, n7658;
  wire n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666;
  wire n7667, n7668, n7671, n7672, n7673, n7674, n7675, n7676;
  wire n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684;
  wire n7685, n7686, n7687, n7688, n7689, n7690, n7692, n7693;
  wire n7694, n7697, n7698, n7699, n7700, n7701, n7702, n7703;
  wire n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711;
  wire n7712, n7713, n7716, n7717, n7718, n7719, n7720, n7721;
  wire n7722, n7723, n7724, n7725, n7728, n7729, n7730, n7731;
  wire n7732, n7733, n7734, n7735, n7736, n7737, n7740, n7741;
  wire n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749;
  wire n7750, n7751, n7754, n7755, n7756, n7757, n7758, n7759;
  wire n7760, n7761, n7762, n7763, n7766, n7767, n7768, n7769;
  wire n7770, n7771, n7772, n7773, n7774, n7775, n7778, n7779;
  wire n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787;
  wire n7788, n7789, n7792, n7793, n7794, n7795, n7796, n7797;
  wire n7798, n7799, n7800, n7801, n7802, n7803, n7806, n7807;
  wire n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815;
  wire n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823;
  wire n7824, n7825, n7826, n7827, n7828, n7829, n7832, n7833;
  wire n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841;
  wire n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849;
  wire n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857;
  wire n7858, n7859, n7860, n7861, n7864, n7865, n7866, n7867;
  wire n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875;
  wire n7876, n7877, n7878, n7879, n7880, n7883, n7884, n7885;
  wire n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893;
  wire n7894, n7895, n7896, n7897, n7898, n7899, n7902, n7903;
  wire n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911;
  wire n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919;
  wire n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927;
  wire n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935;
  wire n7936, n7939, n7940, n7941, n7942, n7943, n7944, n7945;
  wire n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953;
  wire n7954, n7955, n7958, n7959, n7960, n7961, n7962, n7963;
  wire n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971;
  wire n7972, n7973, n7974, n7977, n7978, n7979, n7980, n7981;
  wire n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989;
  wire n7990, n7991, n7992, n7993, n7994, n7995, n7997, n7998;
  wire n7999, n8000, n8003, n8004, n8005, n8006, n8007, n8008;
  wire n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016;
  wire n8017, n8018, n8019, n8020, n8021, n8024, n8025, n8026;
  wire n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034;
  wire n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044;
  wire n8045, n8046, n8049, n8050, n8051, n8052, n8053, n8054;
  wire n8055, n8056, n8057, n8058, n8061, n8062, n8063, n8064;
  wire n8065, n8066, n8067, n8068, n8069, n8070, n8073, n8074;
  wire n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082;
  wire n8083, n8084, n8085, n8086, n8087, n8088, n8091, n8092;
  wire n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100;
  wire n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108;
  wire n8109, n8110, n8113, n8114, n8115, n8116, n8117, n8118;
  wire n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126;
  wire n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134;
  wire n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8144;
  wire n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152;
  wire n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160;
  wire n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170;
  wire n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178;
  wire n8179, n8182, n8183, n8184, n8185, n8186, n8187, n8188;
  wire n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196;
  wire n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8206;
  wire n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214;
  wire n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222;
  wire n8223, n8224, n8225, n8226, n8227, n8230, n8231, n8232;
  wire n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240;
  wire n8241, n8242, n8243, n8244, n8247, n8248, n8249, n8250;
  wire n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258;
  wire n8259, n8260, n8261, n8262, n8263, n8266, n8267, n8268;
  wire n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276;
  wire n8277, n8278, n8279, n8280, n8281, n8284, n8285, n8286;
  wire n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294;
  wire n8295, n8296, n8297, n8298, n8299, n8300, n8302, n8303;
  wire n8304, n8305, n8306, n8307, n8310, n8311, n8312, n8313;
  wire n8314, n8315, n8316, n8317, n8318, n8321, n8322, n8323;
  wire n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331;
  wire n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341;
  wire n8342, n8343, n8344, n8347, n8348, n8349, n8350, n8351;
  wire n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359;
  wire n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367;
  wire n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375;
  wire n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383;
  wire n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391;
  wire n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401;
  wire n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409;
  wire n8410, n8413, n8414, n8415, n8416, n8417, n8418, n8419;
  wire n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427;
  wire n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435;
  wire n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445;
  wire n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453;
  wire n8454, n8457, n8458, n8459, n8460, n8461, n8462, n8463;
  wire n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471;
  wire n8472, n8473, n8476, n8477, n8478, n8479, n8480, n8481;
  wire n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489;
  wire n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497;
  wire n8498, n8499, n8500, n8503, n8504, n8505, n8506, n8507;
  wire n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515;
  wire n8516, n8517, n8518, n8519, n8522, n8523, n8524, n8525;
  wire n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533;
  wire n8534, n8535, n8536, n8537, n8538, n8539, n8542, n8543;
  wire n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551;
  wire n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8561;
  wire n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569;
  wire n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577;
  wire n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587;
  wire n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595;
  wire n8596, n8597, n8600, n8601, n8602, n8603, n8604, n8605;
  wire n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613;
  wire n8614, n8615, n8616, n8619, n8620, n8621, n8622, n8623;
  wire n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631;
  wire n8632, n8633, n8634, n8635, n8636, n8638, n8639, n8640;
  wire n8641, n8644, n8645, n8646, n8647, n8648, n8649, n8650;
  wire n8651, n8652, n8653, n8656, n8657, n8658, n8659, n8660;
  wire n8661, n8662, n8663, n8664, n8665, n8668, n8669, n8670;
  wire n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678;
  wire n8679, n8682, n8683, n8684, n8685, n8686, n8687, n8688;
  wire n8689, n8690, n8691, n8694, n8695, n8696, n8697, n8698;
  wire n8699, n8700, n8701, n8702, n8703, n8706, n8707, n8708;
  wire n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716;
  wire n8717, n8720, n8721, n8722, n8723, n8724, n8725, n8726;
  wire n8727, n8728, n8729, n8730, n8731, n8734, n8735, n8736;
  wire n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744;
  wire n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752;
  wire n8753, n8754, n8755, n8756, n8757, n8760, n8761, n8762;
  wire n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770;
  wire n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778;
  wire n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786;
  wire n8787, n8788, n8789, n8792, n8793, n8794, n8795, n8796;
  wire n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804;
  wire n8805, n8806, n8807, n8808, n8811, n8812, n8813, n8814;
  wire n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822;
  wire n8823, n8824, n8825, n8826, n8827, n8830, n8831, n8832;
  wire n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840;
  wire n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848;
  wire n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856;
  wire n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864;
  wire n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874;
  wire n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882;
  wire n8883, n8886, n8887, n8888, n8889, n8890, n8891, n8892;
  wire n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900;
  wire n8901, n8902, n8905, n8906, n8907, n8908, n8909, n8910;
  wire n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918;
  wire n8919, n8920, n8921, n8924, n8925, n8926, n8927, n8928;
  wire n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936;
  wire n8937, n8938, n8939, n8940, n8943, n8944, n8945, n8946;
  wire n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954;
  wire n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962;
  wire n8964, n8965, n8966, n8967, n8970, n8971, n8972, n8973;
  wire n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981;
  wire n8982, n8983, n8984, n8985, n8986, n8989, n8990, n8991;
  wire n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999;
  wire n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009;
  wire n9010, n9011, n9012, n9015, n9016, n9017, n9018, n9019;
  wire n9020, n9021, n9022, n9023, n9024, n9027, n9028, n9029;
  wire n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9039;
  wire n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047;
  wire n9048, n9051, n9052, n9053, n9054, n9055, n9056, n9057;
  wire n9058, n9059, n9060, n9063, n9064, n9065, n9066, n9067;
  wire n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075;
  wire n9076, n9077, n9078, n9081, n9082, n9083, n9084, n9085;
  wire n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093;
  wire n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9103;
  wire n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111;
  wire n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119;
  wire n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127;
  wire n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135;
  wire n9136, n9137, n9140, n9141, n9142, n9143, n9144, n9145;
  wire n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153;
  wire n9154, n9155, n9156, n9159, n9160, n9161, n9162, n9163;
  wire n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171;
  wire n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179;
  wire n9180, n9183, n9184, n9185, n9186, n9187, n9188, n9189;
  wire n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197;
  wire n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9207;
  wire n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215;
  wire n9216, n9217, n9218, n9219, n9220, n9221, n9224, n9225;
  wire n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233;
  wire n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9243;
  wire n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251;
  wire n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259;
  wire n9260, n9261, n9262, n9263, n9264, n9265, n9268, n9269;
  wire n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277;
  wire n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9286;
  wire n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294;
  wire n9295, n9298, n9299, n9300, n9301, n9302, n9303, n9304;
  wire n9305, n9306, n9307, n9308, n9311, n9312, n9313, n9314;
  wire n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9324;
  wire n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332;
  wire n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340;
  wire n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348;
  wire n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356;
  wire n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364;
  wire n9365, n9366, n9367, n9368, n9371, n9372, n9373, n9374;
  wire n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382;
  wire n9383, n9384, n9385, n9386, n9387, n9390, n9391, n9392;
  wire n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400;
  wire n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408;
  wire n9409, n9410, n9411, n9412, n9415, n9416, n9417, n9418;
  wire n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426;
  wire n9427, n9428, n9429, n9430, n9431, n9434, n9435, n9436;
  wire n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444;
  wire n9445, n9446, n9447, n9448, n9449, n9450, n9453, n9454;
  wire n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462;
  wire n9463, n9464, n9465, n9466, n9467, n9468, n9471, n9472;
  wire n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480;
  wire n9481, n9482, n9483, n9484, n9485, n9488, n9489, n9490;
  wire n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498;
  wire n9499, n9500, n9501, n9502, n9503, n9504, n9507, n9508;
  wire n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516;
  wire n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524;
  wire n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534;
  wire n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542;
  wire n9543, n9546, n9547, n9548, n9549, n9550, n9551, n9552;
  wire n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560;
  wire n9561, n9562, n9565, n9566, n9567, n9568, n9569, n9570;
  wire n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578;
  wire n9579, n9580, n9581, n9584, n9585, n9586, n9587, n9588;
  wire n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596;
  wire n9597, n9598, n9599, n9600, n9601, n9604, n9605, n9606;
  wire n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614;
  wire n9615, n9616, n9617, n9618, n9619, n9622, n9623, n9624;
  wire n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632;
  wire n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9641;
  wire n9642, n9643, n9644, n9645, n9646, n9649, n9650, n9651;
  wire n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9661;
  wire n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669;
  wire n9670, n9673, n9674, n9675, n9676, n9677, n9678, n9679;
  wire n9680, n9681, n9682, n9683, n9684, n9687, n9688, n9689;
  wire n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9699;
  wire n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707;
  wire n9708, n9711, n9712, n9713, n9714, n9715, n9716, n9717;
  wire n9718, n9719, n9722, n9723, n9724, n9725, n9726, n9727;
  wire n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9737;
  wire n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745;
  wire n9746, n9747, n9748, n9751, n9752, n9753, n9754, n9755;
  wire n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763;
  wire n9764, n9765, n9766, n9767, n9770, n9771, n9772, n9773;
  wire n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781;
  wire n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789;
  wire n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797;
  wire n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805;
  wire n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815;
  wire n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823;
  wire n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831;
  wire n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841;
  wire n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849;
  wire n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857;
  wire n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865;
  wire n9866, n9867, n9868, n9871, n9872, n9873, n9874, n9875;
  wire n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883;
  wire n9884, n9885, n9886, n9887, n9890, n9891, n9892, n9893;
  wire n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901;
  wire n9902, n9903, n9904, n9905, n9906, n9909, n9910, n9911;
  wire n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919;
  wire n9920, n9921, n9922, n9923, n9924, n9925, n9928, n9929;
  wire n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937;
  wire n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9947;
  wire n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955;
  wire n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963;
  wire n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973;
  wire n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981;
  wire n9982, n9983, n9985, n9986, n9987, n9988, n9989, n9992;
  wire n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000;
  wire n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10010;
  wire n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018;
  wire n10019, n10020, n10021, n10022, n10025, n10026, n10027, n10028;
  wire n10029, n10030, n10031, n10032, n10033, n10034, n10037, n10038;
  wire n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046;
  wire n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056;
  wire n10057, n10058, n10061, n10062, n10063, n10064, n10065, n10066;
  wire n10067, n10068, n10069, n10070, n10073, n10074, n10075, n10076;
  wire n10077, n10078, n10079, n10080, n10081, n10082, n10085, n10086;
  wire n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094;
  wire n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104;
  wire n10105, n10106, n10109, n10110, n10111, n10112, n10113, n10114;
  wire n10115, n10116, n10117, n10120, n10121, n10122, n10123, n10124;
  wire n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132;
  wire n10133, n10134, n10135, n10138, n10139, n10140, n10141, n10142;
  wire n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150;
  wire n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158;
  wire n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166;
  wire n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174;
  wire n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182;
  wire n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190;
  wire n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198;
  wire n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206;
  wire n10207, n10208, n10209, n10210, n10213, n10214, n10215, n10216;
  wire n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224;
  wire n10225, n10226, n10227, n10228, n10231, n10232, n10233, n10234;
  wire n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242;
  wire n10243, n10244, n10245, n10248, n10249, n10250, n10251, n10252;
  wire n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260;
  wire n10261, n10262, n10263, n10264, n10267, n10268, n10269, n10270;
  wire n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278;
  wire n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286;
  wire n10287, n10288, n10289, n10292, n10293, n10294, n10295, n10296;
  wire n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304;
  wire n10305, n10306, n10307, n10308, n10311, n10312, n10313, n10314;
  wire n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322;
  wire n10323, n10324, n10325, n10326, n10327, n10329, n10330, n10331;
  wire n10332, n10333, n10336, n10337, n10338, n10339, n10340, n10341;
  wire n10342, n10343, n10344, n10345, n10348, n10349, n10350, n10351;
  wire n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359;
  wire n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369;
  wire n10370, n10371, n10374, n10375, n10376, n10377, n10378, n10379;
  wire n10380, n10381, n10382, n10383, n10386, n10387, n10388, n10389;
  wire n10390, n10391, n10392, n10393, n10394, n10395, n10398, n10399;
  wire n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407;
  wire n10408, n10411, n10412, n10413, n10414, n10415, n10416, n10417;
  wire n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425;
  wire n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433;
  wire n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441;
  wire n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449;
  wire n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457;
  wire n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465;
  wire n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473;
  wire n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483;
  wire n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491;
  wire n10492, n10495, n10496, n10497, n10498, n10499, n10500, n10501;
  wire n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509;
  wire n10510, n10511, n10514, n10515, n10516, n10517, n10518, n10519;
  wire n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527;
  wire n10528, n10529, n10530, n10533, n10534, n10535, n10536, n10537;
  wire n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545;
  wire n10546, n10547, n10548, n10549, n10552, n10553, n10554, n10555;
  wire n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563;
  wire n10564, n10565, n10566, n10567, n10568, n10571, n10572, n10573;
  wire n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581;
  wire n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10591;
  wire n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599;
  wire n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607;
  wire n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617;
  wire n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625;
  wire n10626, n10629, n10630, n10631, n10632, n10633, n10634, n10635;
  wire n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643;
  wire n10644, n10645, n10648, n10649, n10650, n10651, n10652, n10653;
  wire n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661;
  wire n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669;
  wire n10670, n10671, n10672, n10673, n10674, n10675, n10678, n10679;
  wire n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687;
  wire n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695;
  wire n10697, n10698, n10699, n10702, n10703, n10704, n10705, n10706;
  wire n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714;
  wire n10715, n10716, n10717, n10718, n10719, n10720, n10723, n10724;
  wire n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732;
  wire n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742;
  wire n10743, n10744, n10747, n10748, n10749, n10750, n10751, n10752;
  wire n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10762;
  wire n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770;
  wire n10771, n10774, n10775, n10776, n10777, n10778, n10779, n10780;
  wire n10781, n10782, n10783, n10786, n10787, n10788, n10789, n10790;
  wire n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798;
  wire n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808;
  wire n10809, n10810, n10811, n10812, n10815, n10816, n10817, n10818;
  wire n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826;
  wire n10827, n10828, n10829, n10830, n10831, n10834, n10835, n10836;
  wire n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844;
  wire n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852;
  wire n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860;
  wire n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868;
  wire n10869, n10872, n10873, n10874, n10875, n10876, n10877, n10878;
  wire n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886;
  wire n10887, n10890, n10891, n10892, n10893, n10894, n10895, n10896;
  wire n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904;
  wire n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914;
  wire n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922;
  wire n10923, n10926, n10927, n10928, n10929, n10930, n10931, n10932;
  wire n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940;
  wire n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948;
  wire n10949, n10950, n10951, n10952, n10953, n10954, n10957, n10958;
  wire n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966;
  wire n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10976;
  wire n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984;
  wire n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992;
  wire n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002;
  wire n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010;
  wire n11011, n11014, n11015, n11016, n11017, n11018, n11019, n11020;
  wire n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028;
  wire n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036;
  wire n11037, n11040, n11041, n11042, n11043, n11044, n11045, n11046;
  wire n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054;
  wire n11055, n11056, n11057, n11058, n11060, n11061, n11062, n11063;
  wire n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073;
  wire n11074, n11075, n11078, n11079, n11080, n11081, n11082, n11083;
  wire n11084, n11085, n11086, n11087, n11090, n11091, n11092, n11093;
  wire n11094, n11095, n11096, n11097, n11098, n11101, n11102, n11103;
  wire n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111;
  wire n11112, n11113, n11116, n11117, n11118, n11119, n11120, n11121;
  wire n11122, n11123, n11124, n11125, n11126, n11129, n11130, n11131;
  wire n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11141;
  wire n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149;
  wire n11150, n11153, n11154, n11155, n11156, n11157, n11158, n11159;
  wire n11160, n11161, n11162, n11165, n11166, n11167, n11168, n11169;
  wire n11170, n11171, n11172, n11173, n11174, n11177, n11178, n11179;
  wire n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187;
  wire n11188, n11189, n11190, n11191, n11192, n11195, n11196, n11197;
  wire n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205;
  wire n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213;
  wire n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223;
  wire n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231;
  wire n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239;
  wire n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247;
  wire n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255;
  wire n11256, n11259, n11260, n11261, n11262, n11263, n11264, n11265;
  wire n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273;
  wire n11274, n11275, n11278, n11279, n11280, n11281, n11282, n11283;
  wire n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291;
  wire n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11301;
  wire n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309;
  wire n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11319;
  wire n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327;
  wire n11328, n11329, n11330, n11331, n11332, n11333, n11336, n11337;
  wire n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345;
  wire n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11355;
  wire n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363;
  wire n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371;
  wire n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379;
  wire n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387;
  wire n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395;
  wire n11396, n11397, n11398, n11399, n11400, n11401, n11404, n11405;
  wire n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413;
  wire n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421;
  wire n11422, n11423, n11425, n11426, n11427, n11430, n11431, n11432;
  wire n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440;
  wire n11441, n11442, n11443, n11444, n11445, n11446, n11449, n11450;
  wire n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458;
  wire n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468;
  wire n11469, n11470, n11473, n11474, n11475, n11476, n11477, n11478;
  wire n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486;
  wire n11487, n11490, n11491, n11492, n11493, n11494, n11495, n11496;
  wire n11497, n11498, n11499, n11500, n11503, n11504, n11505, n11506;
  wire n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11516;
  wire n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524;
  wire n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532;
  wire n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540;
  wire n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548;
  wire n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556;
  wire n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564;
  wire n11565, n11566, n11569, n11570, n11571, n11572, n11573, n11574;
  wire n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582;
  wire n11583, n11584, n11585, n11588, n11589, n11590, n11591, n11592;
  wire n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600;
  wire n11601, n11602, n11603, n11604, n11607, n11608, n11609, n11610;
  wire n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618;
  wire n11619, n11620, n11621, n11622, n11623, n11626, n11627, n11628;
  wire n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636;
  wire n11637, n11638, n11639, n11640, n11641, n11642, n11645, n11646;
  wire n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654;
  wire n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11664;
  wire n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672;
  wire n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11682;
  wire n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690;
  wire n11691, n11692, n11693, n11694, n11695, n11696, n11699, n11700;
  wire n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708;
  wire n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716;
  wire n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726;
  wire n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734;
  wire n11735, n11738, n11739, n11740, n11741, n11742, n11743, n11744;
  wire n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752;
  wire n11753, n11754, n11757, n11758, n11759, n11760, n11761, n11762;
  wire n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770;
  wire n11771, n11772, n11773, n11776, n11777, n11778, n11779, n11780;
  wire n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788;
  wire n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796;
  wire n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804;
  wire n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812;
  wire n11814, n11815, n11816, n11817, n11818, n11819, n11822, n11823;
  wire n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831;
  wire n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841;
  wire n11842, n11843, n11844, n11847, n11848, n11849, n11850, n11851;
  wire n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859;
  wire n11860, n11863, n11864, n11865, n11866, n11867, n11868, n11869;
  wire n11870, n11871, n11874, n11875, n11876, n11877, n11878, n11879;
  wire n11880, n11881, n11882, n11883, n11886, n11887, n11888, n11889;
  wire n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897;
  wire n11898, n11901, n11902, n11903, n11904, n11905, n11906, n11907;
  wire n11908, n11909, n11910, n11911, n11912, n11915, n11916, n11917;
  wire n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925;
  wire n11926, n11927, n11928, n11929, n11930, n11931, n11934, n11935;
  wire n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943;
  wire n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951;
  wire n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959;
  wire n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967;
  wire n11968, n11969, n11972, n11973, n11974, n11975, n11976, n11977;
  wire n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985;
  wire n11986, n11987, n11990, n11991, n11992, n11993, n11994, n11995;
  wire n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003;
  wire n12004, n12007, n12008, n12009, n12010, n12011, n12012, n12013;
  wire n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021;
  wire n12022, n12023, n12026, n12027, n12028, n12029, n12030, n12031;
  wire n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039;
  wire n12040, n12041, n12042, n12045, n12046, n12047, n12048, n12049;
  wire n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057;
  wire n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065;
  wire n12066, n12067, n12070, n12071, n12072, n12073, n12074, n12075;
  wire n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083;
  wire n12084, n12085, n12086, n12089, n12090, n12091, n12092, n12093;
  wire n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101;
  wire n12102, n12103, n12104, n12105, n12108, n12109, n12110, n12111;
  wire n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119;
  wire n12120, n12121, n12122, n12123, n12126, n12127, n12128, n12129;
  wire n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137;
  wire n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145;
  wire n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153;
  wire n12154, n12155, n12158, n12159, n12160, n12161, n12162, n12163;
  wire n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12173;
  wire n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181;
  wire n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189;
  wire n12190, n12191, n12192, n12193, n12194, n12195, n12197, n12198;
  wire n12199, n12200, n12201, n12202, n12205, n12206, n12207, n12208;
  wire n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216;
  wire n12217, n12218, n12219, n12220, n12223, n12224, n12225, n12226;
  wire n12227, n12228, n12229, n12230, n12231, n12232, n12235, n12236;
  wire n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244;
  wire n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254;
  wire n12255, n12256, n12259, n12260, n12261, n12262, n12263, n12264;
  wire n12265, n12266, n12267, n12268, n12269, n12272, n12273, n12274;
  wire n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282;
  wire n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292;
  wire n12293, n12294, n12295, n12298, n12299, n12300, n12301, n12302;
  wire n12303, n12304, n12305, n12306, n12307, n12310, n12311, n12312;
  wire n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12322;
  wire n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330;
  wire n12331, n12334, n12335, n12336, n12337, n12338, n12339, n12340;
  wire n12341, n12342, n12343, n12346, n12347, n12348, n12349, n12350;
  wire n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358;
  wire n12359, n12360, n12361, n12364, n12365, n12366, n12367, n12368;
  wire n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376;
  wire n12377, n12378, n12379, n12380, n12381, n12382, n12385, n12386;
  wire n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394;
  wire n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402;
  wire n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410;
  wire n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418;
  wire n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12428;
  wire n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436;
  wire n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444;
  wire n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454;
  wire n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462;
  wire n12463, n12466, n12467, n12468, n12469, n12470, n12471, n12472;
  wire n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480;
  wire n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12490;
  wire n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498;
  wire n12499, n12500, n12501, n12502, n12503, n12504, n12507, n12508;
  wire n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516;
  wire n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12526;
  wire n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534;
  wire n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542;
  wire n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550;
  wire n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558;
  wire n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566;
  wire n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574;
  wire n12575, n12576, n12577, n12578, n12580, n12581, n12582, n12585;
  wire n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593;
  wire n12594, n12597, n12598, n12599, n12600, n12601, n12602, n12603;
  wire n12604, n12605, n12606, n12609, n12610, n12611, n12612, n12613;
  wire n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621;
  wire n12622, n12623, n12624, n12627, n12628, n12629, n12630, n12631;
  wire n12632, n12633, n12634, n12635, n12636, n12637, n12640, n12641;
  wire n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649;
  wire n12650, n12653, n12654, n12655, n12656, n12657, n12658, n12659;
  wire n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667;
  wire n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675;
  wire n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683;
  wire n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691;
  wire n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699;
  wire n12700, n12701, n12702, n12703, n12706, n12707, n12708, n12709;
  wire n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717;
  wire n12718, n12719, n12720, n12721, n12722, n12725, n12726, n12727;
  wire n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735;
  wire n12736, n12737, n12738, n12739, n12740, n12741, n12744, n12745;
  wire n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753;
  wire n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12763;
  wire n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771;
  wire n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779;
  wire n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789;
  wire n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797;
  wire n12798, n12801, n12802, n12803, n12804, n12805, n12806, n12807;
  wire n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815;
  wire n12816, n12817, n12820, n12821, n12822, n12823, n12824, n12825;
  wire n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833;
  wire n12834, n12835, n12838, n12839, n12840, n12841, n12842, n12843;
  wire n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851;
  wire n12852, n12855, n12856, n12857, n12858, n12859, n12860, n12861;
  wire n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869;
  wire n12870, n12871, n12874, n12875, n12876, n12877, n12878, n12879;
  wire n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887;
  wire n12888, n12889, n12890, n12893, n12894, n12895, n12896, n12897;
  wire n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905;
  wire n12906, n12907, n12908, n12909, n12912, n12913, n12914, n12915;
  wire n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923;
  wire n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931;
  wire n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939;
  wire n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12949;
  wire n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957;
  wire n12958, n12959, n12960, n12963, n12964, n12965, n12966, n12967;
  wire n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975;
  wire n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983;
  wire n12984, n12985, n12986, n12988, n12989, n12990, n12991, n12992;
  wire n12993, n12994, n12997, n12998, n12999, n13000, n13001, n13002;
  wire n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010;
  wire n13011, n13014, n13015, n13016, n13017, n13018, n13019, n13020;
  wire n13021, n13022, n13025, n13026, n13027, n13028, n13029, n13030;
  wire n13031, n13032, n13033, n13034, n13037, n13038, n13039, n13040;
  wire n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048;
  wire n13049, n13052, n13053, n13054, n13055, n13056, n13057, n13058;
  wire n13059, n13060, n13061, n13062, n13063, n13066, n13067, n13068;
  wire n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076;
  wire n13077, n13078, n13079, n13080, n13081, n13082, n13085, n13086;
  wire n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094;
  wire n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102;
  wire n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110;
  wire n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118;
  wire n13119, n13120, n13123, n13124, n13125, n13126, n13127, n13128;
  wire n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136;
  wire n13137, n13138, n13141, n13142, n13143, n13144, n13145, n13146;
  wire n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154;
  wire n13155, n13158, n13159, n13160, n13161, n13162, n13163, n13164;
  wire n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172;
  wire n13173, n13174, n13177, n13178, n13179, n13180, n13181, n13182;
  wire n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190;
  wire n13191, n13192, n13193, n13196, n13197, n13198, n13199, n13200;
  wire n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208;
  wire n13209, n13210, n13211, n13212, n13215, n13216, n13217, n13218;
  wire n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226;
  wire n13227, n13228, n13229, n13230, n13231, n13234, n13235, n13236;
  wire n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244;
  wire n13245, n13246, n13247, n13248, n13249, n13250, n13253, n13254;
  wire n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262;
  wire n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13272;
  wire n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280;
  wire n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13290;
  wire n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298;
  wire n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306;
  wire n13307, n13308, n13309, n13310, n13311, n13314, n13315, n13316;
  wire n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324;
  wire n13325, n13326, n13327, n13328, n13331, n13332, n13333, n13334;
  wire n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342;
  wire n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352;
  wire n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360;
  wire n13361, n13364, n13365, n13366, n13367, n13368, n13369, n13370;
  wire n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378;
  wire n13379, n13380, n13381, n13382, n13383, n13384, n13386, n13387;
  wire n13388, n13389, n13390, n13393, n13394, n13395, n13396, n13397;
  wire n13398, n13399, n13400, n13401, n13402, n13405, n13406, n13407;
  wire n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415;
  wire n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425;
  wire n13426, n13429, n13430, n13431, n13432, n13433, n13434, n13435;
  wire n13436, n13437, n13438, n13439, n13442, n13443, n13444, n13445;
  wire n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13455;
  wire n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463;
  wire n13464, n13467, n13468, n13469, n13470, n13471, n13472, n13473;
  wire n13474, n13475, n13476, n13477, n13480, n13481, n13482, n13483;
  wire n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491;
  wire n13492, n13493, n13494, n13495, n13496, n13499, n13500, n13501;
  wire n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509;
  wire n13510, n13511, n13514, n13515, n13516, n13517, n13518, n13519;
  wire n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527;
  wire n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535;
  wire n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545;
  wire n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553;
  wire n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13563;
  wire n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571;
  wire n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579;
  wire n13580, n13581, n13582, n13583, n13586, n13587, n13588, n13589;
  wire n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597;
  wire n13598, n13599, n13600, n13601, n13602, n13605, n13606, n13607;
  wire n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615;
  wire n13616, n13617, n13618, n13619, n13620, n13621, n13624, n13625;
  wire n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633;
  wire n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641;
  wire n13642, n13643, n13644, n13645, n13646, n13649, n13650, n13651;
  wire n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659;
  wire n13660, n13661, n13662, n13663, n13666, n13667, n13668, n13669;
  wire n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677;
  wire n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685;
  wire n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693;
  wire n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701;
  wire n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709;
  wire n13710, n13713, n13714, n13715, n13716, n13717, n13718, n13719;
  wire n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727;
  wire n13728, n13729, n13732, n13733, n13734, n13735, n13736, n13737;
  wire n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13747;
  wire n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755;
  wire n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13765;
  wire n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773;
  wire n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781;
  wire n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789;
  wire n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798;
  wire n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806;
  wire n13807, n13808, n13809, n13810, n13811, n13812, n13815, n13816;
  wire n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824;
  wire n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834;
  wire n13835, n13836, n13839, n13840, n13841, n13842, n13843, n13844;
  wire n13845, n13846, n13847, n13848, n13851, n13852, n13853, n13854;
  wire n13855, n13856, n13857, n13858, n13859, n13860, n13863, n13864;
  wire n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13874;
  wire n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882;
  wire n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892;
  wire n13893, n13896, n13897, n13898, n13899, n13900, n13901, n13902;
  wire n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13912;
  wire n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920;
  wire n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928;
  wire n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938;
  wire n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946;
  wire n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954;
  wire n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964;
  wire n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972;
  wire n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980;
  wire n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990;
  wire n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998;
  wire n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006;
  wire n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016;
  wire n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024;
  wire n14025, n14028, n14029, n14030, n14031, n14032, n14033, n14034;
  wire n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042;
  wire n14043, n14044, n14047, n14048, n14049, n14050, n14051, n14052;
  wire n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060;
  wire n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068;
  wire n14069, n14070, n14071, n14074, n14075, n14076, n14077, n14078;
  wire n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086;
  wire n14087, n14088, n14089, n14090, n14093, n14094, n14095, n14096;
  wire n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104;
  wire n14105, n14106, n14107, n14108, n14109, n14110, n14113, n14114;
  wire n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122;
  wire n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130;
  wire n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138;
  wire n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146;
  wire n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154;
  wire n14155, n14158, n14159, n14160, n14161, n14162, n14163, n14164;
  wire n14165, n14166, n14167, n14168, n14169, n14170, n14173, n14174;
  wire n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182;
  wire n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190;
  wire n14191, n14192, n14194, n14195, n14196, n14199, n14200, n14201;
  wire n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209;
  wire n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219;
  wire n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14229;
  wire n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237;
  wire n14238, n14239, n14240, n14241, n14242, n14245, n14246, n14247;
  wire n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255;
  wire n14256, n14257, n14258, n14259, n14260, n14261, n14264, n14265;
  wire n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273;
  wire n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14283;
  wire n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291;
  wire n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299;
  wire n14300, n14301, n14302, n14303, n14304, n14307, n14308, n14309;
  wire n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317;
  wire n14318, n14319, n14320, n14321, n14324, n14325, n14326, n14327;
  wire n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335;
  wire n14336, n14337, n14338, n14339, n14342, n14343, n14344, n14345;
  wire n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353;
  wire n14354, n14355, n14356, n14359, n14360, n14361, n14362, n14363;
  wire n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371;
  wire n14372, n14373, n14374, n14375, n14378, n14379, n14380, n14381;
  wire n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389;
  wire n14390, n14391, n14392, n14393, n14394, n14397, n14398, n14399;
  wire n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407;
  wire n14408, n14409, n14410, n14411, n14412, n14413, n14416, n14417;
  wire n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425;
  wire n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14435;
  wire n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443;
  wire n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451;
  wire n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461;
  wire n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469;
  wire n14470, n14473, n14474, n14475, n14476, n14477, n14478, n14479;
  wire n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487;
  wire n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495;
  wire n14496, n14497, n14498, n14501, n14502, n14503, n14504, n14505;
  wire n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513;
  wire n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521;
  wire n14522, n14523, n14526, n14527, n14528, n14529, n14530, n14531;
  wire n14532, n14533, n14534, n14535, n14536, n14537, n14540, n14541;
  wire n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549;
  wire n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14559;
  wire n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567;
  wire n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575;
  wire n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583;
  wire n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14592;
  wire n14593, n14594, n14595, n14598, n14599, n14600, n14601, n14602;
  wire n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610;
  wire n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620;
  wire n14621, n14622, n14623, n14624, n14625, n14628, n14629, n14630;
  wire n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638;
  wire n14639, n14640, n14643, n14644, n14645, n14646, n14647, n14648;
  wire n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14658;
  wire n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666;
  wire n14667, n14668, n14669, n14672, n14673, n14674, n14675, n14676;
  wire n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684;
  wire n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692;
  wire n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14702;
  wire n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710;
  wire n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720;
  wire n14721, n14724, n14725, n14726, n14727, n14728, n14729, n14730;
  wire n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738;
  wire n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746;
  wire n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754;
  wire n14755, n14756, n14757, n14760, n14761, n14762, n14763, n14764;
  wire n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772;
  wire n14773, n14774, n14775, n14778, n14779, n14780, n14781, n14782;
  wire n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790;
  wire n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798;
  wire n14799, n14800, n14801, n14804, n14805, n14806, n14807, n14808;
  wire n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816;
  wire n14817, n14818, n14819, n14820, n14823, n14824, n14825, n14826;
  wire n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834;
  wire n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842;
  wire n14843, n14844, n14845, n14846, n14847, n14850, n14851, n14852;
  wire n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860;
  wire n14861, n14862, n14863, n14864, n14865, n14866, n14869, n14870;
  wire n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878;
  wire n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886;
  wire n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894;
  wire n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902;
  wire n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910;
  wire n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918;
  wire n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926;
  wire n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934;
  wire n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942;
  wire n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950;
  wire n14951, n14954, n14955, n14956, n14957, n14958, n14959, n14960;
  wire n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968;
  wire n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976;
  wire n14977, n14978, n14979, n14981, n14982, n14983, n14984, n14985;
  wire n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995;
  wire n14996, n14997, n14998, n14999, n15000, n15003, n15004, n15005;
  wire n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013;
  wire n15014, n15015, n15016, n15019, n15020, n15021, n15022, n15023;
  wire n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031;
  wire n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039;
  wire n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15049;
  wire n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057;
  wire n15058, n15061, n15062, n15063, n15064, n15065, n15066, n15067;
  wire n15068, n15069, n15072, n15073, n15074, n15075, n15076, n15077;
  wire n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085;
  wire n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093;
  wire n15094, n15095, n15098, n15099, n15100, n15101, n15102, n15103;
  wire n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111;
  wire n15112, n15113, n15114, n15117, n15118, n15119, n15120, n15121;
  wire n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129;
  wire n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137;
  wire n15138, n15139, n15140, n15141, n15144, n15145, n15146, n15147;
  wire n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155;
  wire n15156, n15157, n15158, n15159, n15160, n15163, n15164, n15165;
  wire n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173;
  wire n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15183;
  wire n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191;
  wire n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199;
  wire n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209;
  wire n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217;
  wire n15218, n15221, n15222, n15223, n15224, n15225, n15226, n15227;
  wire n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235;
  wire n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243;
  wire n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251;
  wire n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259;
  wire n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267;
  wire n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277;
  wire n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285;
  wire n15286, n15287, n15288, n15289, n15290, n15293, n15294, n15295;
  wire n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303;
  wire n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311;
  wire n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319;
  wire n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327;
  wire n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335;
  wire n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343;
  wire n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351;
  wire n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359;
  wire n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367;
  wire n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375;
  wire n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384;
  wire n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392;
  wire n15393, n15396, n15397, n15398, n15399, n15400, n15401, n15402;
  wire n15403, n15404, n15405, n15406, n15407, n15408, n15411, n15412;
  wire n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420;
  wire n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428;
  wire n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436;
  wire n15437, n15438, n15439, n15440, n15443, n15444, n15445, n15446;
  wire n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454;
  wire n15455, n15456, n15457, n15460, n15461, n15462, n15463, n15464;
  wire n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472;
  wire n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482;
  wire n15483, n15484, n15485, n15486, n15487, n15490, n15491, n15492;
  wire n15493, n15494, n15495, n15496, n15497, n15498, n15501, n15502;
  wire n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15512;
  wire n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520;
  wire n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530;
  wire n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538;
  wire n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546;
  wire n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556;
  wire n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564;
  wire n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572;
  wire n15573, n15576, n15577, n15578, n15579, n15580, n15581, n15582;
  wire n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590;
  wire n15591, n15592, n15595, n15596, n15597, n15598, n15599, n15600;
  wire n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608;
  wire n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616;
  wire n15617, n15618, n15621, n15622, n15623, n15624, n15625, n15626;
  wire n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634;
  wire n15635, n15636, n15637, n15640, n15641, n15642, n15643, n15644;
  wire n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652;
  wire n15653, n15654, n15655, n15656, n15659, n15660, n15661, n15662;
  wire n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670;
  wire n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678;
  wire n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686;
  wire n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694;
  wire n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702;
  wire n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710;
  wire n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718;
  wire n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726;
  wire n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734;
  wire n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742;
  wire n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750;
  wire n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758;
  wire n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766;
  wire n15768, n15769, n15770, n15771, n15772, n15773, n15776, n15777;
  wire n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785;
  wire n15786, n15787, n15788, n15791, n15792, n15793, n15794, n15795;
  wire n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803;
  wire n15804, n15807, n15808, n15809, n15810, n15811, n15812, n15813;
  wire n15814, n15815, n15816, n15817, n15818, n15819, n15822, n15823;
  wire n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831;
  wire n15832, n15833, n15834, n15835, n15838, n15839, n15840, n15841;
  wire n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849;
  wire n15850, n15853, n15854, n15855, n15856, n15857, n15858, n15859;
  wire n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867;
  wire n15868, n15869, n15870, n15871, n15874, n15875, n15876, n15877;
  wire n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885;
  wire n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893;
  wire n15894, n15895, n15898, n15899, n15900, n15901, n15902, n15903;
  wire n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911;
  wire n15912, n15913, n15914, n15915, n15916, n15917, n15920, n15921;
  wire n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929;
  wire n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15939;
  wire n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947;
  wire n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955;
  wire n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965;
  wire n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973;
  wire n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983;
  wire n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15993;
  wire n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001;
  wire n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009;
  wire n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019;
  wire n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027;
  wire n16028, n16031, n16032, n16033, n16034, n16035, n16036, n16037;
  wire n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045;
  wire n16046, n16049, n16050, n16051, n16052, n16053, n16054, n16055;
  wire n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063;
  wire n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073;
  wire n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081;
  wire n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089;
  wire n16090, n16091, n16094, n16095, n16096, n16097, n16098, n16099;
  wire n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107;
  wire n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115;
  wire n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125;
  wire n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133;
  wire n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141;
  wire n16142, n16143, n16144, n16146, n16147, n16148, n16149, n16150;
  wire n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158;
  wire n16159, n16160, n16161, n16164, n16165, n16166, n16167, n16168;
  wire n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176;
  wire n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184;
  wire n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16194;
  wire n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202;
  wire n16203, n16204, n16205, n16206, n16209, n16210, n16211, n16212;
  wire n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220;
  wire n16221, n16224, n16225, n16226, n16227, n16228, n16229, n16230;
  wire n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238;
  wire n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246;
  wire n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16256;
  wire n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264;
  wire n16265, n16266, n16267, n16268, n16269, n16272, n16273, n16274;
  wire n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282;
  wire n16283, n16284, n16287, n16288, n16289, n16290, n16291, n16292;
  wire n16293, n16294, n16295, n16296, n16297, n16300, n16301, n16302;
  wire n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310;
  wire n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318;
  wire n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326;
  wire n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334;
  wire n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344;
  wire n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352;
  wire n16353, n16356, n16357, n16358, n16359, n16360, n16361, n16362;
  wire n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370;
  wire n16371, n16372, n16375, n16376, n16377, n16378, n16379, n16380;
  wire n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388;
  wire n16389, n16390, n16391, n16394, n16395, n16396, n16397, n16398;
  wire n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406;
  wire n16407, n16408, n16409, n16410, n16411, n16414, n16415, n16416;
  wire n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424;
  wire n16425, n16426, n16427, n16428, n16429, n16430, n16433, n16434;
  wire n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442;
  wire n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16452;
  wire n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460;
  wire n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468;
  wire n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476;
  wire n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484;
  wire n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492;
  wire n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500;
  wire n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508;
  wire n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516;
  wire n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525;
  wire n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533;
  wire n16534, n16537, n16538, n16539, n16540, n16541, n16542, n16543;
  wire n16544, n16545, n16546, n16547, n16548, n16549, n16552, n16553;
  wire n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561;
  wire n16562, n16563, n16564, n16567, n16568, n16569, n16570, n16571;
  wire n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579;
  wire n16580, n16581, n16584, n16585, n16586, n16587, n16588, n16589;
  wire n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16599;
  wire n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607;
  wire n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617;
  wire n16618, n16619, n16622, n16623, n16624, n16625, n16626, n16627;
  wire n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635;
  wire n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643;
  wire n16644, n16647, n16648, n16649, n16650, n16651, n16652, n16653;
  wire n16654, n16655, n16656, n16657, n16658, n16661, n16662, n16663;
  wire n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671;
  wire n16672, n16673, n16674, n16675, n16678, n16679, n16680, n16681;
  wire n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689;
  wire n16690, n16691, n16692, n16693, n16694, n16697, n16698, n16699;
  wire n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707;
  wire n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715;
  wire n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723;
  wire n16724, n16725, n16726, n16727, n16730, n16731, n16732, n16733;
  wire n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741;
  wire n16742, n16743, n16744, n16745, n16746, n16749, n16750, n16751;
  wire n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759;
  wire n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767;
  wire n16768, n16769, n16770, n16771, n16772, n16775, n16776, n16777;
  wire n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785;
  wire n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793;
  wire n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801;
  wire n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809;
  wire n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817;
  wire n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825;
  wire n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833;
  wire n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841;
  wire n16842, n16843, n16846, n16847, n16848, n16849, n16850, n16851;
  wire n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859;
  wire n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867;
  wire n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875;
  wire n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883;
  wire n16884, n16885, n16886, n16887, n16888, n16889, n16891, n16892;
  wire n16893, n16894, n16895, n16896, n16899, n16900, n16901, n16902;
  wire n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910;
  wire n16911, n16912, n16913, n16916, n16917, n16918, n16919, n16920;
  wire n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16930;
  wire n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938;
  wire n16939, n16940, n16941, n16942, n16943, n16946, n16947, n16948;
  wire n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956;
  wire n16957, n16958, n16961, n16962, n16963, n16964, n16965, n16966;
  wire n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974;
  wire n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984;
  wire n16985, n16986, n16987, n16988, n16989, n16990, n16993, n16994;
  wire n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002;
  wire n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17012;
  wire n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020;
  wire n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030;
  wire n17031, n17032, n17033, n17036, n17037, n17038, n17039, n17040;
  wire n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048;
  wire n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056;
  wire n17057, n17058, n17059, n17062, n17063, n17064, n17065, n17066;
  wire n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074;
  wire n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082;
  wire n17083, n17084, n17087, n17088, n17089, n17090, n17091, n17092;
  wire n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100;
  wire n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108;
  wire n17109, n17110, n17111, n17114, n17115, n17116, n17117, n17118;
  wire n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126;
  wire n17127, n17128, n17129, n17130, n17133, n17134, n17135, n17136;
  wire n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144;
  wire n17145, n17146, n17147, n17148, n17149, n17152, n17153, n17154;
  wire n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162;
  wire n17163, n17164, n17165, n17166, n17167, n17170, n17171, n17172;
  wire n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180;
  wire n17181, n17182, n17183, n17184, n17187, n17188, n17189, n17190;
  wire n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198;
  wire n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206;
  wire n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214;
  wire n17215, n17218, n17219, n17220, n17221, n17222, n17223, n17224;
  wire n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232;
  wire n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240;
  wire n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248;
  wire n17249, n17250, n17251, n17252, n17253, n17255, n17256, n17257;
  wire n17258, n17259, n17260, n17263, n17264, n17265, n17266, n17267;
  wire n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275;
  wire n17276, n17279, n17280, n17281, n17282, n17283, n17284, n17285;
  wire n17286, n17287, n17288, n17289, n17290, n17291, n17294, n17295;
  wire n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303;
  wire n17304, n17305, n17306, n17309, n17310, n17311, n17312, n17313;
  wire n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321;
  wire n17322, n17323, n17326, n17327, n17328, n17329, n17330, n17331;
  wire n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17341;
  wire n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349;
  wire n17350, n17353, n17354, n17355, n17356, n17357, n17358, n17359;
  wire n17360, n17361, n17362, n17363, n17366, n17367, n17368, n17369;
  wire n17370, n17371, n17372, n17373, n17374, n17377, n17378, n17379;
  wire n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387;
  wire n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395;
  wire n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403;
  wire n17404, n17407, n17408, n17409, n17410, n17411, n17412, n17413;
  wire n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421;
  wire n17422, n17423, n17426, n17427, n17428, n17429, n17430, n17431;
  wire n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439;
  wire n17440, n17441, n17442, n17445, n17446, n17447, n17448, n17449;
  wire n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457;
  wire n17458, n17459, n17460, n17461, n17464, n17465, n17466, n17467;
  wire n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475;
  wire n17476, n17477, n17478, n17479, n17480, n17483, n17484, n17485;
  wire n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493;
  wire n17494, n17495, n17496, n17497, n17498, n17499, n17502, n17503;
  wire n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511;
  wire n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519;
  wire n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527;
  wire n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535;
  wire n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543;
  wire n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551;
  wire n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559;
  wire n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567;
  wire n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575;
  wire n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583;
  wire n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591;
  wire n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599;
  wire n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607;
  wire n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615;
  wire n17616, n17617, n17618, n17620, n17621, n17622, n17623, n17624;
  wire n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632;
  wire n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640;
  wire n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648;
  wire n17649, n17650, n17651, n17654, n17655, n17656, n17657, n17658;
  wire n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666;
  wire n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676;
  wire n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684;
  wire n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692;
  wire n17693, n17694, n17695, n17696, n17697, n17700, n17701, n17702;
  wire n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710;
  wire n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718;
  wire n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726;
  wire n17727, n17730, n17731, n17732, n17733, n17734, n17735, n17736;
  wire n17737, n17738, n17739, n17742, n17743, n17744, n17745, n17746;
  wire n17747, n17748, n17749, n17750, n17751, n17754, n17755, n17756;
  wire n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17766;
  wire n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774;
  wire n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782;
  wire n17783, n17784, n17785, n17786, n17787, n17790, n17791, n17792;
  wire n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800;
  wire n17801, n17802, n17805, n17806, n17807, n17808, n17809, n17810;
  wire n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818;
  wire n17819, n17820, n17821, n17824, n17825, n17826, n17827, n17828;
  wire n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836;
  wire n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844;
  wire n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852;
  wire n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862;
  wire n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870;
  wire n17871, n17874, n17875, n17876, n17877, n17878, n17879, n17880;
  wire n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888;
  wire n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896;
  wire n17897, n17900, n17901, n17902, n17903, n17904, n17905, n17906;
  wire n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914;
  wire n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922;
  wire n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930;
  wire n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938;
  wire n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946;
  wire n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954;
  wire n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962;
  wire n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17971;
  wire n17972, n17973, n17974, n17975, n17976, n17977, n17980, n17981;
  wire n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989;
  wire n17990, n17991, n17992, n17993, n17996, n17997, n17998, n17999;
  wire n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007;
  wire n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017;
  wire n18018, n18019, n18020, n18021, n18022, n18023, n18026, n18027;
  wire n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035;
  wire n18036, n18037, n18038, n18041, n18042, n18043, n18044, n18045;
  wire n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053;
  wire n18054, n18057, n18058, n18059, n18060, n18061, n18062, n18063;
  wire n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071;
  wire n18072, n18073, n18074, n18077, n18078, n18079, n18080, n18081;
  wire n18082, n18083, n18084, n18085, n18086, n18089, n18090, n18091;
  wire n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099;
  wire n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107;
  wire n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18117;
  wire n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125;
  wire n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133;
  wire n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143;
  wire n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151;
  wire n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159;
  wire n18160, n18163, n18164, n18165, n18166, n18167, n18168, n18169;
  wire n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177;
  wire n18178, n18179, n18182, n18183, n18184, n18185, n18186, n18187;
  wire n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195;
  wire n18196, n18197, n18198, n18201, n18202, n18203, n18204, n18205;
  wire n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213;
  wire n18214, n18215, n18216, n18219, n18220, n18221, n18222, n18223;
  wire n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231;
  wire n18232, n18233, n18236, n18237, n18238, n18239, n18240, n18241;
  wire n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249;
  wire n18250, n18251, n18254, n18255, n18256, n18257, n18258, n18259;
  wire n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267;
  wire n18268, n18269, n18272, n18273, n18274, n18275, n18276, n18277;
  wire n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285;
  wire n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293;
  wire n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301;
  wire n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309;
  wire n18310, n18311, n18312, n18313, n18314, n18315, n18317, n18318;
  wire n18319, n18320, n18321, n18322, n18325, n18326, n18327, n18328;
  wire n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336;
  wire n18337, n18338, n18341, n18342, n18343, n18344, n18345, n18346;
  wire n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354;
  wire n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364;
  wire n18365, n18366, n18367, n18368, n18369, n18370, n18373, n18374;
  wire n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382;
  wire n18383, n18386, n18387, n18388, n18389, n18390, n18391, n18392;
  wire n18393, n18394, n18395, n18398, n18399, n18400, n18401, n18402;
  wire n18403, n18404, n18405, n18406, n18407, n18408, n18411, n18412;
  wire n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18422;
  wire n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430;
  wire n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438;
  wire n18439, n18440, n18443, n18444, n18445, n18446, n18447, n18448;
  wire n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456;
  wire n18457, n18458, n18461, n18462, n18463, n18464, n18465, n18466;
  wire n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474;
  wire n18475, n18476, n18477, n18480, n18481, n18482, n18483, n18484;
  wire n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492;
  wire n18493, n18494, n18495, n18496, n18499, n18500, n18501, n18502;
  wire n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510;
  wire n18511, n18512, n18513, n18514, n18515, n18518, n18519, n18520;
  wire n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528;
  wire n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536;
  wire n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544;
  wire n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552;
  wire n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560;
  wire n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568;
  wire n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576;
  wire n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584;
  wire n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592;
  wire n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600;
  wire n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608;
  wire n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616;
  wire n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624;
  wire n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632;
  wire n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640;
  wire n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648;
  wire n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656;
  wire n18657, n18658, n18659, n18660, n18661, n18663, n18664, n18665;
  wire n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673;
  wire n18674, n18675, n18676, n18677, n18678, n18679, n18682, n18683;
  wire n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691;
  wire n18692, n18693, n18694, n18697, n18698, n18699, n18700, n18701;
  wire n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709;
  wire n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719;
  wire n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727;
  wire n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735;
  wire n18736, n18737, n18738, n18739, n18742, n18743, n18744, n18745;
  wire n18746, n18747, n18748, n18749, n18750, n18751, n18754, n18755;
  wire n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763;
  wire n18764, n18765, n18768, n18769, n18770, n18771, n18772, n18773;
  wire n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781;
  wire n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789;
  wire n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797;
  wire n18798, n18799, n18800, n18801, n18802, n18805, n18806, n18807;
  wire n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815;
  wire n18816, n18817, n18818, n18819, n18820, n18821, n18824, n18825;
  wire n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833;
  wire n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841;
  wire n18842, n18843, n18844, n18847, n18848, n18849, n18850, n18851;
  wire n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859;
  wire n18860, n18861, n18862, n18863, n18864, n18867, n18868, n18869;
  wire n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877;
  wire n18878, n18879, n18880, n18881, n18884, n18885, n18886, n18887;
  wire n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895;
  wire n18896, n18897, n18898, n18899, n18900, n18903, n18904, n18905;
  wire n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913;
  wire n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921;
  wire n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929;
  wire n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937;
  wire n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945;
  wire n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953;
  wire n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961;
  wire n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969;
  wire n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977;
  wire n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985;
  wire n18986, n18987, n18989, n18990, n18991, n18992, n18995, n18996;
  wire n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004;
  wire n19005, n19006, n19007, n19010, n19011, n19012, n19013, n19014;
  wire n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022;
  wire n19023, n19026, n19027, n19028, n19029, n19030, n19031, n19032;
  wire n19033, n19034, n19035, n19036, n19037, n19040, n19041, n19042;
  wire n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050;
  wire n19051, n19052, n19055, n19056, n19057, n19058, n19059, n19060;
  wire n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068;
  wire n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076;
  wire n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084;
  wire n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094;
  wire n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102;
  wire n19103, n19106, n19107, n19108, n19109, n19110, n19111, n19112;
  wire n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120;
  wire n19121, n19122, n19125, n19126, n19127, n19128, n19129, n19130;
  wire n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138;
  wire n19139, n19140, n19141, n19144, n19145, n19146, n19147, n19148;
  wire n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156;
  wire n19157, n19158, n19159, n19160, n19163, n19164, n19165, n19166;
  wire n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174;
  wire n19175, n19176, n19177, n19178, n19179, n19182, n19183, n19184;
  wire n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192;
  wire n19193, n19194, n19195, n19196, n19197, n19200, n19201, n19202;
  wire n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210;
  wire n19211, n19212, n19213, n19214, n19217, n19218, n19219, n19220;
  wire n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228;
  wire n19229, n19230, n19231, n19232, n19235, n19236, n19237, n19238;
  wire n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246;
  wire n19247, n19248, n19249, n19252, n19253, n19254, n19255, n19256;
  wire n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264;
  wire n19265, n19266, n19267, n19268, n19269, n19272, n19273, n19274;
  wire n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282;
  wire n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290;
  wire n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298;
  wire n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306;
  wire n19307, n19308, n19309, n19310, n19311, n19312, n19314, n19315;
  wire n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323;
  wire n19324, n19325, n19326, n19327, n19328, n19329, n19332, n19333;
  wire n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341;
  wire n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349;
  wire n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357;
  wire n19358, n19359, n19360, n19363, n19364, n19365, n19366, n19367;
  wire n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375;
  wire n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385;
  wire n19386, n19387, n19388, n19389, n19390, n19391, n19394, n19395;
  wire n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403;
  wire n19404, n19405, n19406, n19409, n19410, n19411, n19412, n19413;
  wire n19414, n19415, n19416, n19417, n19418, n19419, n19422, n19423;
  wire n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431;
  wire n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441;
  wire n19442, n19443, n19444, n19447, n19448, n19449, n19450, n19451;
  wire n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459;
  wire n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467;
  wire n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475;
  wire n19476, n19477, n19478, n19479, n19480, n19483, n19484, n19485;
  wire n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493;
  wire n19494, n19495, n19496, n19497, n19498, n19499, n19502, n19503;
  wire n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511;
  wire n19512, n19513, n19514, n19515, n19516, n19517, n19520, n19521;
  wire n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529;
  wire n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537;
  wire n19538, n19539, n19540, n19541, n19542, n19543, n19546, n19547;
  wire n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555;
  wire n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563;
  wire n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571;
  wire n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579;
  wire n19580, n19581, n19582, n19583, n19584, n19587, n19588, n19589;
  wire n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597;
  wire n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605;
  wire n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613;
  wire n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621;
  wire n19622, n19623, n19624, n19625, n19626, n19627, n19629, n19630;
  wire n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638;
  wire n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19648;
  wire n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656;
  wire n19657, n19658, n19659, n19660, n19663, n19664, n19665, n19666;
  wire n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674;
  wire n19675, n19676, n19679, n19680, n19681, n19682, n19683, n19684;
  wire n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19694;
  wire n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702;
  wire n19703, n19704, n19705, n19706, n19707, n19710, n19711, n19712;
  wire n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720;
  wire n19721, n19722, n19723, n19726, n19727, n19728, n19729, n19730;
  wire n19731, n19732, n19733, n19734, n19735, n19738, n19739, n19740;
  wire n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748;
  wire n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758;
  wire n19759, n19760, n19763, n19764, n19765, n19766, n19767, n19768;
  wire n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776;
  wire n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784;
  wire n19785, n19786, n19789, n19790, n19791, n19792, n19793, n19794;
  wire n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802;
  wire n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19812;
  wire n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820;
  wire n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828;
  wire n19829, n19830, n19833, n19834, n19835, n19836, n19837, n19838;
  wire n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846;
  wire n19847, n19848, n19851, n19852, n19853, n19854, n19855, n19856;
  wire n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864;
  wire n19865, n19866, n19867, n19868, n19871, n19872, n19873, n19874;
  wire n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882;
  wire n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890;
  wire n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19900;
  wire n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908;
  wire n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916;
  wire n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924;
  wire n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932;
  wire n19933, n19934, n19935, n19936, n19937, n19938, n19940, n19941;
  wire n19942, n19943, n19944, n19945, n19948, n19949, n19950, n19951;
  wire n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959;
  wire n19960, n19963, n19964, n19965, n19966, n19967, n19968, n19969;
  wire n19970, n19971, n19972, n19973, n19974, n19975, n19978, n19979;
  wire n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987;
  wire n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19997;
  wire n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005;
  wire n20006, n20009, n20010, n20011, n20012, n20013, n20014, n20015;
  wire n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023;
  wire n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031;
  wire n20032, n20033, n20034, n20037, n20038, n20039, n20040, n20041;
  wire n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049;
  wire n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057;
  wire n20058, n20059, n20062, n20063, n20064, n20065, n20066, n20067;
  wire n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075;
  wire n20076, n20077, n20078, n20081, n20082, n20083, n20084, n20085;
  wire n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093;
  wire n20094, n20095, n20096, n20097, n20100, n20101, n20102, n20103;
  wire n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111;
  wire n20112, n20113, n20114, n20117, n20118, n20119, n20120, n20121;
  wire n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129;
  wire n20130, n20131, n20132, n20135, n20136, n20137, n20138, n20139;
  wire n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147;
  wire n20148, n20149, n20152, n20153, n20154, n20155, n20156, n20157;
  wire n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165;
  wire n20166, n20167, n20168, n20171, n20172, n20173, n20174, n20175;
  wire n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183;
  wire n20184, n20185, n20186, n20187, n20190, n20191, n20192, n20193;
  wire n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201;
  wire n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209;
  wire n20210, n20213, n20214, n20215, n20216, n20217, n20218, n20219;
  wire n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227;
  wire n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235;
  wire n20236, n20237, n20238, n20239, n20240, n20242, n20243, n20244;
  wire n20245, n20246, n20247, n20250, n20251, n20252, n20253, n20254;
  wire n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262;
  wire n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272;
  wire n20273, n20274, n20275, n20276, n20277, n20280, n20281, n20282;
  wire n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290;
  wire n20291, n20292, n20295, n20296, n20297, n20298, n20299, n20300;
  wire n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20310;
  wire n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318;
  wire n20319, n20320, n20323, n20324, n20325, n20326, n20327, n20328;
  wire n20329, n20330, n20331, n20332, n20335, n20336, n20337, n20338;
  wire n20339, n20340, n20341, n20342, n20343, n20344, n20347, n20348;
  wire n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356;
  wire n20357, n20358, n20359, n20360, n20361, n20362, n20365, n20366;
  wire n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374;
  wire n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382;
  wire n20383, n20384, n20385, n20386, n20387, n20390, n20391, n20392;
  wire n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400;
  wire n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408;
  wire n20409, n20410, n20411, n20412, n20413, n20416, n20417, n20418;
  wire n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426;
  wire n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20436;
  wire n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444;
  wire n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452;
  wire n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460;
  wire n20461, n20462, n20463, n20464, n20465, n20466, n20469, n20470;
  wire n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478;
  wire n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20488;
  wire n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496;
  wire n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504;
  wire n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512;
  wire n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520;
  wire n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528;
  wire n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536;
  wire n20537, n20538, n20540, n20541, n20542, n20543, n20544, n20545;
  wire n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553;
  wire n20554, n20555, n20556, n20559, n20560, n20561, n20562, n20563;
  wire n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571;
  wire n20572, n20575, n20576, n20577, n20578, n20579, n20580, n20581;
  wire n20582, n20583, n20584, n20585, n20586, n20587, n20590, n20591;
  wire n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599;
  wire n20600, n20601, n20602, n20603, n20606, n20607, n20608, n20609;
  wire n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617;
  wire n20618, n20619, n20622, n20623, n20624, n20625, n20626, n20627;
  wire n20628, n20629, n20630, n20631, n20634, n20635, n20636, n20637;
  wire n20638, n20639, n20640, n20641, n20642, n20643, n20646, n20647;
  wire n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655;
  wire n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665;
  wire n20666, n20667, n20668, n20671, n20672, n20673, n20674, n20675;
  wire n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683;
  wire n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691;
  wire n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699;
  wire n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707;
  wire n20708, n20709, n20712, n20713, n20714, n20715, n20716, n20717;
  wire n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725;
  wire n20726, n20727, n20728, n20729, n20730, n20733, n20734, n20735;
  wire n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743;
  wire n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751;
  wire n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759;
  wire n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767;
  wire n20768, n20769, n20770, n20771, n20774, n20775, n20776, n20777;
  wire n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785;
  wire n20786, n20787, n20788, n20789, n20790, n20793, n20794, n20795;
  wire n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803;
  wire n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811;
  wire n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819;
  wire n20820, n20821, n20822, n20823, n20824, n20826, n20827, n20828;
  wire n20829, n20830, n20833, n20834, n20835, n20836, n20837, n20838;
  wire n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20848;
  wire n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856;
  wire n20857, n20858, n20859, n20860, n20861, n20862, n20865, n20866;
  wire n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874;
  wire n20875, n20876, n20879, n20880, n20881, n20882, n20883, n20884;
  wire n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892;
  wire n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900;
  wire n20901, n20902, n20905, n20906, n20907, n20908, n20909, n20910;
  wire n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918;
  wire n20919, n20920, n20921, n20922, n20925, n20926, n20927, n20928;
  wire n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936;
  wire n20937, n20938, n20939, n20940, n20941, n20944, n20945, n20946;
  wire n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954;
  wire n20955, n20956, n20957, n20958, n20959, n20960, n20963, n20964;
  wire n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972;
  wire n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20982;
  wire n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990;
  wire n20991, n20992, n20993, n20994, n20995, n20996, n20999, n21000;
  wire n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008;
  wire n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21018;
  wire n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026;
  wire n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034;
  wire n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044;
  wire n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052;
  wire n21053, n21056, n21057, n21058, n21059, n21060, n21061, n21062;
  wire n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070;
  wire n21071, n21072, n21075, n21076, n21077, n21078, n21079, n21080;
  wire n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088;
  wire n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096;
  wire n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104;
  wire n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21113;
  wire n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121;
  wire n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21131;
  wire n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139;
  wire n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147;
  wire n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155;
  wire n21156, n21157, n21158, n21159, n21162, n21163, n21164, n21165;
  wire n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173;
  wire n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183;
  wire n21184, n21185, n21188, n21189, n21190, n21191, n21192, n21193;
  wire n21194, n21195, n21196, n21197, n21198, n21201, n21202, n21203;
  wire n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211;
  wire n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219;
  wire n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227;
  wire n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235;
  wire n21236, n21237, n21238, n21239, n21240, n21243, n21244, n21245;
  wire n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253;
  wire n21254, n21255, n21256, n21257, n21258, n21259, n21262, n21263;
  wire n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271;
  wire n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279;
  wire n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289;
  wire n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297;
  wire n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305;
  wire n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21315;
  wire n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323;
  wire n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331;
  wire n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341;
  wire n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349;
  wire n21350, n21353, n21354, n21355, n21356, n21357, n21358, n21359;
  wire n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367;
  wire n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375;
  wire n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383;
  wire n21384, n21385, n21387, n21388, n21389, n21390, n21391, n21392;
  wire n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400;
  wire n21401, n21402, n21403, n21406, n21407, n21408, n21409, n21410;
  wire n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418;
  wire n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428;
  wire n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21438;
  wire n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446;
  wire n21447, n21448, n21449, n21450, n21453, n21454, n21455, n21456;
  wire n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21466;
  wire n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474;
  wire n21475, n21476, n21479, n21480, n21481, n21482, n21483, n21484;
  wire n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492;
  wire n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500;
  wire n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508;
  wire n21509, n21510, n21511, n21512, n21515, n21516, n21517, n21518;
  wire n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526;
  wire n21527, n21528, n21529, n21530, n21531, n21534, n21535, n21536;
  wire n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544;
  wire n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552;
  wire n21553, n21554, n21557, n21558, n21559, n21560, n21561, n21562;
  wire n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570;
  wire n21571, n21572, n21573, n21574, n21577, n21578, n21579, n21580;
  wire n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588;
  wire n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596;
  wire n21597, n21600, n21601, n21602, n21603, n21604, n21605, n21606;
  wire n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614;
  wire n21615, n21616, n21619, n21620, n21621, n21622, n21623, n21624;
  wire n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632;
  wire n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640;
  wire n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648;
  wire n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656;
  wire n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21667;
  wire n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675;
  wire n21676, n21677, n21678, n21679, n21680, n21681, n21684, n21685;
  wire n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693;
  wire n21694, n21695, n21698, n21699, n21700, n21701, n21702, n21703;
  wire n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711;
  wire n21712, n21713, n21714, n21715, n21718, n21719, n21720, n21721;
  wire n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729;
  wire n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737;
  wire n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747;
  wire n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755;
  wire n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765;
  wire n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21775;
  wire n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783;
  wire n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791;
  wire n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21801;
  wire n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809;
  wire n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817;
  wire n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827;
  wire n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835;
  wire n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845;
  wire n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21855;
  wire n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863;
  wire n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871;
  wire n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881;
  wire n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889;
  wire n21890, n21893, n21894, n21895, n21896, n21897, n21898, n21899;
  wire n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907;
  wire n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915;
  wire n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21924;
  wire n21925, n21926, n21927, n21928, n21929, n21932, n21933, n21934;
  wire n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942;
  wire n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950;
  wire n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958;
  wire n21959, n21960, n21963, n21964, n21965, n21966, n21967, n21968;
  wire n21969, n21970, n21971, n21972, n21975, n21976, n21977, n21978;
  wire n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986;
  wire n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994;
  wire n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002;
  wire n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010;
  wire n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020;
  wire n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028;
  wire n22029, n22032, n22033, n22034, n22035, n22036, n22037, n22038;
  wire n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046;
  wire n22047, n22048, n22051, n22052, n22053, n22054, n22055, n22056;
  wire n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064;
  wire n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072;
  wire n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080;
  wire n22081, n22082, n22085, n22086, n22087, n22088, n22089, n22090;
  wire n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098;
  wire n22099, n22100, n22101, n22104, n22105, n22106, n22107, n22108;
  wire n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116;
  wire n22117, n22118, n22119, n22120, n22123, n22124, n22125, n22126;
  wire n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134;
  wire n22135, n22136, n22137, n22138, n22141, n22142, n22143, n22144;
  wire n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152;
  wire n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160;
  wire n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168;
  wire n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176;
  wire n22177, n22178, n22179, n22180, n22181, n22182, n22184, n22185;
  wire n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193;
  wire n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22203;
  wire n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211;
  wire n22212, n22213, n22214, n22215, n22218, n22219, n22220, n22221;
  wire n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229;
  wire n22230, n22231, n22234, n22235, n22236, n22237, n22238, n22239;
  wire n22240, n22241, n22242, n22243, n22246, n22247, n22248, n22249;
  wire n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22259;
  wire n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267;
  wire n22268, n22269, n22272, n22273, n22274, n22275, n22276, n22277;
  wire n22278, n22279, n22280, n22281, n22284, n22285, n22286, n22287;
  wire n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295;
  wire n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303;
  wire n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311;
  wire n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319;
  wire n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327;
  wire n22328, n22331, n22332, n22333, n22334, n22335, n22336, n22337;
  wire n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345;
  wire n22346, n22347, n22348, n22351, n22352, n22353, n22354, n22355;
  wire n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363;
  wire n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371;
  wire n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381;
  wire n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389;
  wire n22390, n22393, n22394, n22395, n22396, n22397, n22398, n22399;
  wire n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407;
  wire n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415;
  wire n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423;
  wire n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431;
  wire n22433, n22434, n22435, n22436, n22437, n22440, n22441, n22442;
  wire n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450;
  wire n22451, n22452, n22455, n22456, n22457, n22458, n22459, n22460;
  wire n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468;
  wire n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478;
  wire n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486;
  wire n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494;
  wire n22495, n22496, n22499, n22500, n22501, n22502, n22503, n22504;
  wire n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512;
  wire n22513, n22514, n22517, n22518, n22519, n22520, n22521, n22522;
  wire n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530;
  wire n22531, n22532, n22533, n22536, n22537, n22538, n22539, n22540;
  wire n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548;
  wire n22549, n22550, n22551, n22552, n22555, n22556, n22557, n22558;
  wire n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566;
  wire n22567, n22568, n22569, n22570, n22573, n22574, n22575, n22576;
  wire n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584;
  wire n22585, n22586, n22587, n22590, n22591, n22592, n22593, n22594;
  wire n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602;
  wire n22603, n22604, n22605, n22606, n22609, n22610, n22611, n22612;
  wire n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620;
  wire n22621, n22622, n22623, n22624, n22625, n22628, n22629, n22630;
  wire n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638;
  wire n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646;
  wire n22647, n22648, n22649, n22650, n22653, n22654, n22655, n22656;
  wire n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664;
  wire n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672;
  wire n22673, n22674, n22676, n22677, n22678, n22679, n22680, n22681;
  wire n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689;
  wire n22690, n22691, n22692, n22695, n22696, n22697, n22698, n22699;
  wire n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707;
  wire n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717;
  wire n22718, n22719, n22722, n22723, n22724, n22725, n22726, n22727;
  wire n22728, n22729, n22730, n22731, n22734, n22735, n22736, n22737;
  wire n22738, n22739, n22740, n22741, n22742, n22743, n22746, n22747;
  wire n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755;
  wire n22756, n22757, n22758, n22759, n22760, n22761, n22764, n22765;
  wire n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773;
  wire n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781;
  wire n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22791;
  wire n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799;
  wire n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807;
  wire n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815;
  wire n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22825;
  wire n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833;
  wire n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841;
  wire n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851;
  wire n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859;
  wire n22860, n22863, n22864, n22865, n22866, n22867, n22868, n22869;
  wire n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877;
  wire n22878, n22881, n22882, n22883, n22884, n22885, n22886, n22887;
  wire n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895;
  wire n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903;
  wire n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911;
  wire n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920;
  wire n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928;
  wire n22929, n22932, n22933, n22934, n22935, n22936, n22937, n22938;
  wire n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946;
  wire n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956;
  wire n22957, n22958, n22961, n22962, n22963, n22964, n22965, n22966;
  wire n22967, n22968, n22969, n22970, n22971, n22974, n22975, n22976;
  wire n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984;
  wire n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994;
  wire n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002;
  wire n23003, n23004, n23005, n23006, n23007, n23010, n23011, n23012;
  wire n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020;
  wire n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23030;
  wire n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038;
  wire n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046;
  wire n23047, n23048, n23051, n23052, n23053, n23054, n23055, n23056;
  wire n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064;
  wire n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23074;
  wire n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082;
  wire n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090;
  wire n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100;
  wire n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108;
  wire n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116;
  wire n23117, n23118, n23119, n23120, n23121, n23124, n23125, n23126;
  wire n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134;
  wire n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142;
  wire n23143, n23144, n23145, n23146, n23148, n23149, n23150, n23151;
  wire n23152, n23155, n23156, n23157, n23158, n23159, n23160, n23161;
  wire n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23171;
  wire n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179;
  wire n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187;
  wire n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195;
  wire n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205;
  wire n23206, n23207, n23208, n23209, n23212, n23213, n23214, n23215;
  wire n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223;
  wire n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231;
  wire n23232, n23233, n23234, n23237, n23238, n23239, n23240, n23241;
  wire n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249;
  wire n23250, n23251, n23252, n23255, n23256, n23257, n23258, n23259;
  wire n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267;
  wire n23268, n23269, n23272, n23273, n23274, n23275, n23276, n23277;
  wire n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285;
  wire n23286, n23287, n23288, n23291, n23292, n23293, n23294, n23295;
  wire n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303;
  wire n23304, n23305, n23306, n23307, n23310, n23311, n23312, n23313;
  wire n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321;
  wire n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329;
  wire n23330, n23331, n23332, n23335, n23336, n23337, n23338, n23339;
  wire n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347;
  wire n23348, n23349, n23350, n23351, n23352, n23355, n23356, n23357;
  wire n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365;
  wire n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23374;
  wire n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382;
  wire n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23392;
  wire n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400;
  wire n23401, n23404, n23405, n23406, n23407, n23408, n23409, n23410;
  wire n23411, n23412, n23413, n23416, n23417, n23418, n23419, n23420;
  wire n23421, n23422, n23423, n23424, n23425, n23428, n23429, n23430;
  wire n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438;
  wire n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23448;
  wire n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456;
  wire n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464;
  wire n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472;
  wire n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480;
  wire n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23490;
  wire n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498;
  wire n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506;
  wire n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516;
  wire n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524;
  wire n23525, n23528, n23529, n23530, n23531, n23532, n23533, n23534;
  wire n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542;
  wire n23543, n23546, n23547, n23548, n23549, n23550, n23551, n23552;
  wire n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560;
  wire n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568;
  wire n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578;
  wire n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586;
  wire n23587, n23588, n23589, n23590, n23591, n23592, n23594, n23595;
  wire n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603;
  wire n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611;
  wire n23612, n23615, n23616, n23617, n23618, n23619, n23620, n23621;
  wire n23622, n23623, n23624, n23627, n23628, n23629, n23630, n23631;
  wire n23632, n23633, n23634, n23635, n23636, n23637, n23640, n23641;
  wire n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649;
  wire n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659;
  wire n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667;
  wire n23668, n23669, n23670, n23671, n23672, n23673, n23676, n23677;
  wire n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685;
  wire n23686, n23687, n23688, n23691, n23692, n23693, n23694, n23695;
  wire n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703;
  wire n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711;
  wire n23712, n23713, n23714, n23715, n23716, n23717, n23720, n23721;
  wire n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729;
  wire n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23739;
  wire n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747;
  wire n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755;
  wire n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763;
  wire n23764, n23765, n23766, n23767, n23770, n23771, n23772, n23773;
  wire n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781;
  wire n23782, n23783, n23784, n23785, n23786, n23789, n23790, n23791;
  wire n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799;
  wire n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807;
  wire n23808, n23810, n23811, n23812, n23813, n23814, n23815, n23818;
  wire n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826;
  wire n23827, n23828, n23831, n23832, n23833, n23834, n23835, n23836;
  wire n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844;
  wire n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852;
  wire n23853, n23854, n23855, n23858, n23859, n23860, n23861, n23862;
  wire n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23872;
  wire n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880;
  wire n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888;
  wire n23889, n23890, n23891, n23892, n23893, n23894, n23897, n23898;
  wire n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906;
  wire n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23916;
  wire n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924;
  wire n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932;
  wire n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942;
  wire n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950;
  wire n23951, n23954, n23955, n23956, n23957, n23958, n23959, n23960;
  wire n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968;
  wire n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976;
  wire n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986;
  wire n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994;
  wire n23995, n23996, n23999, n24000, n24001, n24002, n24003, n24004;
  wire n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012;
  wire n24013, n24014, n24015, n24016, n24018, n24019, n24020, n24021;
  wire n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029;
  wire n24030, n24031, n24032, n24033, n24036, n24037, n24038, n24039;
  wire n24040, n24041, n24042, n24043, n24044, n24045, n24048, n24049;
  wire n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057;
  wire n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067;
  wire n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075;
  wire n24076, n24077, n24080, n24081, n24082, n24083, n24084, n24085;
  wire n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093;
  wire n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101;
  wire n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109;
  wire n24110, n24113, n24114, n24115, n24116, n24117, n24118, n24119;
  wire n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127;
  wire n24128, n24129, n24132, n24133, n24134, n24135, n24136, n24137;
  wire n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145;
  wire n24146, n24147, n24148, n24151, n24152, n24153, n24154, n24155;
  wire n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163;
  wire n24164, n24165, n24166, n24169, n24170, n24171, n24172, n24173;
  wire n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181;
  wire n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189;
  wire n24190, n24191, n24194, n24195, n24196, n24197, n24198, n24199;
  wire n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207;
  wire n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215;
  wire n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224;
  wire n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232;
  wire n24233, n24234, n24235, n24238, n24239, n24240, n24241, n24242;
  wire n24243, n24244, n24245, n24246, n24247, n24250, n24251, n24252;
  wire n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260;
  wire n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270;
  wire n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278;
  wire n24279, n24280, n24281, n24282, n24283, n24284, n24287, n24288;
  wire n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296;
  wire n24297, n24298, n24299, n24302, n24303, n24304, n24305, n24306;
  wire n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314;
  wire n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322;
  wire n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332;
  wire n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340;
  wire n24341, n24344, n24345, n24346, n24347, n24348, n24349, n24350;
  wire n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358;
  wire n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366;
  wire n24367, n24368, n24369, n24370, n24371, n24372, n24375, n24376;
  wire n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384;
  wire n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24394;
  wire n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402;
  wire n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410;
  wire n24411, n24413, n24414, n24415, n24416, n24417, n24420, n24421;
  wire n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429;
  wire n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437;
  wire n24438, n24439, n24440, n24441, n24444, n24445, n24446, n24447;
  wire n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455;
  wire n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465;
  wire n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473;
  wire n24474, n24475, n24476, n24479, n24480, n24481, n24482, n24483;
  wire n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491;
  wire n24492, n24493, n24494, n24495, n24498, n24499, n24500, n24501;
  wire n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509;
  wire n24510, n24511, n24512, n24513, n24514, n24517, n24518, n24519;
  wire n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527;
  wire n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535;
  wire n24536, n24537, n24540, n24541, n24542, n24543, n24544, n24545;
  wire n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553;
  wire n24554, n24555, n24556, n24559, n24560, n24561, n24562, n24563;
  wire n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571;
  wire n24572, n24573, n24574, n24575, n24578, n24579, n24580, n24581;
  wire n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589;
  wire n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597;
  wire n24598, n24600, n24601, n24602, n24603, n24604, n24605, n24606;
  wire n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614;
  wire n24615, n24618, n24619, n24620, n24621, n24622, n24623, n24624;
  wire n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632;
  wire n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640;
  wire n24641, n24642, n24643, n24646, n24647, n24648, n24649, n24650;
  wire n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658;
  wire n24659, n24660, n24661, n24662, n24665, n24666, n24667, n24668;
  wire n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676;
  wire n24677, n24678, n24679, n24680, n24681, n24684, n24685, n24686;
  wire n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694;
  wire n24695, n24696, n24697, n24698, n24699, n24700, n24703, n24704;
  wire n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712;
  wire n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720;
  wire n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730;
  wire n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738;
  wire n24739, n24742, n24743, n24744, n24745, n24746, n24747, n24748;
  wire n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756;
  wire n24757, n24758, n24761, n24762, n24763, n24764, n24765, n24766;
  wire n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774;
  wire n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24783;
  wire n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791;
  wire n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799;
  wire n24800, n24803, n24804, n24805, n24806, n24807, n24808, n24809;
  wire n24810, n24811, n24812, n24815, n24816, n24817, n24818, n24819;
  wire n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827;
  wire n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835;
  wire n24836, n24839, n24840, n24841, n24842, n24843, n24844, n24845;
  wire n24846, n24847, n24848, n24849, n24850, n24851, n24854, n24855;
  wire n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863;
  wire n24864, n24865, n24866, n24867, n24868, n24869, n24872, n24873;
  wire n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881;
  wire n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24891;
  wire n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899;
  wire n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907;
  wire n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915;
  wire n24916, n24917, n24918, n24919, n24922, n24923, n24924, n24925;
  wire n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933;
  wire n24934, n24935, n24936, n24937, n24938, n24941, n24942, n24943;
  wire n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951;
  wire n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24960;
  wire n24961, n24962, n24963, n24964, n24967, n24968, n24969, n24970;
  wire n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978;
  wire n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986;
  wire n24987, n24988, n24989, n24992, n24993, n24994, n24995, n24996;
  wire n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004;
  wire n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014;
  wire n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022;
  wire n25023, n25024, n25025, n25028, n25029, n25030, n25031, n25032;
  wire n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040;
  wire n25041, n25042, n25043, n25044, n25047, n25048, n25049, n25050;
  wire n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058;
  wire n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066;
  wire n25067, n25070, n25071, n25072, n25073, n25074, n25075, n25076;
  wire n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084;
  wire n25085, n25086, n25089, n25090, n25091, n25092, n25093, n25094;
  wire n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102;
  wire n25103, n25104, n25105, n25108, n25109, n25110, n25111, n25112;
  wire n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120;
  wire n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128;
  wire n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137;
  wire n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145;
  wire n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153;
  wire n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161;
  wire n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169;
  wire n25170, n25171, n25174, n25175, n25176, n25177, n25178, n25179;
  wire n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187;
  wire n25188, n25189, n25190, n25193, n25194, n25195, n25196, n25197;
  wire n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205;
  wire n25206, n25207, n25208, n25209, n25212, n25213, n25214, n25215;
  wire n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223;
  wire n25224, n25225, n25226, n25227, n25228, n25229, n25232, n25233;
  wire n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241;
  wire n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25251;
  wire n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259;
  wire n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267;
  wire n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277;
  wire n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285;
  wire n25286, n25287, n25288, n25289, n25290, n25292, n25293, n25294;
  wire n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302;
  wire n25303, n25304, n25305, n25306, n25307, n25308, n25311, n25312;
  wire n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320;
  wire n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330;
  wire n25331, n25332, n25335, n25336, n25337, n25338, n25339, n25340;
  wire n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348;
  wire n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356;
  wire n25357, n25360, n25361, n25362, n25363, n25364, n25365, n25366;
  wire n25367, n25368, n25369, n25370, n25371, n25374, n25375, n25376;
  wire n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384;
  wire n25385, n25386, n25387, n25388, n25391, n25392, n25393, n25394;
  wire n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402;
  wire n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410;
  wire n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418;
  wire n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426;
  wire n25427, n25428, n25429, n25432, n25433, n25434, n25435, n25436;
  wire n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444;
  wire n25445, n25446, n25447, n25448, n25449, n25451, n25452, n25453;
  wire n25454, n25457, n25458, n25459, n25460, n25461, n25462, n25463;
  wire n25464, n25465, n25466, n25469, n25470, n25471, n25472, n25473;
  wire n25474, n25475, n25476, n25477, n25478, n25479, n25482, n25483;
  wire n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491;
  wire n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499;
  wire n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509;
  wire n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517;
  wire n25518, n25521, n25522, n25523, n25524, n25525, n25526, n25527;
  wire n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535;
  wire n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543;
  wire n25544, n25545, n25546, n25549, n25550, n25551, n25552, n25553;
  wire n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561;
  wire n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569;
  wire n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577;
  wire n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587;
  wire n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595;
  wire n25596, n25597, n25598, n25599, n25600, n25602, n25603, n25604;
  wire n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612;
  wire n25613, n25614, n25615, n25616, n25617, n25620, n25621, n25622;
  wire n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630;
  wire n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638;
  wire n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646;
  wire n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654;
  wire n25655, n25656, n25657, n25660, n25661, n25662, n25663, n25664;
  wire n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672;
  wire n25673, n25674, n25675, n25676, n25679, n25680, n25681, n25682;
  wire n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690;
  wire n25691, n25692, n25693, n25694, n25695, n25698, n25699, n25700;
  wire n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708;
  wire n25709, n25710, n25711, n25712, n25713, n25716, n25717, n25718;
  wire n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726;
  wire n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734;
  wire n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742;
  wire n25743, n25745, n25746, n25747, n25748, n25749, n25750, n25751;
  wire n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759;
  wire n25760, n25761, n25764, n25765, n25766, n25767, n25768, n25769;
  wire n25770, n25771, n25772, n25773, n25776, n25777, n25778, n25779;
  wire n25780, n25781, n25782, n25783, n25784, n25785, n25788, n25789;
  wire n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797;
  wire n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807;
  wire n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815;
  wire n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823;
  wire n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831;
  wire n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839;
  wire n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847;
  wire n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855;
  wire n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863;
  wire n25864, n25865, n25866, n25869, n25870, n25871, n25872, n25873;
  wire n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881;
  wire n25882, n25883, n25884, n25885, n25886, n25888, n25889, n25890;
  wire n25891, n25894, n25895, n25896, n25897, n25898, n25899, n25900;
  wire n25901, n25902, n25903, n25906, n25907, n25908, n25909, n25910;
  wire n25911, n25912, n25913, n25914, n25915, n25918, n25919, n25920;
  wire n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25930;
  wire n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938;
  wire n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946;
  wire n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954;
  wire n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964;
  wire n25965, n25966, n25967, n25968, n25969, n25972, n25973, n25974;
  wire n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982;
  wire n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990;
  wire n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998;
  wire n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006;
  wire n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014;
  wire n26015, n26016, n26018, n26019, n26020, n26021, n26022, n26023;
  wire n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031;
  wire n26032, n26033, n26036, n26037, n26038, n26039, n26040, n26041;
  wire n26042, n26043, n26044, n26045, n26046, n26049, n26050, n26051;
  wire n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26061;
  wire n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069;
  wire n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077;
  wire n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087;
  wire n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095;
  wire n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103;
  wire n26104, n26105, n26106, n26107, n26108, n26109, n26112, n26113;
  wire n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121;
  wire n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129;
  wire n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137;
  wire n26138, n26139, n26141, n26142, n26143, n26146, n26147, n26148;
  wire n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26158;
  wire n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166;
  wire n26167, n26170, n26171, n26172, n26173, n26174, n26175, n26176;
  wire n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184;
  wire n26185, n26186, n26187, n26188, n26189, n26190, n26193, n26194;
  wire n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202;
  wire n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210;
  wire n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218;
  wire n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226;
  wire n26227, n26228, n26231, n26232, n26233, n26234, n26235, n26236;
  wire n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244;
  wire n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252;
  wire n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260;
  wire n26261, n26262, n26264, n26265, n26266, n26269, n26270, n26271;
  wire n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26281;
  wire n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289;
  wire n26290, n26293, n26294, n26295, n26296, n26297, n26298, n26299;
  wire n26300, n26301, n26302, n26303, n26306, n26307, n26308, n26309;
  wire n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317;
  wire n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325;
  wire n26326, n26327, n26328, n26329, n26330, n26331, n26334, n26335;
  wire n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343;
  wire n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351;
  wire n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359;
  wire n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367;
  wire n26368, n26369, n26370, n26371, n26372, n26374, n26375, n26376;
  wire n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384;
  wire n26385, n26386, n26389, n26390, n26391, n26392, n26393, n26394;
  wire n26395, n26396, n26397, n26398, n26401, n26402, n26403, n26404;
  wire n26405, n26406, n26407, n26408, n26409, n26410, n26413, n26414;
  wire n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422;
  wire n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430;
  wire n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438;
  wire n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446;
  wire n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454;
  wire n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462;
  wire n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470;
  wire n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26479;
  wire n26480, n26481, n26484, n26485, n26486, n26487, n26488, n26489;
  wire n26490, n26491, n26492, n26493, n26496, n26497, n26498, n26499;
  wire n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507;
  wire n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515;
  wire n26516, n26517, n26518, n26519, n26522, n26523, n26524, n26525;
  wire n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533;
  wire n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541;
  wire n26542, n26543, n26544, n26547, n26548, n26549, n26550, n26551;
  wire n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559;
  wire n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567;
  wire n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575;
  wire n26576, n26577, n26578, n26580, n26581, n26582, n26583, n26586;
  wire n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594;
  wire n26595, n26598, n26599, n26600, n26601, n26602, n26603, n26604;
  wire n26605, n26606, n26609, n26610, n26611, n26612, n26613, n26614;
  wire n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622;
  wire n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630;
  wire n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638;
  wire n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646;
  wire n26647, n26648, n26649, n26652, n26653, n26654, n26655, n26656;
  wire n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664;
  wire n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672;
  wire n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681;
  wire n26682, n26683, n26684, n26685, n26686, n26689, n26690, n26691;
  wire n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26701;
  wire n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709;
  wire n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717;
  wire n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727;
  wire n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735;
  wire n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743;
  wire n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751;
  wire n26752, n26753, n26754, n26755, n26756, n26758, n26759, n26760;
  wire n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768;
  wire n26769, n26770, n26771, n26772, n26773, n26776, n26777, n26778;
  wire n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786;
  wire n26787, n26790, n26791, n26792, n26793, n26794, n26795, n26796;
  wire n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804;
  wire n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814;
  wire n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822;
  wire n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830;
  wire n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838;
  wire n26840, n26841, n26842, n26843, n26844, n26845, n26848, n26849;
  wire n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857;
  wire n26858, n26859, n26860, n26861, n26862, n26865, n26866, n26867;
  wire n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875;
  wire n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26885;
  wire n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893;
  wire n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901;
  wire n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909;
  wire n26910, n26911, n26912, n26913, n26915, n26916, n26917, n26918;
  wire n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926;
  wire n26927, n26930, n26931, n26932, n26933, n26934, n26935, n26936;
  wire n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944;
  wire n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952;
  wire n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960;
  wire n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968;
  wire n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976;
  wire n26977, n26978, n26979, n26980, n26981, n26982, n26984, n26985;
  wire n26986, n26989, n26990, n26991, n26992, n26993, n26994, n26995;
  wire n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003;
  wire n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011;
  wire n27012, n27015, n27016, n27017, n27018, n27019, n27020, n27021;
  wire n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029;
  wire n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037;
  wire n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045;
  wire n27046, n27048, n27049, n27050, n27051, n27054, n27055, n27056;
  wire n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064;
  wire n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072;
  wire n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080;
  wire n27081, n27084, n27085, n27086, n27087, n27088, n27089, n27090;
  wire n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098;
  wire n27099, n27100, n27101, n27102, n27103, n27104, n27106, n27107;
  wire n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115;
  wire n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123;
  wire n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131;
  wire n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139;
  wire n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147;
  wire n27148, n27149, n27150, n27152, n27153, n27154, n27155, n27156;
  wire n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164;
  wire n27165, n27166, n27167, n27168, n27171, n27172, n27173, n27174;
  wire n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182;
  wire n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190;
  wire n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27199;
  wire n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207;
  wire n27208, n27209, n27210, n27211, n27212, n27213, n27216, n27217;
  wire n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225;
  wire n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233;
  wire n27234, n27235, n27237, n27238, n27239, n27240, n27241, n27242;
  wire n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250;
  wire n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258;
  wire n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27267;
  wire n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275;
  wire n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283;
  wire n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291;
  wire n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300;
  wire n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308;
  wire n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317;
  wire n_4, n_5, n_6, n_7, n_8, n_10, n_11, n_12;
  wire n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21;
  wire n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29;
  wire n_34, n_35, n_36, n_37, n_38, n_39, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_59, n_61, n_62, n_63;
  wire n_64, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_89, n_90, n_91, n_92, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_215, n_216, n_217, n_218, n_223;
  wire n_224, n_225, n_226, n_228, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_321, n_322;
  wire n_323, n_324, n_326, n_327, n_328, n_329, n_330, n_331;
  wire n_332, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372;
  wire n_373, n_374, n_375, n_376, n_381, n_382, n_383, n_384;
  wire n_385, n_390, n_391, n_392, n_393, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451;
  wire n_452, n_453, n_454, n_459, n_460, n_461, n_462, n_467;
  wire n_468, n_469, n_470, n_471, n_472, n_473, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_503, n_504, n_505, n_506, n_507;
  wire n_508, n_509, n_511, n_512, n_513, n_514, n_515, n_516;
  wire n_517, n_518, n_519, n_520, n_521, n_522, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_535, n_536, n_537;
  wire n_538, n_543, n_544, n_545, n_546, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_579, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_604, n_605, n_606, n_607, n_608, n_613, n_614;
  wire n_615, n_616, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_658, n_659, n_660;
  wire n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668;
  wire n_669, n_674, n_675, n_676, n_677, n_678, n_679, n_680;
  wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_699, n_700, n_701;
  wire n_702, n_703, n_704, n_705, n_707, n_708, n_709, n_710;
  wire n_715, n_716, n_717, n_718, n_723, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_734, n_735, n_736, n_737, n_738;
  wire n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_750;
  wire n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758;
  wire n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766;
  wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
  wire n_775, n_776, n_777, n_778, n_783, n_784, n_785, n_786;
  wire n_787, n_788, n_789, n_791, n_792, n_793, n_794, n_799;
  wire n_800, n_801, n_802, n_807, n_808, n_809, n_810, n_815;
  wire n_816, n_817, n_818, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_831, n_832, n_833, n_834, n_835, n_836;
  wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868;
  wire n_869, n_870, n_875, n_876, n_877, n_878, n_879, n_880;
  wire n_881, n_883, n_884, n_885, n_886, n_891, n_892, n_893;
  wire n_894, n_899, n_900, n_901, n_902, n_907, n_908, n_909;
  wire n_910, n_911, n_916, n_917, n_918, n_919, n_922, n_923;
  wire n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931;
  wire n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939;
  wire n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947;
  wire n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955;
  wire n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963;
  wire n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971;
  wire n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979;
  wire n_980, n_985, n_986, n_987, n_988, n_989, n_990, n_991;
  wire n_993, n_994, n_995, n_996, n_1001, n_1002, n_1003, n_1004;
  wire n_1009, n_1010, n_1011, n_1012, n_1017, n_1018, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1044;
  wire n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052;
  wire n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060;
  wire n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068;
  wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1077, n_1078, n_1079, n_1080, n_1085, n_1086, n_1087, n_1088;
  wire n_1093, n_1094, n_1095, n_1096, n_1101, n_1102, n_1103, n_1104;
  wire n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1117;
  wire n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125;
  wire n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1137;
  wire n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153;
  wire n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161;
  wire n_1162, n_1163, n_1164, n_1169, n_1170, n_1171, n_1172, n_1173;
  wire n_1174, n_1175, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182;
  wire n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1193, n_1194;
  wire n_1195, n_1196, n_1197, n_1202, n_1203, n_1204, n_1205, n_1206;
  wire n_1211, n_1212, n_1213, n_1214, n_1217, n_1218, n_1219, n_1220;
  wire n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228;
  wire n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236;
  wire n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244;
  wire n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264;
  wire n_1265, n_1266, n_1267, n_1272, n_1273, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1304, n_1305;
  wire n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313;
  wire n_1314, n_1315, n_1320, n_1321, n_1322, n_1323, n_1328, n_1329;
  wire n_1330, n_1331, n_1336, n_1337, n_1338, n_1339, n_1340, n_1345;
  wire n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377;
  wire n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385;
  wire n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393;
  wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
  wire n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1413;
  wire n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1421, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430;
  wire n_1431, n_1432, n_1433, n_1438, n_1439, n_1440, n_1441, n_1446;
  wire n_1447, n_1448, n_1449, n_1454, n_1455, n_1456, n_1457, n_1459;
  wire n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1470, n_1471;
  wire n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1490, n_1491;
  wire n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499;
  wire n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507;
  wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1517, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527;
  wire n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1538, n_1539;
  wire n_1540, n_1541, n_1542, n_1543, n_1544, n_1546, n_1547, n_1548;
  wire n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556;
  wire n_1557, n_1562, n_1563, n_1564, n_1565, n_1566, n_1571, n_1572;
  wire n_1573, n_1574, n_1575, n_1580, n_1581, n_1582, n_1583, n_1586;
  wire n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594;
  wire n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602;
  wire n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610;
  wire n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618;
  wire n_1619, n_1620, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630;
  wire n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1641, n_1642;
  wire n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650;
  wire n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658;
  wire n_1659, n_1660, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670;
  wire n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1681, n_1682;
  wire n_1683, n_1684, n_1685, n_1686, n_1687, n_1689, n_1690, n_1691;
  wire n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699;
  wire n_1700, n_1705, n_1706, n_1707, n_1708, n_1713, n_1714, n_1715;
  wire n_1716, n_1721, n_1722, n_1723, n_1724, n_1725, n_1730, n_1731;
  wire n_1732, n_1733, n_1734, n_1735, n_1736, n_1741, n_1742, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763;
  wire n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771;
  wire n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779;
  wire n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787;
  wire n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1810, n_1815, n_1816, n_1817, n_1818, n_1819;
  wire n_1820, n_1821, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1839, n_1840;
  wire n_1841, n_1842, n_1847, n_1848, n_1849, n_1850, n_1855, n_1856;
  wire n_1857, n_1858, n_1863, n_1864, n_1865, n_1866, n_1868, n_1869;
  wire n_1870, n_1871, n_1872, n_1873, n_1874, n_1879, n_1880, n_1881;
  wire n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889;
  wire n_1890, n_1891, n_1892, n_1893, n_1894, n_1899, n_1900, n_1901;
  wire n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909;
  wire n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917;
  wire n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925;
  wire n_1926, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937;
  wire n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945;
  wire n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1956, n_1957;
  wire n_1958, n_1959, n_1960, n_1961, n_1962, n_1964, n_1965, n_1966;
  wire n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974;
  wire n_1975, n_1976, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986;
  wire n_1987, n_1989, n_1990, n_1991, n_1992, n_1997, n_1998, n_1999;
  wire n_2000, n_2001, n_2006, n_2007, n_2008, n_2009, n_2010, n_2015;
  wire n_2016, n_2017, n_2018, n_2021, n_2022, n_2023, n_2024, n_2025;
  wire n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033;
  wire n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041;
  wire n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049;
  wire n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2060, n_2061;
  wire n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069;
  wire n_2070, n_2071, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081;
  wire n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089;
  wire n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2100, n_2101;
  wire n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109;
  wire n_2110, n_2111, n_2112, n_2117, n_2118, n_2119, n_2120, n_2121;
  wire n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129;
  wire n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137;
  wire n_2142, n_2143, n_2144, n_2145, n_2150, n_2151, n_2152, n_2153;
  wire n_2154, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165;
  wire n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177;
  wire n_2178, n_2179, n_2180, n_2181, n_2186, n_2187, n_2188, n_2189;
  wire n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197;
  wire n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205;
  wire n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213;
  wire n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225;
  wire n_2226, n_2227, n_2228, n_2229, n_2234, n_2235, n_2236, n_2237;
  wire n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245;
  wire n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257;
  wire n_2258, n_2259, n_2260, n_2261, n_2266, n_2267, n_2268, n_2269;
  wire n_2270, n_2271, n_2272, n_2274, n_2275, n_2276, n_2277, n_2278;
  wire n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2290;
  wire n_2291, n_2292, n_2293, n_2298, n_2299, n_2300, n_2301, n_2306;
  wire n_2307, n_2308, n_2309, n_2314, n_2315, n_2316, n_2317, n_2319;
  wire n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2330, n_2331;
  wire n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339;
  wire n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2350, n_2351;
  wire n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359;
  wire n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367;
  wire n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375;
  wire n_2376, n_2377, n_2378, n_2383, n_2384, n_2385, n_2386, n_2387;
  wire n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2399;
  wire n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407;
  wire n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415;
  wire n_2416, n_2417, n_2418, n_2419, n_2424, n_2425, n_2426, n_2427;
  wire n_2428, n_2429, n_2430, n_2432, n_2433, n_2434, n_2435, n_2436;
  wire n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2448;
  wire n_2449, n_2450, n_2451, n_2452, n_2457, n_2458, n_2459, n_2460;
  wire n_2461, n_2466, n_2467, n_2468, n_2469, n_2472, n_2473, n_2474;
  wire n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482;
  wire n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490;
  wire n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498;
  wire n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506;
  wire n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518;
  wire n_2519, n_2520, n_2521, n_2522, n_2527, n_2528, n_2529, n_2530;
  wire n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538;
  wire n_2539, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550;
  wire n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2561, n_2562;
  wire n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, n_2570;
  wire n_2571, n_2572, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582;
  wire n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590;
  wire n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2601, n_2602;
  wire n_2603, n_2604, n_2605, n_2606, n_2607, n_2609, n_2610, n_2611;
  wire n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619;
  wire n_2620, n_2625, n_2626, n_2627, n_2628, n_2633, n_2634, n_2635;
  wire n_2636, n_2641, n_2642, n_2643, n_2644, n_2645, n_2650, n_2651;
  wire n_2652, n_2653, n_2654, n_2655, n_2656, n_2661, n_2662, n_2663;
  wire n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671;
  wire n_2672, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683;
  wire n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691;
  wire n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699;
  wire n_2700, n_2701, n_2702, n_2703, n_2704, n_2709, n_2710, n_2711;
  wire n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719;
  wire n_2720, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731;
  wire n_2732, n_2733, n_2734, n_2735, n_2736, n_2741, n_2742, n_2743;
  wire n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751;
  wire n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759;
  wire n_2760, n_2761, n_2762, n_2767, n_2768, n_2769, n_2770, n_2771;
  wire n_2772, n_2773, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780;
  wire n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2792;
  wire n_2793, n_2794, n_2795, n_2800, n_2801, n_2802, n_2803, n_2808;
  wire n_2809, n_2810, n_2811, n_2813, n_2814, n_2815, n_2816, n_2817;
  wire n_2818, n_2819, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829;
  wire n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837;
  wire n_2838, n_2839, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849;
  wire n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857;
  wire n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865;
  wire n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2876, n_2877;
  wire n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885;
  wire n_2886, n_2887, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897;
  wire n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2908, n_2909;
  wire n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917;
  wire n_2918, n_2919, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929;
  wire n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2940, n_2941;
  wire n_2942, n_2943, n_2944, n_2945, n_2946, n_2948, n_2949, n_2950;
  wire n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958;
  wire n_2959, n_2964, n_2965, n_2966, n_2967, n_2968, n_2973, n_2974;
  wire n_2975, n_2976, n_2977, n_2982, n_2983, n_2984, n_2985, n_2988;
  wire n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996;
  wire n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004;
  wire n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012;
  wire n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020;
  wire n_3021, n_3022, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032;
  wire n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3043, n_3044;
  wire n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052;
  wire n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060;
  wire n_3061, n_3062, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072;
  wire n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3083, n_3084;
  wire n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092;
  wire n_3093, n_3094, n_3095, n_3100, n_3101, n_3102, n_3103, n_3104;
  wire n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3116;
  wire n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124;
  wire n_3125, n_3126, n_3127, n_3132, n_3133, n_3134, n_3135, n_3136;
  wire n_3137, n_3138, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145;
  wire n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3156, n_3157;
  wire n_3158, n_3159, n_3164, n_3165, n_3166, n_3167, n_3168, n_3173;
  wire n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3184, n_3185;
  wire n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193;
  wire n_3194, n_3195, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205;
  wire n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3217;
  wire n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225;
  wire n_3226, n_3227, n_3228, n_3233, n_3234, n_3235, n_3236, n_3237;
  wire n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245;
  wire n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3257;
  wire n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265;
  wire n_3266, n_3267, n_3268, n_3273, n_3274, n_3275, n_3276, n_3277;
  wire n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285;
  wire n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3297;
  wire n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305;
  wire n_3306, n_3307, n_3308, n_3313, n_3314, n_3315, n_3316, n_3317;
  wire n_3318, n_3319, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326;
  wire n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3338;
  wire n_3339, n_3340, n_3341, n_3346, n_3347, n_3348, n_3349, n_3354;
  wire n_3355, n_3356, n_3357, n_3359, n_3360, n_3361, n_3362, n_3363;
  wire n_3364, n_3365, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375;
  wire n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383;
  wire n_3384, n_3385, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395;
  wire n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3406, n_3407;
  wire n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415;
  wire n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423;
  wire n_3424, n_3425, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435;
  wire n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3446, n_3447;
  wire n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455;
  wire n_3456, n_3457, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467;
  wire n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475;
  wire n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3486, n_3487;
  wire n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495;
  wire n_3496, n_3497, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507;
  wire n_3508, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516;
  wire n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3527, n_3528;
  wire n_3529, n_3530, n_3531, n_3536, n_3537, n_3538, n_3539, n_3540;
  wire n_3545, n_3546, n_3547, n_3548, n_3551, n_3552, n_3553, n_3554;
  wire n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562;
  wire n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570;
  wire n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578;
  wire n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586;
  wire n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3598;
  wire n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606;
  wire n_3607, n_3608, n_3609, n_3614, n_3615, n_3616, n_3617, n_3618;
  wire n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626;
  wire n_3627, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638;
  wire n_3639, n_3640, n_3641, n_3642, n_3643, n_3648, n_3649, n_3650;
  wire n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658;
  wire n_3659, n_3660, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670;
  wire n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3681, n_3682;
  wire n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690;
  wire n_3691, n_3692, n_3693, n_3698, n_3699, n_3700, n_3701, n_3702;
  wire n_3703, n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3714;
  wire n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3722, n_3723;
  wire n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731;
  wire n_3732, n_3733, n_3734, n_3739, n_3740, n_3741, n_3742, n_3747;
  wire n_3748, n_3749, n_3750, n_3755, n_3756, n_3757, n_3758, n_3763;
  wire n_3764, n_3765, n_3766, n_3771, n_3772, n_3773, n_3774, n_3775;
  wire n_3776, n_3777, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787;
  wire n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3798, n_3799;
  wire n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3807;
  wire n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815;
  wire n_3816, n_3817, n_3818, n_3819, n_3824, n_3825, n_3826, n_3827;
  wire n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835;
  wire n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, n_3843;
  wire n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855;
  wire n_3856, n_3857, n_3858, n_3859, n_3864, n_3865, n_3866, n_3867;
  wire n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875;
  wire n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883;
  wire n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, n_3890, n_3891;
  wire n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903;
  wire n_3904, n_3905, n_3906, n_3907, n_3912, n_3913, n_3914, n_3915;
  wire n_3916, n_3917, n_3918, n_3920, n_3921, n_3922, n_3923, n_3924;
  wire n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, n_3931, n_3936;
  wire n_3937, n_3938, n_3939, n_3944, n_3945, n_3946, n_3947, n_3952;
  wire n_3953, n_3954, n_3955, n_3960, n_3961, n_3962, n_3963, n_3965;
  wire n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3976, n_3977;
  wire n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985;
  wire n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3996, n_3997;
  wire n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005;
  wire n_4006, n_4007, n_4012, n_4013, n_4014, n_4015, n_4016, n_4017;
  wire n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024, n_4025;
  wire n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4036, n_4037;
  wire n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045;
  wire n_4046, n_4047, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057;
  wire n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4068, n_4069;
  wire n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077;
  wire n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085;
  wire n_4086, n_4087, n_4092, n_4093, n_4094, n_4095, n_4096, n_4097;
  wire n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, n_4105;
  wire n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4116, n_4117;
  wire n_4118, n_4119, n_4120, n_4121, n_4122, n_4124, n_4125, n_4126;
  wire n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134;
  wire n_4135, n_4136, n_4141, n_4142, n_4143, n_4144, n_4149, n_4150;
  wire n_4151, n_4152, n_4153, n_4158, n_4159, n_4160, n_4161, n_4166;
  wire n_4167, n_4168, n_4169, n_4174, n_4175, n_4176, n_4177, n_4178;
  wire n_4183, n_4184, n_4185, n_4186, n_4187, n_4192, n_4193, n_4194;
  wire n_4195, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204;
  wire n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212;
  wire n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220;
  wire n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, n_4228;
  wire n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236;
  wire n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244;
  wire n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252;
  wire n_4253, n_4254, n_4255, n_4256, n_4257, n_4262, n_4263, n_4264;
  wire n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272;
  wire n_4273, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284;
  wire n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4295, n_4296;
  wire n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, n_4304;
  wire n_4305, n_4306, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316;
  wire n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324;
  wire n_4325, n_4326, n_4327, n_4328, n_4329, n_4330, n_4331, n_4332;
  wire n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4343, n_4344;
  wire n_4345, n_4346, n_4347, n_4348, n_4349, n_4351, n_4352, n_4353;
  wire n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360, n_4361;
  wire n_4362, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373;
  wire n_4375, n_4376, n_4377, n_4378, n_4383, n_4384, n_4385, n_4386;
  wire n_4391, n_4392, n_4393, n_4394, n_4399, n_4400, n_4401, n_4402;
  wire n_4407, n_4408, n_4409, n_4410, n_4415, n_4416, n_4417, n_4418;
  wire n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4434;
  wire n_4435, n_4436, n_4437, n_4438, n_4439, n_4440, n_4441, n_4442;
  wire n_4443, n_4444, n_4445, n_4450, n_4451, n_4452, n_4453, n_4454;
  wire n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462;
  wire n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470;
  wire n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481, n_4482;
  wire n_4483, n_4484, n_4485, n_4486, n_4487, n_4488, n_4489, n_4490;
  wire n_4491, n_4492, n_4493, n_4494, n_4499, n_4500, n_4501, n_4502;
  wire n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509, n_4510;
  wire n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521, n_4522;
  wire n_4523, n_4524, n_4525, n_4526, n_4531, n_4532, n_4533, n_4534;
  wire n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542;
  wire n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4550;
  wire n_4551, n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558;
  wire n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565, n_4566;
  wire n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574;
  wire n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, n_4585, n_4587;
  wire n_4588, n_4589, n_4590, n_4595, n_4596, n_4597, n_4598, n_4603;
  wire n_4604, n_4605, n_4606, n_4611, n_4612, n_4613, n_4614, n_4619;
  wire n_4620, n_4621, n_4622, n_4624, n_4625, n_4626, n_4627, n_4628;
  wire n_4629, n_4630, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640;
  wire n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648;
  wire n_4649, n_4650, n_4651, n_4656, n_4657, n_4658, n_4659, n_4660;
  wire n_4661, n_4662, n_4663, n_4664, n_4665, n_4666, n_4667, n_4672;
  wire n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680;
  wire n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688;
  wire n_4689, n_4690, n_4691, n_4696, n_4697, n_4698, n_4699, n_4700;
  wire n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, n_4712;
  wire n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720;
  wire n_4721, n_4722, n_4723, n_4728, n_4729, n_4730, n_4731, n_4732;
  wire n_4733, n_4734, n_4735, n_4736, n_4737, n_4738, n_4739, n_4740;
  wire n_4741, n_4742, n_4743, n_4744, n_4745, n_4746, n_4747, n_4752;
  wire n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760;
  wire n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768;
  wire n_4769, n_4770, n_4771, n_4776, n_4777, n_4778, n_4779, n_4780;
  wire n_4781, n_4782, n_4783, n_4784, n_4785, n_4786, n_4787, n_4788;
  wire n_4789, n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4800;
  wire n_4801, n_4802, n_4803, n_4804, n_4809, n_4810, n_4811, n_4812;
  wire n_4813, n_4818, n_4819, n_4820, n_4821, n_4826, n_4827, n_4828;
  wire n_4829, n_4834, n_4835, n_4836, n_4837, n_4838, n_4843, n_4844;
  wire n_4845, n_4846, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854;
  wire n_4855, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862;
  wire n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870;
  wire n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877, n_4878;
  wire n_4879, n_4880, n_4881, n_4882, n_4883, n_4888, n_4889, n_4890;
  wire n_4891, n_4892, n_4893, n_4894, n_4895, n_4896, n_4897, n_4898;
  wire n_4899, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4910;
  wire n_4911, n_4912, n_4913, n_4914, n_4915, n_4916, n_4917, n_4918;
  wire n_4919, n_4920, n_4921, n_4922, n_4923, n_4924, n_4929, n_4930;
  wire n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938;
  wire n_4939, n_4940, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950;
  wire n_4951, n_4952, n_4953, n_4954, n_4955, n_4956, n_4961, n_4962;
  wire n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970;
  wire n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978;
  wire n_4979, n_4980, n_4981, n_4986, n_4987, n_4988, n_4989, n_4990;
  wire n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997, n_4998;
  wire n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, n_5005, n_5006;
  wire n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, n_5018;
  wire n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5026, n_5027;
  wire n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035;
  wire n_5036, n_5037, n_5038, n_5043, n_5044, n_5045, n_5046, n_5051;
  wire n_5052, n_5053, n_5054, n_5059, n_5060, n_5061, n_5062, n_5067;
  wire n_5068, n_5069, n_5070, n_5075, n_5076, n_5077, n_5078, n_5083;
  wire n_5084, n_5085, n_5086, n_5091, n_5092, n_5093, n_5094, n_5099;
  wire n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5110, n_5111;
  wire n_5112, n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119;
  wire n_5120, n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127;
  wire n_5128, n_5129, n_5130, n_5135, n_5136, n_5137, n_5138, n_5139;
  wire n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147;
  wire n_5148, n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155;
  wire n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163;
  wire n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5175;
  wire n_5176, n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183;
  wire n_5184, n_5185, n_5186, n_5191, n_5192, n_5193, n_5194, n_5195;
  wire n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203;
  wire n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211;
  wire n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219;
  wire n_5220, n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5231;
  wire n_5232, n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239;
  wire n_5240, n_5241, n_5242, n_5247, n_5248, n_5249, n_5250, n_5251;
  wire n_5252, n_5253, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260;
  wire n_5261, n_5262, n_5263, n_5264, n_5265, n_5266, n_5271, n_5272;
  wire n_5273, n_5274, n_5275, n_5280, n_5281, n_5282, n_5283, n_5288;
  wire n_5289, n_5290, n_5291, n_5296, n_5297, n_5298, n_5299, n_5304;
  wire n_5305, n_5306, n_5307, n_5312, n_5313, n_5314, n_5315, n_5317;
  wire n_5318, n_5319, n_5320, n_5321, n_5322, n_5323, n_5328, n_5329;
  wire n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336, n_5337;
  wire n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5348, n_5349;
  wire n_5350, n_5351, n_5352, n_5353, n_5354, n_5355, n_5356, n_5357;
  wire n_5358, n_5359, n_5360, n_5361, n_5362, n_5363, n_5364, n_5365;
  wire n_5366, n_5367, n_5368, n_5373, n_5374, n_5375, n_5376, n_5377;
  wire n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384, n_5385;
  wire n_5390, n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397;
  wire n_5398, n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405;
  wire n_5406, n_5407, n_5408, n_5409, n_5414, n_5415, n_5416, n_5417;
  wire n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424, n_5425;
  wire n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432, n_5433;
  wire n_5438, n_5439, n_5440, n_5441, n_5442, n_5443, n_5444, n_5445;
  wire n_5446, n_5447, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453;
  wire n_5454, n_5455, n_5456, n_5457, n_5462, n_5463, n_5464, n_5465;
  wire n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472, n_5473;
  wire n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480, n_5481;
  wire n_5482, n_5487, n_5488, n_5489, n_5490, n_5491, n_5492, n_5493;
  wire n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5501, n_5502;
  wire n_5503, n_5504, n_5505, n_5506, n_5507, n_5512, n_5513, n_5514;
  wire n_5515, n_5516, n_5517, n_5518, n_5520, n_5521, n_5522, n_5523;
  wire n_5528, n_5529, n_5530, n_5531, n_5532, n_5537, n_5538, n_5539;
  wire n_5540, n_5545, n_5546, n_5547, n_5548, n_5553, n_5554, n_5555;
  wire n_5556, n_5557, n_5562, n_5563, n_5564, n_5565, n_5568, n_5569;
  wire n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576, n_5577;
  wire n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584, n_5585;
  wire n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592, n_5593;
  wire n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600, n_5601;
  wire n_5602, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613;
  wire n_5614, n_5615, n_5616, n_5617, n_5618, n_5623, n_5624, n_5625;
  wire n_5626, n_5627, n_5628, n_5629, n_5630, n_5631, n_5632, n_5633;
  wire n_5634, n_5635, n_5636, n_5637, n_5638, n_5639, n_5640, n_5641;
  wire n_5642, n_5643, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653;
  wire n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5664, n_5665;
  wire n_5666, n_5667, n_5668, n_5669, n_5670, n_5671, n_5672, n_5673;
  wire n_5674, n_5675, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685;
  wire n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693;
  wire n_5694, n_5695, n_5696, n_5697, n_5698, n_5699, n_5700, n_5705;
  wire n_5706, n_5707, n_5708, n_5709, n_5710, n_5711, n_5712, n_5713;
  wire n_5714, n_5715, n_5716, n_5717, n_5718, n_5719, n_5720, n_5721;
  wire n_5722, n_5723, n_5724, n_5725, n_5730, n_5731, n_5732, n_5733;
  wire n_5734, n_5735, n_5736, n_5737, n_5738, n_5739, n_5740, n_5741;
  wire n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, n_5752, n_5753;
  wire n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760, n_5761;
  wire n_5762, n_5763, n_5764, n_5765, n_5770, n_5771, n_5772, n_5773;
  wire n_5778, n_5779, n_5780, n_5781, n_5786, n_5787, n_5788, n_5789;
  wire n_5794, n_5795, n_5796, n_5797, n_5802, n_5803, n_5804, n_5805;
  wire n_5810, n_5811, n_5812, n_5813, n_5818, n_5819, n_5820, n_5821;
  wire n_5826, n_5827, n_5828, n_5829, n_5834, n_5835, n_5836, n_5837;
  wire n_5838, n_5839, n_5840, n_5845, n_5846, n_5847, n_5848, n_5849;
  wire n_5850, n_5851, n_5852, n_5853, n_5854, n_5855, n_5856, n_5857;
  wire n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5864, n_5865;
  wire n_5870, n_5871, n_5872, n_5873, n_5874, n_5875, n_5876, n_5877;
  wire n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884, n_5885;
  wire n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892, n_5893;
  wire n_5894, n_5895, n_5896, n_5897, n_5898, n_5899, n_5900, n_5901;
  wire n_5902, n_5903, n_5904, n_5905, n_5910, n_5911, n_5912, n_5913;
  wire n_5914, n_5915, n_5916, n_5917, n_5918, n_5919, n_5920, n_5921;
  wire n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932, n_5933;
  wire n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940, n_5941;
  wire n_5942, n_5943, n_5944, n_5945, n_5946, n_5947, n_5948, n_5949;
  wire n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956, n_5957;
  wire n_5958, n_5959, n_5960, n_5961, n_5966, n_5967, n_5968, n_5969;
  wire n_5970, n_5971, n_5972, n_5973, n_5974, n_5975, n_5976, n_5977;
  wire n_5978, n_5979, n_5980, n_5981, n_5982, n_5983, n_5984, n_5985;
  wire n_5986, n_5991, n_5992, n_5993, n_5994, n_5995, n_5996, n_5997;
  wire n_5999, n_6000, n_6001, n_6002, n_6003, n_6004, n_6005, n_6006;
  wire n_6007, n_6008, n_6009, n_6010, n_6011, n_6016, n_6017, n_6018;
  wire n_6019, n_6024, n_6025, n_6026, n_6027, n_6032, n_6033, n_6034;
  wire n_6035, n_6040, n_6041, n_6042, n_6043, n_6048, n_6049, n_6050;
  wire n_6051, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059;
  wire n_6064, n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071;
  wire n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079;
  wire n_6084, n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091;
  wire n_6092, n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099;
  wire n_6100, n_6101, n_6102, n_6103, n_6104, n_6109, n_6110, n_6111;
  wire n_6112, n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119;
  wire n_6120, n_6121, n_6126, n_6127, n_6128, n_6129, n_6130, n_6131;
  wire n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6139;
  wire n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6150, n_6151;
  wire n_6152, n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6159;
  wire n_6160, n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167;
  wire n_6168, n_6169, n_6174, n_6175, n_6176, n_6177, n_6178, n_6179;
  wire n_6180, n_6181, n_6182, n_6183, n_6184, n_6185, n_6186, n_6187;
  wire n_6188, n_6189, n_6190, n_6191, n_6192, n_6193, n_6198, n_6199;
  wire n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207;
  wire n_6208, n_6209, n_6214, n_6215, n_6216, n_6217, n_6218, n_6219;
  wire n_6220, n_6221, n_6222, n_6223, n_6224, n_6225, n_6230, n_6231;
  wire n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239;
  wire n_6240, n_6241, n_6246, n_6247, n_6248, n_6249, n_6250, n_6251;
  wire n_6252, n_6254, n_6255, n_6256, n_6257, n_6258, n_6259, n_6260;
  wire n_6261, n_6262, n_6263, n_6264, n_6265, n_6270, n_6271, n_6272;
  wire n_6273, n_6274, n_6279, n_6280, n_6281, n_6282, n_6287, n_6288;
  wire n_6289, n_6290, n_6295, n_6296, n_6297, n_6298, n_6299, n_6304;
  wire n_6305, n_6306, n_6307, n_6310, n_6311, n_6312, n_6313, n_6314;
  wire n_6315, n_6316, n_6317, n_6318, n_6319, n_6320, n_6321, n_6322;
  wire n_6323, n_6324, n_6325, n_6326, n_6327, n_6328, n_6329, n_6330;
  wire n_6331, n_6332, n_6333, n_6334, n_6335, n_6336, n_6337, n_6338;
  wire n_6339, n_6340, n_6341, n_6342, n_6343, n_6344, n_6349, n_6350;
  wire n_6351, n_6352, n_6353, n_6354, n_6355, n_6356, n_6357, n_6358;
  wire n_6359, n_6360, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370;
  wire n_6371, n_6372, n_6373, n_6374, n_6375, n_6376, n_6377, n_6378;
  wire n_6379, n_6380, n_6381, n_6382, n_6383, n_6384, n_6385, n_6390;
  wire n_6391, n_6392, n_6393, n_6394, n_6395, n_6396, n_6397, n_6398;
  wire n_6399, n_6400, n_6401, n_6406, n_6407, n_6408, n_6409, n_6410;
  wire n_6411, n_6412, n_6413, n_6414, n_6415, n_6416, n_6417, n_6422;
  wire n_6423, n_6424, n_6425, n_6426, n_6427, n_6428, n_6429, n_6430;
  wire n_6431, n_6432, n_6433, n_6434, n_6435, n_6436, n_6437, n_6438;
  wire n_6439, n_6440, n_6441, n_6442, n_6447, n_6448, n_6449, n_6450;
  wire n_6451, n_6452, n_6453, n_6454, n_6455, n_6456, n_6457, n_6458;
  wire n_6459, n_6460, n_6461, n_6462, n_6463, n_6464, n_6465, n_6466;
  wire n_6467, n_6472, n_6473, n_6474, n_6475, n_6476, n_6477, n_6478;
  wire n_6479, n_6480, n_6481, n_6482, n_6483, n_6488, n_6489, n_6490;
  wire n_6491, n_6492, n_6493, n_6494, n_6495, n_6496, n_6497, n_6498;
  wire n_6499, n_6504, n_6505, n_6506, n_6507, n_6508, n_6509, n_6510;
  wire n_6511, n_6512, n_6513, n_6514, n_6515, n_6516, n_6521, n_6522;
  wire n_6523, n_6524, n_6525, n_6526, n_6527, n_6529, n_6530, n_6531;
  wire n_6532, n_6533, n_6534, n_6535, n_6536, n_6537, n_6538, n_6539;
  wire n_6540, n_6545, n_6546, n_6547, n_6548, n_6549, n_6550, n_6551;
  wire n_6553, n_6554, n_6555, n_6556, n_6561, n_6562, n_6563, n_6564;
  wire n_6569, n_6570, n_6571, n_6572, n_6577, n_6578, n_6579, n_6580;
  wire n_6585, n_6586, n_6587, n_6588, n_6593, n_6594, n_6595, n_6596;
  wire n_6601, n_6602, n_6603, n_6604, n_6609, n_6610, n_6611, n_6612;
  wire n_6613, n_6614, n_6615, n_6620, n_6621, n_6622, n_6623, n_6624;
  wire n_6625, n_6626, n_6627, n_6628, n_6629, n_6630, n_6631, n_6632;
  wire n_6633, n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640;
  wire n_6645, n_6646, n_6647, n_6648, n_6649, n_6650, n_6651, n_6652;
  wire n_6653, n_6654, n_6655, n_6656, n_6657, n_6658, n_6659, n_6660;
  wire n_6661, n_6662, n_6663, n_6664, n_6665, n_6666, n_6667, n_6668;
  wire n_6669, n_6670, n_6671, n_6672, n_6673, n_6678, n_6679, n_6680;
  wire n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687, n_6688;
  wire n_6689, n_6690, n_6695, n_6696, n_6697, n_6698, n_6699, n_6700;
  wire n_6701, n_6702, n_6703, n_6704, n_6705, n_6706, n_6711, n_6712;
  wire n_6713, n_6714, n_6715, n_6716, n_6717, n_6718, n_6719, n_6720;
  wire n_6721, n_6722, n_6723, n_6724, n_6725, n_6726, n_6727, n_6728;
  wire n_6729, n_6730, n_6731, n_6732, n_6733, n_6734, n_6735, n_6736;
  wire n_6737, n_6738, n_6739, n_6740, n_6741, n_6742, n_6743, n_6744;
  wire n_6745, n_6746, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756;
  wire n_6757, n_6758, n_6759, n_6760, n_6761, n_6762, n_6767, n_6768;
  wire n_6769, n_6770, n_6771, n_6772, n_6773, n_6774, n_6775, n_6776;
  wire n_6777, n_6778, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788;
  wire n_6789, n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796;
  wire n_6797, n_6798, n_6799, n_6800, n_6801, n_6802, n_6807, n_6808;
  wire n_6809, n_6810, n_6811, n_6812, n_6813, n_6815, n_6816, n_6817;
  wire n_6818, n_6823, n_6824, n_6825, n_6826, n_6831, n_6832, n_6833;
  wire n_6834, n_6839, n_6840, n_6841, n_6842, n_6847, n_6848, n_6849;
  wire n_6850, n_6855, n_6856, n_6857, n_6858, n_6860, n_6861, n_6862;
  wire n_6863, n_6864, n_6865, n_6866, n_6871, n_6872, n_6873, n_6874;
  wire n_6875, n_6876, n_6877, n_6878, n_6879, n_6880, n_6881, n_6882;
  wire n_6883, n_6884, n_6885, n_6886, n_6891, n_6892, n_6893, n_6894;
  wire n_6895, n_6896, n_6897, n_6898, n_6899, n_6900, n_6901, n_6902;
  wire n_6903, n_6904, n_6905, n_6906, n_6907, n_6908, n_6909, n_6910;
  wire n_6911, n_6912, n_6913, n_6914, n_6915, n_6916, n_6917, n_6918;
  wire n_6923, n_6924, n_6925, n_6926, n_6927, n_6928, n_6929, n_6930;
  wire n_6931, n_6932, n_6933, n_6934, n_6939, n_6940, n_6941, n_6942;
  wire n_6943, n_6944, n_6945, n_6946, n_6947, n_6948, n_6949, n_6950;
  wire n_6955, n_6956, n_6957, n_6958, n_6959, n_6960, n_6961, n_6962;
  wire n_6963, n_6964, n_6965, n_6966, n_6967, n_6968, n_6969, n_6970;
  wire n_6971, n_6972, n_6973, n_6974, n_6979, n_6980, n_6981, n_6982;
  wire n_6983, n_6984, n_6985, n_6986, n_6987, n_6988, n_6989, n_6990;
  wire n_6991, n_6992, n_6993, n_6994, n_6995, n_6996, n_6997, n_6998;
  wire n_7003, n_7004, n_7005, n_7006, n_7007, n_7008, n_7009, n_7010;
  wire n_7011, n_7012, n_7013, n_7014, n_7019, n_7020, n_7021, n_7022;
  wire n_7023, n_7024, n_7025, n_7026, n_7027, n_7028, n_7029, n_7030;
  wire n_7035, n_7036, n_7037, n_7038, n_7039, n_7040, n_7041, n_7042;
  wire n_7043, n_7044, n_7045, n_7046, n_7051, n_7052, n_7053, n_7054;
  wire n_7055, n_7056, n_7057, n_7058, n_7059, n_7060, n_7061, n_7062;
  wire n_7063, n_7064, n_7065, n_7066, n_7067, n_7068, n_7069, n_7070;
  wire n_7071, n_7076, n_7077, n_7078, n_7079, n_7084, n_7085, n_7086;
  wire n_7087, n_7092, n_7093, n_7094, n_7095, n_7096, n_7101, n_7102;
  wire n_7103, n_7104, n_7107, n_7108, n_7109, n_7110, n_7111, n_7112;
  wire n_7113, n_7114, n_7115, n_7116, n_7117, n_7118, n_7119, n_7120;
  wire n_7121, n_7122, n_7123, n_7124, n_7125, n_7126, n_7127, n_7128;
  wire n_7129, n_7130, n_7131, n_7132, n_7133, n_7134, n_7135, n_7136;
  wire n_7137, n_7138, n_7139, n_7140, n_7141, n_7146, n_7147, n_7148;
  wire n_7149, n_7150, n_7151, n_7152, n_7153, n_7154, n_7155, n_7156;
  wire n_7157, n_7162, n_7163, n_7164, n_7165, n_7166, n_7167, n_7168;
  wire n_7169, n_7170, n_7171, n_7172, n_7173, n_7174, n_7175, n_7176;
  wire n_7177, n_7178, n_7179, n_7180, n_7181, n_7186, n_7187, n_7188;
  wire n_7189, n_7190, n_7191, n_7192, n_7193, n_7194, n_7195, n_7196;
  wire n_7197, n_7202, n_7203, n_7204, n_7205, n_7206, n_7207, n_7208;
  wire n_7209, n_7210, n_7211, n_7212, n_7213, n_7218, n_7219, n_7220;
  wire n_7221, n_7222, n_7223, n_7224, n_7225, n_7226, n_7227, n_7228;
  wire n_7229, n_7230, n_7231, n_7232, n_7233, n_7234, n_7235, n_7236;
  wire n_7237, n_7238, n_7243, n_7244, n_7245, n_7246, n_7247, n_7248;
  wire n_7249, n_7250, n_7251, n_7252, n_7253, n_7254, n_7255, n_7260;
  wire n_7261, n_7262, n_7263, n_7264, n_7265, n_7266, n_7267, n_7268;
  wire n_7269, n_7270, n_7271, n_7272, n_7277, n_7278, n_7279, n_7280;
  wire n_7281, n_7282, n_7283, n_7284, n_7285, n_7286, n_7287, n_7288;
  wire n_7293, n_7294, n_7295, n_7296, n_7297, n_7298, n_7299, n_7300;
  wire n_7301, n_7302, n_7303, n_7304, n_7309, n_7310, n_7311, n_7312;
  wire n_7313, n_7314, n_7315, n_7316, n_7317, n_7318, n_7319, n_7320;
  wire n_7321, n_7326, n_7327, n_7328, n_7329, n_7330, n_7331, n_7332;
  wire n_7333, n_7334, n_7335, n_7336, n_7337, n_7342, n_7343, n_7344;
  wire n_7345, n_7346, n_7347, n_7348, n_7350, n_7351, n_7352, n_7353;
  wire n_7354, n_7355, n_7356, n_7357, n_7358, n_7359, n_7360, n_7361;
  wire n_7366, n_7367, n_7368, n_7369, n_7374, n_7375, n_7376, n_7377;
  wire n_7382, n_7383, n_7384, n_7385, n_7390, n_7391, n_7392, n_7393;
  wire n_7398, n_7399, n_7400, n_7401, n_7406, n_7407, n_7408, n_7409;
  wire n_7414, n_7415, n_7416, n_7417, n_7418, n_7419, n_7420, n_7425;
  wire n_7426, n_7427, n_7428, n_7429, n_7430, n_7431, n_7432, n_7433;
  wire n_7434, n_7435, n_7436, n_7437, n_7438, n_7439, n_7440, n_7441;
  wire n_7442, n_7443, n_7444, n_7445, n_7450, n_7451, n_7452, n_7453;
  wire n_7454, n_7455, n_7456, n_7457, n_7458, n_7459, n_7460, n_7461;
  wire n_7462, n_7463, n_7464, n_7465, n_7466, n_7467, n_7468, n_7469;
  wire n_7470, n_7471, n_7472, n_7473, n_7474, n_7475, n_7476, n_7477;
  wire n_7478, n_7483, n_7484, n_7485, n_7486, n_7487, n_7488, n_7489;
  wire n_7490, n_7491, n_7492, n_7493, n_7494, n_7495, n_7500, n_7501;
  wire n_7502, n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509;
  wire n_7510, n_7511, n_7516, n_7517, n_7518, n_7519, n_7520, n_7521;
  wire n_7522, n_7523, n_7524, n_7525, n_7526, n_7527, n_7528, n_7529;
  wire n_7530, n_7531, n_7532, n_7533, n_7534, n_7535, n_7536, n_7537;
  wire n_7538, n_7539, n_7540, n_7541, n_7542, n_7543, n_7544, n_7545;
  wire n_7546, n_7547, n_7548, n_7549, n_7550, n_7551, n_7556, n_7557;
  wire n_7558, n_7559, n_7560, n_7561, n_7562, n_7563, n_7564, n_7565;
  wire n_7566, n_7567, n_7572, n_7573, n_7574, n_7575, n_7576, n_7577;
  wire n_7578, n_7579, n_7580, n_7581, n_7582, n_7583, n_7588, n_7589;
  wire n_7590, n_7591, n_7592, n_7593, n_7594, n_7595, n_7596, n_7597;
  wire n_7598, n_7599, n_7604, n_7605, n_7606, n_7607, n_7608, n_7609;
  wire n_7610, n_7611, n_7612, n_7613, n_7614, n_7615, n_7616, n_7621;
  wire n_7622, n_7623, n_7624, n_7625, n_7626, n_7627, n_7629, n_7630;
  wire n_7631, n_7632, n_7633, n_7634, n_7635, n_7636, n_7637, n_7638;
  wire n_7639, n_7640, n_7645, n_7646, n_7647, n_7648, n_7649, n_7650;
  wire n_7651, n_7653, n_7654, n_7655, n_7656, n_7661, n_7662, n_7663;
  wire n_7664, n_7669, n_7670, n_7671, n_7672, n_7677, n_7678, n_7679;
  wire n_7680, n_7685, n_7686, n_7687, n_7688, n_7693, n_7694, n_7695;
  wire n_7696, n_7701, n_7702, n_7703, n_7704, n_7709, n_7710, n_7711;
  wire n_7712, n_7714, n_7715, n_7716, n_7717, n_7718, n_7719, n_7720;
  wire n_7725, n_7726, n_7727, n_7728, n_7729, n_7730, n_7731, n_7732;
  wire n_7733, n_7734, n_7735, n_7736, n_7737, n_7738, n_7739, n_7740;
  wire n_7745, n_7746, n_7747, n_7748, n_7749, n_7750, n_7751, n_7752;
  wire n_7753, n_7754, n_7755, n_7756, n_7757, n_7758, n_7759, n_7760;
  wire n_7761, n_7762, n_7763, n_7764, n_7765, n_7766, n_7767, n_7768;
  wire n_7769, n_7770, n_7771, n_7772, n_7773, n_7774, n_7775, n_7776;
  wire n_7777, n_7778, n_7779, n_7780, n_7785, n_7786, n_7787, n_7788;
  wire n_7789, n_7790, n_7791, n_7792, n_7793, n_7794, n_7795, n_7796;
  wire n_7801, n_7802, n_7803, n_7804, n_7805, n_7806, n_7807, n_7808;
  wire n_7809, n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816;
  wire n_7817, n_7818, n_7819, n_7820, n_7825, n_7826, n_7827, n_7828;
  wire n_7829, n_7830, n_7831, n_7832, n_7833, n_7834, n_7835, n_7836;
  wire n_7837, n_7838, n_7839, n_7840, n_7841, n_7842, n_7843, n_7844;
  wire n_7849, n_7850, n_7851, n_7852, n_7853, n_7854, n_7855, n_7856;
  wire n_7857, n_7858, n_7859, n_7860, n_7865, n_7866, n_7867, n_7868;
  wire n_7869, n_7870, n_7871, n_7872, n_7873, n_7874, n_7875, n_7876;
  wire n_7881, n_7882, n_7883, n_7884, n_7885, n_7886, n_7887, n_7888;
  wire n_7889, n_7890, n_7891, n_7892, n_7893, n_7894, n_7895, n_7896;
  wire n_7897, n_7898, n_7899, n_7900, n_7905, n_7906, n_7907, n_7908;
  wire n_7909, n_7910, n_7911, n_7912, n_7913, n_7914, n_7915, n_7916;
  wire n_7917, n_7918, n_7919, n_7920, n_7921, n_7922, n_7923, n_7924;
  wire n_7925, n_7930, n_7931, n_7932, n_7933, n_7938, n_7939, n_7940;
  wire n_7941, n_7942, n_7947, n_7948, n_7949, n_7950, n_7953, n_7954;
  wire n_7955, n_7956, n_7957, n_7958, n_7959, n_7960, n_7961, n_7962;
  wire n_7963, n_7964, n_7965, n_7966, n_7967, n_7968, n_7969, n_7970;
  wire n_7971, n_7972, n_7973, n_7974, n_7975, n_7976, n_7977, n_7978;
  wire n_7979, n_7980, n_7981, n_7982, n_7983, n_7984, n_7985, n_7986;
  wire n_7987, n_7992, n_7993, n_7994, n_7995, n_7996, n_7997, n_7998;
  wire n_7999, n_8000, n_8001, n_8002, n_8003, n_8008, n_8009, n_8010;
  wire n_8011, n_8012, n_8013, n_8014, n_8015, n_8016, n_8017, n_8018;
  wire n_8019, n_8020, n_8021, n_8022, n_8023, n_8024, n_8025, n_8026;
  wire n_8027, n_8032, n_8033, n_8034, n_8035, n_8036, n_8037, n_8038;
  wire n_8039, n_8040, n_8041, n_8042, n_8043, n_8048, n_8049, n_8050;
  wire n_8051, n_8052, n_8053, n_8054, n_8055, n_8056, n_8057, n_8058;
  wire n_8059, n_8060, n_8065, n_8066, n_8067, n_8068, n_8069, n_8070;
  wire n_8071, n_8072, n_8073, n_8074, n_8075, n_8076, n_8081, n_8082;
  wire n_8083, n_8084, n_8085, n_8086, n_8087, n_8088, n_8089, n_8090;
  wire n_8091, n_8092, n_8097, n_8098, n_8099, n_8100, n_8101, n_8102;
  wire n_8103, n_8104, n_8105, n_8106, n_8107, n_8108, n_8113, n_8114;
  wire n_8115, n_8116, n_8117, n_8118, n_8119, n_8120, n_8121, n_8122;
  wire n_8123, n_8124, n_8125, n_8130, n_8131, n_8132, n_8133, n_8134;
  wire n_8135, n_8136, n_8137, n_8138, n_8139, n_8140, n_8141, n_8146;
  wire n_8147, n_8148, n_8149, n_8150, n_8151, n_8152, n_8153, n_8154;
  wire n_8155, n_8156, n_8157, n_8162, n_8163, n_8164, n_8165, n_8166;
  wire n_8167, n_8168, n_8169, n_8170, n_8171, n_8172, n_8173, n_8178;
  wire n_8179, n_8180, n_8181, n_8182, n_8183, n_8184, n_8185, n_8186;
  wire n_8187, n_8188, n_8189, n_8190, n_8191, n_8196, n_8197, n_8198;
  wire n_8199, n_8200, n_8201, n_8202, n_8203, n_8204, n_8205, n_8206;
  wire n_8207, n_8212, n_8213, n_8214, n_8215, n_8216, n_8217, n_8218;
  wire n_8220, n_8221, n_8222, n_8223, n_8224, n_8225, n_8226, n_8227;
  wire n_8228, n_8229, n_8230, n_8231, n_8232, n_8237, n_8238, n_8239;
  wire n_8240, n_8245, n_8246, n_8247, n_8248, n_8253, n_8254, n_8255;
  wire n_8256, n_8257, n_8262, n_8263, n_8264, n_8265, n_8270, n_8271;
  wire n_8272, n_8273, n_8278, n_8279, n_8280, n_8281, n_8286, n_8287;
  wire n_8288, n_8289, n_8294, n_8295, n_8296, n_8297, n_8298, n_8299;
  wire n_8300, n_8305, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311;
  wire n_8312, n_8313, n_8314, n_8315, n_8316, n_8321, n_8322, n_8323;
  wire n_8324, n_8325, n_8326, n_8327, n_8328, n_8329, n_8330, n_8331;
  wire n_8332, n_8333, n_8334, n_8335, n_8336, n_8337, n_8338, n_8339;
  wire n_8340, n_8341, n_8342, n_8343, n_8344, n_8345, n_8346, n_8347;
  wire n_8348, n_8349, n_8350, n_8351, n_8352, n_8353, n_8354, n_8355;
  wire n_8356, n_8357, n_8362, n_8363, n_8364, n_8365, n_8366, n_8367;
  wire n_8368, n_8369, n_8370, n_8371, n_8372, n_8373, n_8374, n_8375;
  wire n_8376, n_8377, n_8378, n_8379, n_8380, n_8381, n_8382, n_8383;
  wire n_8388, n_8389, n_8390, n_8391, n_8392, n_8393, n_8394, n_8395;
  wire n_8396, n_8397, n_8398, n_8399, n_8400, n_8401, n_8402, n_8403;
  wire n_8404, n_8405, n_8406, n_8407, n_8408, n_8409, n_8410, n_8411;
  wire n_8412, n_8413, n_8414, n_8415, n_8416, n_8417, n_8418, n_8419;
  wire n_8420, n_8421, n_8422, n_8423, n_8428, n_8429, n_8430, n_8431;
  wire n_8432, n_8433, n_8434, n_8435, n_8436, n_8437, n_8438, n_8439;
  wire n_8444, n_8445, n_8446, n_8447, n_8448, n_8449, n_8450, n_8451;
  wire n_8452, n_8453, n_8454, n_8455, n_8460, n_8461, n_8462, n_8463;
  wire n_8464, n_8465, n_8466, n_8467, n_8468, n_8469, n_8470, n_8471;
  wire n_8476, n_8477, n_8478, n_8479, n_8480, n_8481, n_8482, n_8483;
  wire n_8484, n_8485, n_8486, n_8487, n_8488, n_8493, n_8494, n_8495;
  wire n_8496, n_8497, n_8498, n_8499, n_8500, n_8501, n_8502, n_8503;
  wire n_8504, n_8509, n_8510, n_8511, n_8512, n_8513, n_8514, n_8515;
  wire n_8517, n_8518, n_8519, n_8520, n_8521, n_8522, n_8523, n_8524;
  wire n_8525, n_8526, n_8527, n_8528, n_8529, n_8534, n_8535, n_8536;
  wire n_8537, n_8538, n_8539, n_8540, n_8542, n_8543, n_8544, n_8545;
  wire n_8550, n_8551, n_8552, n_8553, n_8558, n_8559, n_8560, n_8561;
  wire n_8566, n_8567, n_8568, n_8569, n_8574, n_8575, n_8576, n_8577;
  wire n_8582, n_8583, n_8584, n_8585, n_8590, n_8591, n_8592, n_8593;
  wire n_8598, n_8599, n_8600, n_8601, n_8606, n_8607, n_8608, n_8609;
  wire n_8614, n_8615, n_8616, n_8617, n_8622, n_8623, n_8624, n_8625;
  wire n_8627, n_8628, n_8629, n_8630, n_8631, n_8632, n_8633, n_8638;
  wire n_8639, n_8640, n_8641, n_8642, n_8643, n_8644, n_8645, n_8646;
  wire n_8647, n_8648, n_8649, n_8650, n_8651, n_8652, n_8653, n_8654;
  wire n_8655, n_8656, n_8657, n_8658, n_8659, n_8660, n_8661, n_8662;
  wire n_8663, n_8664, n_8665, n_8666, n_8667, n_8668, n_8669, n_8670;
  wire n_8671, n_8672, n_8673, n_8674, n_8675, n_8676, n_8677, n_8678;
  wire n_8679, n_8680, n_8681, n_8682, n_8683, n_8684, n_8685, n_8686;
  wire n_8687, n_8688, n_8689, n_8690, n_8691, n_8692, n_8693, n_8694;
  wire n_8695, n_8696, n_8697, n_8698, n_8699, n_8700, n_8701, n_8702;
  wire n_8703, n_8704, n_8705, n_8706, n_8707, n_8708, n_8709, n_8710;
  wire n_8711, n_8712, n_8713, n_8714, n_8715, n_8716, n_8717, n_8722;
  wire n_8723, n_8724, n_8725, n_8726, n_8727, n_8728, n_8729, n_8730;
  wire n_8731, n_8732, n_8733, n_8738, n_8739, n_8740, n_8741, n_8742;
  wire n_8743, n_8744, n_8745, n_8746, n_8747, n_8748, n_8749, n_8754;
  wire n_8755, n_8756, n_8757, n_8758, n_8759, n_8760, n_8761, n_8762;
  wire n_8763, n_8764, n_8765, n_8770, n_8771, n_8772, n_8773, n_8774;
  wire n_8775, n_8776, n_8777, n_8778, n_8779, n_8780, n_8781, n_8782;
  wire n_8783, n_8784, n_8785, n_8786, n_8787, n_8788, n_8789, n_8790;
  wire n_8795, n_8796, n_8797, n_8798, n_8799, n_8800, n_8801, n_8802;
  wire n_8803, n_8804, n_8805, n_8806, n_8807, n_8812, n_8813, n_8814;
  wire n_8815, n_8816, n_8817, n_8818, n_8819, n_8820, n_8821, n_8822;
  wire n_8823, n_8824, n_8825, n_8826, n_8827, n_8828, n_8829, n_8830;
  wire n_8831, n_8836, n_8837, n_8838, n_8839, n_8844, n_8845, n_8846;
  wire n_8847, n_8852, n_8853, n_8854, n_8855, n_8860, n_8861, n_8862;
  wire n_8863, n_8868, n_8869, n_8870, n_8871, n_8876, n_8877, n_8878;
  wire n_8879, n_8880, n_8885, n_8886, n_8887, n_8888, n_8891, n_8892;
  wire n_8893, n_8894, n_8895, n_8896, n_8897, n_8898, n_8899, n_8900;
  wire n_8901, n_8902, n_8903, n_8904, n_8905, n_8906, n_8907, n_8908;
  wire n_8909, n_8910, n_8911, n_8912, n_8913, n_8914, n_8915, n_8916;
  wire n_8917, n_8918, n_8919, n_8920, n_8921, n_8922, n_8923, n_8924;
  wire n_8925, n_8926, n_8927, n_8928, n_8929, n_8930, n_8931, n_8932;
  wire n_8933, n_8934, n_8935, n_8936, n_8937, n_8938, n_8939, n_8940;
  wire n_8941, n_8942, n_8943, n_8944, n_8945, n_8946, n_8947, n_8948;
  wire n_8949, n_8954, n_8955, n_8956, n_8957, n_8958, n_8959, n_8960;
  wire n_8961, n_8962, n_8963, n_8964, n_8965, n_8970, n_8971, n_8972;
  wire n_8973, n_8974, n_8975, n_8976, n_8977, n_8978, n_8979, n_8980;
  wire n_8981, n_8982, n_8987, n_8988, n_8989, n_8990, n_8991, n_8992;
  wire n_8993, n_8994, n_8995, n_8996, n_8997, n_8998, n_9003, n_9004;
  wire n_9005, n_9006, n_9007, n_9008, n_9009, n_9010, n_9011, n_9012;
  wire n_9013, n_9014, n_9019, n_9020, n_9021, n_9022, n_9023, n_9024;
  wire n_9025, n_9026, n_9027, n_9028, n_9029, n_9030, n_9035, n_9036;
  wire n_9037, n_9038, n_9039, n_9040, n_9041, n_9042, n_9043, n_9044;
  wire n_9045, n_9046, n_9047, n_9052, n_9053, n_9054, n_9055, n_9056;
  wire n_9057, n_9058, n_9059, n_9060, n_9061, n_9062, n_9063, n_9068;
  wire n_9069, n_9070, n_9071, n_9072, n_9073, n_9074, n_9075, n_9076;
  wire n_9077, n_9078, n_9079, n_9084, n_9085, n_9086, n_9087, n_9088;
  wire n_9089, n_9090, n_9091, n_9092, n_9093, n_9094, n_9095, n_9100;
  wire n_9101, n_9102, n_9103, n_9104, n_9105, n_9106, n_9107, n_9108;
  wire n_9109, n_9110, n_9111, n_9112, n_9113, n_9114, n_9115, n_9116;
  wire n_9117, n_9118, n_9119, n_9120, n_9121, n_9122, n_9123, n_9124;
  wire n_9125, n_9126, n_9127, n_9132, n_9133, n_9134, n_9135, n_9136;
  wire n_9137, n_9138, n_9140, n_9141, n_9142, n_9143, n_9144, n_9145;
  wire n_9146, n_9147, n_9148, n_9149, n_9150, n_9151, n_9156, n_9157;
  wire n_9158, n_9159, n_9160, n_9161, n_9162, n_9164, n_9165, n_9166;
  wire n_9167, n_9168, n_9173, n_9174, n_9175, n_9176, n_9181, n_9182;
  wire n_9183, n_9184, n_9189, n_9190, n_9191, n_9192, n_9197, n_9198;
  wire n_9199, n_9200, n_9205, n_9206, n_9207, n_9208, n_9213, n_9214;
  wire n_9215, n_9216, n_9221, n_9222, n_9223, n_9224, n_9225, n_9226;
  wire n_9227, n_9232, n_9233, n_9234, n_9235, n_9236, n_9237, n_9238;
  wire n_9239, n_9240, n_9241, n_9242, n_9243, n_9248, n_9249, n_9250;
  wire n_9251, n_9252, n_9253, n_9254, n_9255, n_9256, n_9257, n_9258;
  wire n_9259, n_9260, n_9261, n_9262, n_9263, n_9264, n_9265, n_9266;
  wire n_9267, n_9268, n_9269, n_9270, n_9271, n_9272, n_9273, n_9274;
  wire n_9275, n_9276, n_9277, n_9278, n_9279, n_9280, n_9281, n_9282;
  wire n_9283, n_9284, n_9289, n_9290, n_9291, n_9292, n_9293, n_9294;
  wire n_9295, n_9296, n_9297, n_9298, n_9299, n_9300, n_9301, n_9306;
  wire n_9307, n_9308, n_9309, n_9310, n_9311, n_9312, n_9313, n_9314;
  wire n_9315, n_9316, n_9317, n_9322, n_9323, n_9324, n_9325, n_9326;
  wire n_9327, n_9328, n_9329, n_9330, n_9331, n_9332, n_9333, n_9338;
  wire n_9339, n_9340, n_9341, n_9342, n_9343, n_9344, n_9345, n_9346;
  wire n_9347, n_9348, n_9349, n_9350, n_9351, n_9352, n_9353, n_9354;
  wire n_9355, n_9356, n_9357, n_9358, n_9359, n_9360, n_9361, n_9362;
  wire n_9363, n_9364, n_9365, n_9370, n_9371, n_9372, n_9373, n_9374;
  wire n_9375, n_9376, n_9377, n_9378, n_9379, n_9380, n_9381, n_9386;
  wire n_9387, n_9388, n_9389, n_9390, n_9391, n_9392, n_9393, n_9394;
  wire n_9395, n_9396, n_9397, n_9402, n_9403, n_9404, n_9405, n_9406;
  wire n_9407, n_9408, n_9409, n_9410, n_9411, n_9412, n_9413, n_9418;
  wire n_9419, n_9420, n_9421, n_9422, n_9423, n_9424, n_9425, n_9426;
  wire n_9427, n_9428, n_9429, n_9430, n_9431, n_9432, n_9433, n_9434;
  wire n_9435, n_9436, n_9437, n_9438, n_9439, n_9444, n_9445, n_9446;
  wire n_9447, n_9448, n_9449, n_9450, n_9451, n_9452, n_9453, n_9454;
  wire n_9455, n_9456, n_9457, n_9458, n_9459, n_9460, n_9461, n_9462;
  wire n_9463, n_9468, n_9469, n_9470, n_9471, n_9476, n_9477, n_9478;
  wire n_9479, n_9484, n_9485, n_9486, n_9487, n_9492, n_9493, n_9494;
  wire n_9495, n_9500, n_9501, n_9502, n_9503, n_9504, n_9509, n_9510;
  wire n_9511, n_9512, n_9517, n_9518, n_9519, n_9520, n_9525, n_9526;
  wire n_9527, n_9528, n_9533, n_9534, n_9535, n_9536, n_9541, n_9542;
  wire n_9543, n_9544, n_9546, n_9547, n_9548, n_9549, n_9550, n_9551;
  wire n_9552, n_9557, n_9558, n_9559, n_9560, n_9561, n_9562, n_9563;
  wire n_9564, n_9565, n_9566, n_9567, n_9568, n_9569, n_9570, n_9571;
  wire n_9572, n_9577, n_9578, n_9579, n_9580, n_9581, n_9582, n_9583;
  wire n_9584, n_9585, n_9586, n_9587, n_9588, n_9589, n_9590, n_9591;
  wire n_9592, n_9593, n_9594, n_9595, n_9596, n_9597, n_9598, n_9599;
  wire n_9600, n_9601, n_9602, n_9603, n_9604, n_9605, n_9606, n_9607;
  wire n_9608, n_9609, n_9610, n_9611, n_9612, n_9613, n_9614, n_9615;
  wire n_9616, n_9617, n_9618, n_9619, n_9620, n_9625, n_9626, n_9627;
  wire n_9628, n_9629, n_9630, n_9631, n_9632, n_9633, n_9634, n_9635;
  wire n_9636, n_9641, n_9642, n_9643, n_9644, n_9645, n_9646, n_9647;
  wire n_9648, n_9649, n_9650, n_9651, n_9652, n_9653, n_9654, n_9655;
  wire n_9656, n_9657, n_9658, n_9659, n_9660, n_9665, n_9666, n_9667;
  wire n_9668, n_9669, n_9670, n_9671, n_9672, n_9673, n_9674, n_9675;
  wire n_9676, n_9681, n_9682, n_9683, n_9684, n_9685, n_9686, n_9687;
  wire n_9688, n_9689, n_9690, n_9691, n_9692, n_9697, n_9698, n_9699;
  wire n_9700, n_9701, n_9702, n_9703, n_9704, n_9705, n_9706, n_9707;
  wire n_9708, n_9713, n_9714, n_9715, n_9716, n_9717, n_9718, n_9719;
  wire n_9720, n_9721, n_9722, n_9723, n_9724, n_9725, n_9726, n_9727;
  wire n_9728, n_9729, n_9730, n_9731, n_9732, n_9733, n_9734, n_9735;
  wire n_9736, n_9737, n_9738, n_9739, n_9740, n_9741, n_9742, n_9743;
  wire n_9744, n_9745, n_9746, n_9747, n_9748, n_9749, n_9750, n_9751;
  wire n_9752, n_9753, n_9754, n_9755, n_9756, n_9757, n_9762, n_9763;
  wire n_9764, n_9765, n_9766, n_9767, n_9768, n_9770, n_9771, n_9772;
  wire n_9773, n_9774, n_9775, n_9776, n_9777, n_9778, n_9779, n_9780;
  wire n_9781, n_9782, n_9787, n_9788, n_9789, n_9790, n_9791, n_9792;
  wire n_9793, n_9795, n_9796, n_9797, n_9798, n_9803, n_9804, n_9805;
  wire n_9806, n_9811, n_9812, n_9813, n_9814, n_9819, n_9820, n_9821;
  wire n_9822, n_9827, n_9828, n_9829, n_9830, n_9831, n_9836, n_9837;
  wire n_9838, n_9839, n_9840, n_9845, n_9846, n_9847, n_9848, n_9851;
  wire n_9852, n_9853, n_9854, n_9855, n_9856, n_9857, n_9858, n_9859;
  wire n_9860, n_9861, n_9862, n_9863, n_9864, n_9865, n_9866, n_9867;
  wire n_9868, n_9869, n_9870, n_9871, n_9872, n_9873, n_9874, n_9875;
  wire n_9876, n_9877, n_9878, n_9879, n_9880, n_9881, n_9882, n_9883;
  wire n_9884, n_9885, n_9886, n_9887, n_9888, n_9889, n_9890, n_9891;
  wire n_9892, n_9893, n_9898, n_9899, n_9900, n_9901, n_9902, n_9903;
  wire n_9904, n_9905, n_9906, n_9907, n_9908, n_9909, n_9914, n_9915;
  wire n_9916, n_9917, n_9918, n_9919, n_9920, n_9921, n_9922, n_9923;
  wire n_9924, n_9925, n_9926, n_9931, n_9932, n_9933, n_9934, n_9935;
  wire n_9936, n_9937, n_9938, n_9939, n_9940, n_9941, n_9942, n_9947;
  wire n_9948, n_9949, n_9950, n_9951, n_9952, n_9953, n_9954, n_9955;
  wire n_9956, n_9957, n_9958, n_9959, n_9964, n_9965, n_9966, n_9967;
  wire n_9968, n_9969, n_9970, n_9971, n_9972, n_9973, n_9974, n_9975;
  wire n_9980, n_9981, n_9982, n_9983, n_9984, n_9985, n_9986, n_9987;
  wire n_9988, n_9989, n_9990, n_9991, n_9996, n_9997, n_9998, n_9999;
  wire n_10000, n_10001, n_10002, n_10003, n_10004, n_10005, n_10006,
       n_10007;
  wire n_10012, n_10013, n_10014, n_10015, n_10016, n_10017, n_10018,
       n_10019;
  wire n_10020, n_10021, n_10022, n_10023, n_10024, n_10029, n_10030,
       n_10031;
  wire n_10032, n_10033, n_10034, n_10035, n_10036, n_10037, n_10038,
       n_10039;
  wire n_10040, n_10045, n_10046, n_10047, n_10048, n_10049, n_10050,
       n_10051;
  wire n_10052, n_10053, n_10054, n_10055, n_10056, n_10061, n_10062,
       n_10063;
  wire n_10064, n_10065, n_10066, n_10067, n_10068, n_10069, n_10070,
       n_10071;
  wire n_10072, n_10077, n_10078, n_10079, n_10080, n_10081, n_10082,
       n_10083;
  wire n_10084, n_10085, n_10086, n_10087, n_10088, n_10089, n_10090,
       n_10091;
  wire n_10092, n_10093, n_10094, n_10095, n_10096, n_10097, n_10098,
       n_10099;
  wire n_10100, n_10101, n_10102, n_10103, n_10104, n_10105, n_10106,
       n_10107;
  wire n_10108, n_10109, n_10110, n_10111, n_10112, n_10113, n_10114,
       n_10115;
  wire n_10116, n_10117, n_10118, n_10119, n_10120, n_10125, n_10126,
       n_10127;
  wire n_10128, n_10133, n_10134, n_10135, n_10136, n_10141, n_10142,
       n_10143;
  wire n_10144, n_10145, n_10150, n_10151, n_10152, n_10153, n_10158,
       n_10159;
  wire n_10160, n_10161, n_10166, n_10167, n_10168, n_10169, n_10174,
       n_10175;
  wire n_10176, n_10177, n_10178, n_10179, n_10180, n_10185, n_10186,
       n_10187;
  wire n_10188, n_10189, n_10190, n_10191, n_10192, n_10193, n_10194,
       n_10195;
  wire n_10196, n_10201, n_10202, n_10203, n_10204, n_10205, n_10206,
       n_10207;
  wire n_10208, n_10209, n_10210, n_10211, n_10212, n_10213, n_10214,
       n_10215;
  wire n_10216, n_10217, n_10218, n_10219, n_10220, n_10221, n_10222,
       n_10223;
  wire n_10224, n_10225, n_10226, n_10227, n_10228, n_10229, n_10230,
       n_10231;
  wire n_10232, n_10233, n_10234, n_10235, n_10236, n_10237, n_10242,
       n_10243;
  wire n_10244, n_10245, n_10246, n_10247, n_10248, n_10249, n_10250,
       n_10251;
  wire n_10252, n_10253, n_10254, n_10259, n_10260, n_10261, n_10262,
       n_10263;
  wire n_10264, n_10265, n_10266, n_10267, n_10268, n_10269, n_10270,
       n_10275;
  wire n_10276, n_10277, n_10278, n_10279, n_10280, n_10281, n_10282,
       n_10283;
  wire n_10284, n_10285, n_10286, n_10291, n_10292, n_10293, n_10294,
       n_10295;
  wire n_10296, n_10297, n_10298, n_10299, n_10300, n_10301, n_10302,
       n_10307;
  wire n_10308, n_10309, n_10310, n_10311, n_10312, n_10313, n_10314,
       n_10315;
  wire n_10316, n_10317, n_10318, n_10319, n_10320, n_10321, n_10322,
       n_10323;
  wire n_10324, n_10325, n_10326, n_10331, n_10332, n_10333, n_10334,
       n_10335;
  wire n_10336, n_10337, n_10338, n_10339, n_10340, n_10341, n_10342,
       n_10347;
  wire n_10348, n_10349, n_10350, n_10351, n_10352, n_10353, n_10354,
       n_10355;
  wire n_10356, n_10357, n_10358, n_10363, n_10364, n_10365, n_10366,
       n_10367;
  wire n_10368, n_10369, n_10370, n_10371, n_10372, n_10373, n_10374,
       n_10375;
  wire n_10380, n_10381, n_10382, n_10383, n_10384, n_10385, n_10386,
       n_10387;
  wire n_10388, n_10389, n_10390, n_10391, n_10392, n_10393, n_10394,
       n_10395;
  wire n_10396, n_10397, n_10398, n_10399, n_10400, n_10401, n_10402,
       n_10403;
  wire n_10404, n_10405, n_10406, n_10407, n_10408, n_10413, n_10414,
       n_10415;
  wire n_10416, n_10417, n_10418, n_10419, n_10420, n_10421, n_10426,
       n_10427;
  wire n_10428, n_10429, n_10430, n_10431, n_10432, n_10434, n_10435,
       n_10436;
  wire n_10437, n_10438, n_10439, n_10440, n_10441, n_10442, n_10443,
       n_10444;
  wire n_10445, n_10446, n_10447, n_10448, n_10449, n_10450, n_10451,
       n_10456;
  wire n_10457, n_10458, n_10459, n_10460, n_10461, n_10462, n_10464,
       n_10465;
  wire n_10466, n_10467, n_10472, n_10473, n_10474, n_10475, n_10480,
       n_10481;
  wire n_10482, n_10483, n_10488, n_10489, n_10490, n_10491, n_10496,
       n_10497;
  wire n_10498, n_10499, n_10500, n_10505, n_10506, n_10507, n_10508,
       n_10513;
  wire n_10514, n_10515, n_10516, n_10517, n_10522, n_10523, n_10524,
       n_10525;
  wire n_10530, n_10531, n_10532, n_10533, n_10538, n_10539, n_10540,
       n_10541;
  wire n_10546, n_10547, n_10548, n_10549, n_10554, n_10555, n_10556,
       n_10557;
  wire n_10559, n_10560, n_10561, n_10562, n_10563, n_10564, n_10565,
       n_10570;
  wire n_10571, n_10572, n_10573, n_10574, n_10575, n_10576, n_10577,
       n_10578;
  wire n_10579, n_10580, n_10581, n_10582, n_10583, n_10584, n_10585,
       n_10590;
  wire n_10591, n_10592, n_10593, n_10594, n_10595, n_10596, n_10597,
       n_10598;
  wire n_10599, n_10600, n_10601, n_10602, n_10603, n_10604, n_10605,
       n_10606;
  wire n_10607, n_10608, n_10609, n_10610, n_10611, n_10612, n_10613,
       n_10614;
  wire n_10615, n_10616, n_10617, n_10618, n_10619, n_10620, n_10621,
       n_10622;
  wire n_10623, n_10624, n_10625, n_10626, n_10627, n_10628, n_10629,
       n_10630;
  wire n_10631, n_10632, n_10633, n_10638, n_10639, n_10640, n_10641,
       n_10642;
  wire n_10643, n_10644, n_10645, n_10646, n_10647, n_10648, n_10649,
       n_10654;
  wire n_10655, n_10656, n_10657, n_10658, n_10659, n_10660, n_10661,
       n_10662;
  wire n_10663, n_10664, n_10665, n_10670, n_10671, n_10672, n_10673,
       n_10674;
  wire n_10675, n_10676, n_10677, n_10678, n_10679, n_10680, n_10681,
       n_10682;
  wire n_10683, n_10684, n_10685, n_10686, n_10687, n_10688, n_10689,
       n_10694;
  wire n_10695, n_10696, n_10697, n_10698, n_10699, n_10700, n_10701,
       n_10702;
  wire n_10703, n_10704, n_10705, n_10710, n_10711, n_10712, n_10713,
       n_10714;
  wire n_10715, n_10716, n_10717, n_10718, n_10719, n_10720, n_10721,
       n_10726;
  wire n_10727, n_10728, n_10729, n_10730, n_10731, n_10732, n_10733,
       n_10734;
  wire n_10735, n_10736, n_10737, n_10738, n_10739, n_10740, n_10741,
       n_10742;
  wire n_10743, n_10744, n_10745, n_10746, n_10747, n_10748, n_10749,
       n_10750;
  wire n_10751, n_10752, n_10753, n_10754, n_10755, n_10756, n_10757,
       n_10758;
  wire n_10759, n_10760, n_10761, n_10762, n_10763, n_10764, n_10765,
       n_10766;
  wire n_10767, n_10768, n_10769, n_10770, n_10771, n_10772, n_10773,
       n_10774;
  wire n_10775, n_10776, n_10777, n_10778, n_10779, n_10780, n_10781,
       n_10782;
  wire n_10783, n_10784, n_10785, n_10790, n_10791, n_10792, n_10793,
       n_10798;
  wire n_10799, n_10800, n_10801, n_10806, n_10807, n_10808, n_10809,
       n_10810;
  wire n_10815, n_10816, n_10817, n_10818, n_10819, n_10824, n_10825,
       n_10826;
  wire n_10827, n_10828, n_10833, n_10834, n_10835, n_10836, n_10839,
       n_10840;
  wire n_10841, n_10842, n_10843, n_10844, n_10845, n_10846, n_10847,
       n_10848;
  wire n_10849, n_10850, n_10851, n_10852, n_10853, n_10854, n_10855,
       n_10856;
  wire n_10857, n_10858, n_10859, n_10860, n_10861, n_10862, n_10863,
       n_10864;
  wire n_10865, n_10866, n_10867, n_10868, n_10869, n_10870, n_10871,
       n_10872;
  wire n_10873, n_10874, n_10875, n_10876, n_10877, n_10878, n_10879,
       n_10880;
  wire n_10881, n_10886, n_10887, n_10888, n_10889, n_10890, n_10891,
       n_10892;
  wire n_10893, n_10894, n_10895, n_10896, n_10897, n_10902, n_10903,
       n_10904;
  wire n_10905, n_10906, n_10907, n_10908, n_10909, n_10910, n_10911,
       n_10912;
  wire n_10913, n_10914, n_10919, n_10920, n_10921, n_10922, n_10923,
       n_10924;
  wire n_10925, n_10926, n_10927, n_10928, n_10929, n_10930, n_10935,
       n_10936;
  wire n_10937, n_10938, n_10939, n_10940, n_10941, n_10942, n_10943,
       n_10944;
  wire n_10945, n_10946, n_10947, n_10952, n_10953, n_10954, n_10955,
       n_10956;
  wire n_10957, n_10958, n_10959, n_10960, n_10961, n_10962, n_10963,
       n_10968;
  wire n_10969, n_10970, n_10971, n_10972, n_10973, n_10974, n_10975,
       n_10976;
  wire n_10977, n_10978, n_10979, n_10984, n_10985, n_10986, n_10987,
       n_10988;
  wire n_10989, n_10990, n_10991, n_10992, n_10993, n_10994, n_10995,
       n_11000;
  wire n_11001, n_11002, n_11003, n_11004, n_11005, n_11006, n_11007,
       n_11008;
  wire n_11009, n_11010, n_11011, n_11016, n_11017, n_11018, n_11019,
       n_11020;
  wire n_11021, n_11022, n_11023, n_11024, n_11025, n_11026, n_11027,
       n_11032;
  wire n_11033, n_11034, n_11035, n_11036, n_11037, n_11038, n_11039,
       n_11040;
  wire n_11041, n_11042, n_11043, n_11048, n_11049, n_11050, n_11051,
       n_11052;
  wire n_11053, n_11054, n_11055, n_11056, n_11057, n_11058, n_11059,
       n_11064;
  wire n_11065, n_11066, n_11067, n_11068, n_11069, n_11070, n_11071,
       n_11072;
  wire n_11073, n_11074, n_11075, n_11076, n_11077, n_11078, n_11079,
       n_11080;
  wire n_11081, n_11082, n_11083, n_11084, n_11085, n_11086, n_11087,
       n_11088;
  wire n_11089, n_11090, n_11091, n_11092, n_11093, n_11094, n_11095,
       n_11096;
  wire n_11097, n_11098, n_11099, n_11104, n_11105, n_11106, n_11107,
       n_11108;
  wire n_11109, n_11110, n_11111, n_11116, n_11117, n_11118, n_11119,
       n_11120;
  wire n_11121, n_11122, n_11124, n_11125, n_11126, n_11127, n_11128,
       n_11129;
  wire n_11130, n_11131, n_11132, n_11133, n_11134, n_11135, n_11136,
       n_11137;
  wire n_11138, n_11139, n_11144, n_11145, n_11146, n_11147, n_11148,
       n_11153;
  wire n_11154, n_11155, n_11156, n_11161, n_11162, n_11163, n_11164,
       n_11169;
  wire n_11170, n_11171, n_11172, n_11177, n_11178, n_11179, n_11180,
       n_11181;
  wire n_11182, n_11183, n_11188, n_11189, n_11190, n_11191, n_11192,
       n_11193;
  wire n_11194, n_11195, n_11196, n_11197, n_11198, n_11199, n_11204,
       n_11205;
  wire n_11206, n_11207, n_11208, n_11209, n_11210, n_11211, n_11212,
       n_11213;
  wire n_11214, n_11215, n_11216, n_11217, n_11218, n_11219, n_11220,
       n_11221;
  wire n_11222, n_11223, n_11224, n_11225, n_11226, n_11227, n_11228,
       n_11229;
  wire n_11230, n_11231, n_11232, n_11233, n_11234, n_11235, n_11236,
       n_11237;
  wire n_11238, n_11239, n_11240, n_11245, n_11246, n_11247, n_11248,
       n_11249;
  wire n_11250, n_11251, n_11252, n_11253, n_11254, n_11255, n_11256,
       n_11257;
  wire n_11262, n_11263, n_11264, n_11265, n_11266, n_11267, n_11268,
       n_11269;
  wire n_11270, n_11271, n_11272, n_11273, n_11278, n_11279, n_11280,
       n_11281;
  wire n_11282, n_11283, n_11284, n_11285, n_11286, n_11287, n_11288,
       n_11289;
  wire n_11294, n_11295, n_11296, n_11297, n_11298, n_11299, n_11300,
       n_11301;
  wire n_11302, n_11303, n_11304, n_11305, n_11310, n_11311, n_11312,
       n_11313;
  wire n_11314, n_11315, n_11316, n_11317, n_11318, n_11319, n_11320,
       n_11321;
  wire n_11326, n_11327, n_11328, n_11329, n_11330, n_11331, n_11332,
       n_11333;
  wire n_11334, n_11335, n_11336, n_11337, n_11338, n_11343, n_11344,
       n_11345;
  wire n_11346, n_11347, n_11348, n_11349, n_11350, n_11351, n_11352,
       n_11353;
  wire n_11354, n_11359, n_11360, n_11361, n_11362, n_11363, n_11364,
       n_11365;
  wire n_11366, n_11367, n_11368, n_11369, n_11370, n_11375, n_11376,
       n_11377;
  wire n_11378, n_11379, n_11380, n_11381, n_11382, n_11383, n_11384,
       n_11385;
  wire n_11386, n_11387, n_11392, n_11393, n_11394, n_11395, n_11396,
       n_11397;
  wire n_11398, n_11399, n_11400, n_11401, n_11402, n_11403, n_11404,
       n_11405;
  wire n_11406, n_11407, n_11408, n_11409, n_11410, n_11411, n_11416,
       n_11417;
  wire n_11418, n_11419, n_11420, n_11421, n_11422, n_11423, n_11424,
       n_11425;
  wire n_11426, n_11427, n_11432, n_11433, n_11434, n_11435, n_11436,
       n_11437;
  wire n_11438, n_11439, n_11444, n_11445, n_11446, n_11447, n_11448,
       n_11449;
  wire n_11450, n_11451, n_11452, n_11453, n_11454, n_11455, n_11460,
       n_11461;
  wire n_11462, n_11463, n_11464, n_11465, n_11466, n_11468, n_11469,
       n_11470;
  wire n_11471, n_11472, n_11473, n_11474, n_11475, n_11476, n_11477,
       n_11478;
  wire n_11479, n_11480, n_11481, n_11482, n_11483, n_11484, n_11489,
       n_11490;
  wire n_11491, n_11492, n_11497, n_11498, n_11499, n_11500, n_11501,
       n_11506;
  wire n_11507, n_11508, n_11509, n_11514, n_11515, n_11516, n_11517,
       n_11522;
  wire n_11523, n_11524, n_11525, n_11526, n_11531, n_11532, n_11533,
       n_11534;
  wire n_11539, n_11540, n_11541, n_11542, n_11547, n_11548, n_11549,
       n_11550;
  wire n_11552, n_11553, n_11554, n_11555, n_11556, n_11557, n_11558,
       n_11563;
  wire n_11564, n_11565, n_11566, n_11567, n_11568, n_11569, n_11570,
       n_11571;
  wire n_11576, n_11577, n_11578, n_11579, n_11580, n_11581, n_11582,
       n_11583;
  wire n_11584, n_11585, n_11586, n_11587, n_11588, n_11589, n_11590,
       n_11591;
  wire n_11592, n_11593, n_11594, n_11595, n_11600, n_11601, n_11602,
       n_11603;
  wire n_11604, n_11605, n_11606, n_11607, n_11608, n_11609, n_11610,
       n_11611;
  wire n_11612, n_11613, n_11614, n_11615, n_11616, n_11617, n_11618,
       n_11619;
  wire n_11624, n_11625, n_11626, n_11627, n_11628, n_11629, n_11630,
       n_11631;
  wire n_11632, n_11633, n_11634, n_11635, n_11636, n_11637, n_11638,
       n_11639;
  wire n_11640, n_11641, n_11642, n_11643, n_11648, n_11649, n_11650,
       n_11651;
  wire n_11652, n_11653, n_11654, n_11655, n_11656, n_11657, n_11658,
       n_11659;
  wire n_11664, n_11665, n_11666, n_11667, n_11668, n_11669, n_11670,
       n_11671;
  wire n_11672, n_11673, n_11674, n_11675, n_11680, n_11681, n_11682,
       n_11683;
  wire n_11684, n_11685, n_11686, n_11687, n_11688, n_11689, n_11690,
       n_11691;
  wire n_11692, n_11693, n_11694, n_11695, n_11696, n_11697, n_11698,
       n_11699;
  wire n_11704, n_11705, n_11706, n_11707, n_11708, n_11709, n_11710,
       n_11711;
  wire n_11712, n_11713, n_11714, n_11715, n_11720, n_11721, n_11722,
       n_11723;
  wire n_11724, n_11725, n_11726, n_11727, n_11728, n_11729, n_11730,
       n_11731;
  wire n_11732, n_11733, n_11734, n_11735, n_11736, n_11737, n_11738,
       n_11739;
  wire n_11740, n_11741, n_11742, n_11743, n_11744, n_11745, n_11746,
       n_11747;
  wire n_11748, n_11749, n_11750, n_11751, n_11752, n_11753, n_11754,
       n_11755;
  wire n_11756, n_11757, n_11758, n_11759, n_11760, n_11761, n_11762,
       n_11763;
  wire n_11768, n_11769, n_11770, n_11771, n_11772, n_11773, n_11774,
       n_11775;
  wire n_11776, n_11777, n_11778, n_11779, n_11784, n_11785, n_11786,
       n_11787;
  wire n_11788, n_11789, n_11790, n_11791, n_11796, n_11797, n_11798,
       n_11799;
  wire n_11800, n_11801, n_11802, n_11803, n_11804, n_11805, n_11806,
       n_11807;
  wire n_11812, n_11813, n_11814, n_11815, n_11816, n_11817, n_11818,
       n_11820;
  wire n_11821, n_11822, n_11823, n_11824, n_11825, n_11826, n_11827,
       n_11828;
  wire n_11829, n_11830, n_11831, n_11832, n_11833, n_11834, n_11835,
       n_11836;
  wire n_11837, n_11838, n_11839, n_11840, n_11841, n_11842, n_11843,
       n_11844;
  wire n_11845, n_11846, n_11847, n_11848, n_11849, n_11854, n_11855,
       n_11856;
  wire n_11857, n_11862, n_11863, n_11864, n_11865, n_11870, n_11871,
       n_11872;
  wire n_11873, n_11878, n_11879, n_11880, n_11881, n_11886, n_11887,
       n_11888;
  wire n_11889, n_11894, n_11895, n_11896, n_11897, n_11902, n_11903,
       n_11904;
  wire n_11905, n_11910, n_11911, n_11912, n_11913, n_11914, n_11915,
       n_11920;
  wire n_11921, n_11922, n_11923, n_11924, n_11925, n_11926, n_11927,
       n_11928;
  wire n_11929, n_11930, n_11931, n_11932, n_11937, n_11938, n_11939,
       n_11940;
  wire n_11941, n_11942, n_11943, n_11944, n_11945, n_11946, n_11947,
       n_11948;
  wire n_11949, n_11950, n_11951, n_11952, n_11953, n_11954, n_11955,
       n_11956;
  wire n_11957, n_11962, n_11963, n_11964, n_11965, n_11966, n_11967,
       n_11968;
  wire n_11969, n_11970, n_11971, n_11972, n_11973, n_11974, n_11975,
       n_11976;
  wire n_11977, n_11978, n_11979, n_11980, n_11981, n_11986, n_11987,
       n_11988;
  wire n_11989, n_11990, n_11991, n_11992, n_11993, n_11994, n_11995,
       n_11996;
  wire n_11997, n_11998, n_11999, n_12000, n_12001, n_12002, n_12003,
       n_12004;
  wire n_12005, n_12010, n_12011, n_12012, n_12013, n_12014, n_12015,
       n_12016;
  wire n_12017, n_12018, n_12019, n_12020, n_12021, n_12026, n_12027,
       n_12028;
  wire n_12029, n_12030, n_12031, n_12032, n_12033, n_12034, n_12035,
       n_12036;
  wire n_12037, n_12042, n_12043, n_12044, n_12045, n_12046, n_12047,
       n_12048;
  wire n_12049, n_12050, n_12051, n_12052, n_12053, n_12054, n_12055,
       n_12056;
  wire n_12057, n_12058, n_12059, n_12060, n_12061, n_12062, n_12067,
       n_12068;
  wire n_12069, n_12070, n_12071, n_12072, n_12073, n_12074, n_12075,
       n_12076;
  wire n_12077, n_12078, n_12083, n_12084, n_12085, n_12086, n_12087,
       n_12088;
  wire n_12089, n_12090, n_12091, n_12092, n_12093, n_12094, n_12095,
       n_12100;
  wire n_12101, n_12102, n_12103, n_12104, n_12105, n_12106, n_12107,
       n_12108;
  wire n_12109, n_12110, n_12111, n_12112, n_12113, n_12114, n_12115,
       n_12116;
  wire n_12117, n_12118, n_12119, n_12120, n_12121, n_12122, n_12123,
       n_12124;
  wire n_12125, n_12126, n_12127, n_12128, n_12129, n_12130, n_12131,
       n_12132;
  wire n_12133, n_12134, n_12135, n_12136, n_12137, n_12138, n_12139,
       n_12140;
  wire n_12141, n_12142, n_12143, n_12148, n_12149, n_12150, n_12151,
       n_12152;
  wire n_12153, n_12154, n_12155, n_12160, n_12161, n_12162, n_12163,
       n_12164;
  wire n_12165, n_12166, n_12167, n_12168, n_12169, n_12170, n_12171,
       n_12172;
  wire n_12173, n_12174, n_12175, n_12176, n_12177, n_12178, n_12179,
       n_12180;
  wire n_12181, n_12182, n_12183, n_12188, n_12189, n_12190, n_12191,
       n_12196;
  wire n_12197, n_12198, n_12199, n_12204, n_12205, n_12206, n_12207,
       n_12208;
  wire n_12209, n_12214, n_12215, n_12216, n_12217, n_12218, n_12219,
       n_12220;
  wire n_12221, n_12222, n_12223, n_12224, n_12225, n_12226, n_12231,
       n_12232;
  wire n_12233, n_12234, n_12235, n_12236, n_12237, n_12238, n_12239,
       n_12240;
  wire n_12241, n_12242, n_12247, n_12248, n_12249, n_12250, n_12251,
       n_12252;
  wire n_12253, n_12254, n_12255, n_12256, n_12257, n_12258, n_12259,
       n_12260;
  wire n_12261, n_12262, n_12263, n_12264, n_12265, n_12266, n_12271,
       n_12272;
  wire n_12273, n_12274, n_12275, n_12276, n_12277, n_12278, n_12279,
       n_12280;
  wire n_12281, n_12282, n_12287, n_12288, n_12289, n_12290, n_12291,
       n_12292;
  wire n_12293, n_12294, n_12295, n_12296, n_12297, n_12298, n_12303,
       n_12304;
  wire n_12305, n_12306, n_12307, n_12308, n_12309, n_12310, n_12311,
       n_12312;
  wire n_12313, n_12314, n_12319, n_12320, n_12321, n_12322, n_12323,
       n_12324;
  wire n_12325, n_12326, n_12327, n_12328, n_12329, n_12330, n_12335,
       n_12336;
  wire n_12337, n_12338, n_12339, n_12340, n_12341, n_12342, n_12343,
       n_12344;
  wire n_12345, n_12346, n_12351, n_12352, n_12353, n_12354, n_12355,
       n_12356;
  wire n_12357, n_12358, n_12359, n_12360, n_12361, n_12362, n_12367,
       n_12368;
  wire n_12369, n_12370, n_12371, n_12372, n_12373, n_12374, n_12375,
       n_12376;
  wire n_12377, n_12378, n_12379, n_12384, n_12385, n_12386, n_12387,
       n_12388;
  wire n_12389, n_12390, n_12391, n_12392, n_12393, n_12394, n_12395,
       n_12400;
  wire n_12401, n_12402, n_12403, n_12404, n_12405, n_12406, n_12407,
       n_12408;
  wire n_12409, n_12410, n_12411, n_12416, n_12417, n_12418, n_12419,
       n_12420;
  wire n_12421, n_12422, n_12423, n_12424, n_12425, n_12426, n_12427,
       n_12428;
  wire n_12429, n_12430, n_12431, n_12432, n_12433, n_12434, n_12435,
       n_12436;
  wire n_12437, n_12438, n_12443, n_12444, n_12445, n_12446, n_12447,
       n_12448;
  wire n_12449, n_12450, n_12451, n_12452, n_12453, n_12454, n_12455,
       n_12456;
  wire n_12457, n_12458, n_12459, n_12460, n_12461, n_12462, n_12467,
       n_12468;
  wire n_12469, n_12470, n_12471, n_12472, n_12473, n_12474, n_12479,
       n_12480;
  wire n_12481, n_12482, n_12483, n_12484, n_12485, n_12486, n_12487,
       n_12488;
  wire n_12489, n_12490, n_12495, n_12496, n_12497, n_12498, n_12499,
       n_12500;
  wire n_12501, n_12502, n_12503, n_12504, n_12505, n_12506, n_12507,
       n_12508;
  wire n_12509, n_12510, n_12511, n_12512, n_12513, n_12514, n_12515,
       n_12516;
  wire n_12517, n_12518, n_12519, n_12520, n_12521, n_12522, n_12523,
       n_12524;
  wire n_12529, n_12530, n_12531, n_12532, n_12533, n_12534, n_12535,
       n_12536;
  wire n_12537, n_12542, n_12543, n_12544, n_12545, n_12546, n_12547,
       n_12548;
  wire n_12549, n_12554, n_12555, n_12556, n_12557, n_12558, n_12559,
       n_12560;
  wire n_12561, n_12566, n_12567, n_12568, n_12569, n_12570, n_12571,
       n_12572;
  wire n_12573, n_12578, n_12579, n_12580, n_12581, n_12582, n_12583,
       n_12584;
  wire n_12585, n_12590, n_12591, n_12592, n_12593, n_12594, n_12595,
       n_12596;
  wire n_12597, n_12598, n_12599, n_12600, n_12601, n_12602, n_12603,
       n_12604;
  wire n_12605, n_12606, n_12607, n_12608, n_12609, n_12610, n_12611,
       n_12616;
  wire n_12617, n_12618, n_12619, n_12624, n_12625, n_12626, n_12627,
       n_12632;
  wire n_12633, n_12634, n_12635, n_12636, n_12637, n_12638, n_12639,
       n_12640;
  wire n_12641, n_12642, n_12643, n_12644, n_12645, n_12646, n_12647,
       n_12648;
  wire n_12649, n_12650, n_12651, n_12652, n_12653, n_12654, n_12655,
       n_12656;
  wire n_12657, n_12658, n_12663, n_12664, n_12665, n_12666, n_12667,
       n_12668;
  wire n_12669, n_12670, n_12671, n_12672, n_12673, n_12674, n_12679,
       n_12680;
  wire n_12681, n_12682, n_12683, n_12684, n_12685, n_12686, n_12687,
       n_12688;
  wire n_12689, n_12690, n_12691, n_12692, n_12693, n_12694, n_12695,
       n_12696;
  wire n_12697, n_12698, n_12699, n_12704, n_12705, n_12706, n_12707,
       n_12708;
  wire n_12709, n_12710, n_12711, n_12712, n_12713, n_12714, n_12715,
       n_12720;
  wire n_12721, n_12722, n_12723, n_12724, n_12725, n_12726, n_12727,
       n_12728;
  wire n_12729, n_12730, n_12731, n_12732, n_12733, n_12734, n_12735,
       n_12736;
  wire n_12737, n_12738, n_12739, n_12740, n_12745, n_12746, n_12747,
       n_12748;
  wire n_12749, n_12750, n_12751, n_12752, n_12753, n_12754, n_12755,
       n_12756;
  wire n_12761, n_12762, n_12763, n_12764, n_12765, n_12766, n_12767,
       n_12768;
  wire n_12769, n_12770, n_12771, n_12772, n_12773, n_12774, n_12775,
       n_12776;
  wire n_12777, n_12778, n_12779, n_12780, n_12781, n_12782, n_12783,
       n_12784;
  wire n_12785, n_12786, n_12787, n_12788, n_12789, n_12790, n_12791,
       n_12792;
  wire n_12793, n_12794, n_12795, n_12796, n_12797, n_12798, n_12799,
       n_12800;
  wire n_12801, n_12802, n_12803, n_12804, n_12805, n_12806, n_12807,
       n_12808;
  wire n_12809, n_12810, n_12811, n_12812, n_12813, n_12814, n_12815,
       n_12816;
  wire n_12817, n_12818, n_12819, n_12820, n_12821, n_12822, n_12823,
       n_12824;
  wire n_12825, n_12826, n_12827, n_12828, n_12829, n_12830, n_12831,
       n_12832;
  wire n_12833, n_12834, n_12835, n_12836, n_12837, n_12838, n_12839,
       n_12844;
  wire n_12845, n_12846, n_12847, n_12848, n_12849, n_12850, n_12851,
       n_12852;
  wire n_12853, n_12854, n_12855, n_12856, n_12857, n_12858, n_12859,
       n_12860;
  wire n_12861, n_12862, n_12863, n_12864, n_12865, n_12866, n_12867,
       n_12868;
  wire n_12869, n_12870, n_12875, n_12876, n_12877, n_12878, n_12879,
       n_12880;
  wire n_12881, n_12882, n_12887, n_12888, n_12889, n_12890, n_12891,
       n_12892;
  wire n_12893, n_12894, n_12895, n_12900, n_12901, n_12902, n_12903,
       n_12904;
  wire n_12905, n_12906, n_12907, n_12908, n_12909, n_12910, n_12911,
       n_12912;
  wire n_12913, n_12914, n_12915, n_12916, n_12917, n_12918, n_12919,
       n_12920;
  wire n_12925, n_12926, n_12927, n_12928, n_12933, n_12934, n_12935,
       n_12936;
  wire n_12941, n_12942, n_12943, n_12944, n_12945, n_12946, n_12947,
       n_12948;
  wire n_12949, n_12950, n_12951, n_12952, n_12953, n_12954, n_12955,
       n_12956;
  wire n_12957, n_12958, n_12959, n_12964, n_12965, n_12966, n_12967,
       n_12968;
  wire n_12969, n_12970, n_12971, n_12972, n_12973, n_12974, n_12975,
       n_12980;
  wire n_12981, n_12982, n_12983, n_12984, n_12985, n_12986, n_12987,
       n_12988;
  wire n_12989, n_12990, n_12991, n_12992, n_12993, n_12994, n_12995,
       n_12996;
  wire n_12997, n_12998, n_12999, n_13000, n_13005, n_13006, n_13007,
       n_13008;
  wire n_13009, n_13010, n_13011, n_13012, n_13013, n_13014, n_13015,
       n_13016;
  wire n_13021, n_13022, n_13023, n_13024, n_13025, n_13026, n_13027,
       n_13028;
  wire n_13029, n_13030, n_13031, n_13032, n_13033, n_13038, n_13039,
       n_13040;
  wire n_13041, n_13042, n_13043, n_13044, n_13045, n_13046, n_13047,
       n_13048;
  wire n_13049, n_13050, n_13055, n_13056, n_13057, n_13058, n_13059,
       n_13060;
  wire n_13061, n_13062, n_13063, n_13064, n_13065, n_13066, n_13071,
       n_13072;
  wire n_13073, n_13074, n_13075, n_13076, n_13077, n_13078, n_13079,
       n_13080;
  wire n_13081, n_13082, n_13083, n_13084, n_13085, n_13086, n_13087,
       n_13088;
  wire n_13089, n_13090, n_13091, n_13092, n_13093, n_13094, n_13095,
       n_13096;
  wire n_13097, n_13098, n_13099, n_13100, n_13101, n_13102, n_13103,
       n_13104;
  wire n_13105, n_13106, n_13107, n_13108, n_13109, n_13110, n_13111,
       n_13112;
  wire n_13113, n_13118, n_13119, n_13120, n_13121, n_13122, n_13123,
       n_13124;
  wire n_13125, n_13126, n_13127, n_13128, n_13129, n_13130, n_13131,
       n_13132;
  wire n_13133, n_13134, n_13139, n_13140, n_13141, n_13142, n_13143,
       n_13144;
  wire n_13145, n_13146, n_13147, n_13148, n_13149, n_13150, n_13151,
       n_13152;
  wire n_13153, n_13154, n_13155, n_13156, n_13157, n_13158, n_13159,
       n_13160;
  wire n_13161, n_13162, n_13163, n_13164, n_13165, n_13166, n_13167,
       n_13168;
  wire n_13169, n_13170, n_13171, n_13172, n_13173, n_13174, n_13175,
       n_13176;
  wire n_13177, n_13178, n_13179, n_13180, n_13181, n_13182, n_13183,
       n_13184;
  wire n_13185, n_13186, n_13187, n_13188, n_13189, n_13190, n_13191,
       n_13192;
  wire n_13193, n_13194, n_13195, n_13196, n_13197, n_13198, n_13199,
       n_13200;
  wire n_13201, n_13202, n_13203, n_13204, n_13205, n_13206, n_13207,
       n_13208;
  wire n_13209, n_13210, n_13211, n_13212, n_13213, n_13214, n_13215,
       n_13216;
  wire n_13217, n_13218, n_13219, n_13220, n_13221, n_13222, n_13223,
       n_13224;
  wire n_13225, n_13226, n_13227, n_13228, n_13229, n_13230, n_13235,
       n_13236;
  wire n_13237, n_13238, n_13239, n_13240, n_13241, n_13242, n_13247,
       n_13248;
  wire n_13249, n_13250, n_13251, n_13252, n_13253, n_13254, n_13255,
       n_13256;
  wire n_13257, n_13258, n_13259, n_13260, n_13261, n_13262, n_13263,
       n_13264;
  wire n_13265, n_13266, n_13267, n_13268, n_13269, n_13270, n_13275,
       n_13276;
  wire n_13277, n_13278, n_13279, n_13280, n_13281, n_13282, n_13283,
       n_13284;
  wire n_13289, n_13290, n_13291, n_13292, n_13293, n_13294, n_13295,
       n_13296;
  wire n_13301, n_13302, n_13303, n_13304, n_13305, n_13306, n_13307,
       n_13308;
  wire n_13313, n_13314, n_13315, n_13316, n_13321, n_13322, n_13323,
       n_13324;
  wire n_13329, n_13330, n_13331, n_13332, n_13337, n_13338, n_13339,
       n_13340;
  wire n_13341, n_13342, n_13343, n_13344, n_13345, n_13346, n_13347,
       n_13348;
  wire n_13349, n_13350, n_13351, n_13352, n_13353, n_13354, n_13355,
       n_13360;
  wire n_13361, n_13362, n_13363, n_13364, n_13365, n_13366, n_13367,
       n_13368;
  wire n_13369, n_13370, n_13371, n_13372, n_13373, n_13374, n_13375,
       n_13376;
  wire n_13377, n_13378, n_13379, n_13380, n_13385, n_13386, n_13387,
       n_13388;
  wire n_13389, n_13390, n_13391, n_13392, n_13393, n_13394, n_13395,
       n_13396;
  wire n_13397, n_13402, n_13403, n_13404, n_13405, n_13406, n_13407,
       n_13408;
  wire n_13409, n_13410, n_13411, n_13412, n_13413, n_13414, n_13415,
       n_13416;
  wire n_13417, n_13418, n_13419, n_13420, n_13421, n_13426, n_13427,
       n_13428;
  wire n_13429, n_13430, n_13431, n_13432, n_13433, n_13434, n_13435,
       n_13436;
  wire n_13437, n_13442, n_13443, n_13444, n_13445, n_13446, n_13447,
       n_13448;
  wire n_13449, n_13450, n_13451, n_13452, n_13453, n_13458, n_13459,
       n_13460;
  wire n_13461, n_13462, n_13463, n_13464, n_13465, n_13466, n_13467,
       n_13468;
  wire n_13469, n_13470, n_13471, n_13472, n_13473, n_13474, n_13475,
       n_13476;
  wire n_13477, n_13478, n_13479, n_13480, n_13481, n_13482, n_13483,
       n_13484;
  wire n_13485, n_13486, n_13487, n_13488, n_13489, n_13490, n_13491,
       n_13492;
  wire n_13493, n_13494, n_13495, n_13496, n_13497, n_13498, n_13499,
       n_13500;
  wire n_13501, n_13502, n_13503, n_13504, n_13505, n_13506, n_13507,
       n_13508;
  wire n_13509, n_13510, n_13511, n_13512, n_13513, n_13514, n_13515,
       n_13516;
  wire n_13517, n_13518, n_13519, n_13520, n_13521, n_13522, n_13523,
       n_13524;
  wire n_13525, n_13526, n_13527, n_13528, n_13529, n_13530, n_13531,
       n_13532;
  wire n_13533, n_13534, n_13535, n_13536, n_13537, n_13538, n_13539,
       n_13540;
  wire n_13541, n_13542, n_13543, n_13544, n_13545, n_13546, n_13547,
       n_13548;
  wire n_13549, n_13550, n_13551, n_13552, n_13553, n_13554, n_13555,
       n_13556;
  wire n_13557, n_13558, n_13559, n_13560, n_13561, n_13562, n_13563,
       n_13564;
  wire n_13569, n_13570, n_13571, n_13572, n_13573, n_13574, n_13575,
       n_13576;
  wire n_13577, n_13582, n_13583, n_13584, n_13585, n_13586, n_13587,
       n_13588;
  wire n_13589, n_13594, n_13595, n_13596, n_13597, n_13598, n_13599,
       n_13600;
  wire n_13601, n_13602, n_13607, n_13608, n_13609, n_13610, n_13611,
       n_13612;
  wire n_13613, n_13614, n_13619, n_13620, n_13621, n_13622, n_13623,
       n_13624;
  wire n_13625, n_13626, n_13627, n_13632, n_13633, n_13634, n_13635,
       n_13636;
  wire n_13637, n_13638, n_13639, n_13644, n_13645, n_13646, n_13647,
       n_13648;
  wire n_13649, n_13650, n_13651, n_13652, n_13653, n_13654, n_13655,
       n_13656;
  wire n_13657, n_13658, n_13659, n_13664, n_13665, n_13666, n_13667,
       n_13668;
  wire n_13669, n_13670, n_13671, n_13672, n_13673, n_13674, n_13675,
       n_13676;
  wire n_13677, n_13678, n_13679, n_13680, n_13685, n_13686, n_13687,
       n_13688;
  wire n_13689, n_13690, n_13691, n_13692, n_13693, n_13694, n_13695,
       n_13696;
  wire n_13697, n_13702, n_13703, n_13704, n_13705, n_13706, n_13707,
       n_13708;
  wire n_13709, n_13710, n_13711, n_13712, n_13713, n_13718, n_13719,
       n_13720;
  wire n_13721, n_13722, n_13723, n_13724, n_13725, n_13726, n_13727,
       n_13728;
  wire n_13729, n_13734, n_13735, n_13736, n_13737, n_13738, n_13739,
       n_13740;
  wire n_13741, n_13742, n_13743, n_13744, n_13745, n_13750, n_13751,
       n_13752;
  wire n_13753, n_13754, n_13755, n_13756, n_13757, n_13758, n_13759,
       n_13760;
  wire n_13761, n_13766, n_13767, n_13768, n_13769, n_13770, n_13771,
       n_13772;
  wire n_13773, n_13774, n_13775, n_13776, n_13777, n_13782, n_13783,
       n_13784;
  wire n_13785, n_13786, n_13787, n_13788, n_13789, n_13790, n_13791,
       n_13792;
  wire n_13793, n_13794, n_13799, n_13800, n_13801, n_13802, n_13803,
       n_13804;
  wire n_13805, n_13806, n_13807, n_13808, n_13809, n_13810, n_13815,
       n_13816;
  wire n_13817, n_13818, n_13819, n_13820, n_13821, n_13822, n_13823,
       n_13824;
  wire n_13825, n_13826, n_13827, n_13828, n_13829, n_13830, n_13831,
       n_13832;
  wire n_13833, n_13834, n_13835, n_13836, n_13837, n_13838, n_13843,
       n_13844;
  wire n_13845, n_13846, n_13847, n_13848, n_13849, n_13850, n_13851,
       n_13852;
  wire n_13853, n_13854, n_13855, n_13856, n_13857, n_13858, n_13859,
       n_13860;
  wire n_13865, n_13866, n_13867, n_13868, n_13869, n_13870, n_13871,
       n_13872;
  wire n_13873, n_13874, n_13875, n_13876, n_13877, n_13878, n_13879,
       n_13880;
  wire n_13881, n_13882, n_13883, n_13884, n_13885, n_13886, n_13887,
       n_13888;
  wire n_13889, n_13890, n_13891, n_13892, n_13893, n_13894, n_13895,
       n_13896;
  wire n_13897, n_13898, n_13899, n_13900, n_13901, n_13902, n_13903,
       n_13904;
  wire n_13909, n_13910, n_13911, n_13912, n_13913, n_13914, n_13915,
       n_13916;
  wire n_13917, n_13918, n_13919, n_13920, n_13921, n_13922, n_13923,
       n_13924;
  wire n_13925, n_13926, n_13927, n_13928, n_13933, n_13934, n_13935,
       n_13936;
  wire n_13937, n_13938, n_13939, n_13940, n_13945, n_13946, n_13947,
       n_13948;
  wire n_13949, n_13950, n_13951, n_13952, n_13957, n_13958, n_13959,
       n_13960;
  wire n_13961, n_13962, n_13963, n_13964, n_13965, n_13966, n_13967,
       n_13968;
  wire n_13969, n_13970, n_13971, n_13972, n_13973, n_13974, n_13975,
       n_13976;
  wire n_13977, n_13978, n_13979, n_13984, n_13985, n_13986, n_13987,
       n_13988;
  wire n_13989, n_13990, n_13991, n_13992, n_13997, n_13998, n_13999,
       n_14000;
  wire n_14001, n_14002, n_14003, n_14004, n_14009, n_14010, n_14011,
       n_14012;
  wire n_14013, n_14018, n_14019, n_14020, n_14021, n_14022, n_14023,
       n_14024;
  wire n_14025, n_14026, n_14027, n_14028, n_14029, n_14030, n_14031,
       n_14032;
  wire n_14033, n_14034, n_14035, n_14036, n_14037, n_14038, n_14039,
       n_14040;
  wire n_14041, n_14042, n_14043, n_14044, n_14045, n_14050, n_14051,
       n_14052;
  wire n_14053, n_14054, n_14055, n_14056, n_14057, n_14058, n_14059,
       n_14060;
  wire n_14061, n_14066, n_14067, n_14068, n_14069, n_14070, n_14071,
       n_14072;
  wire n_14073, n_14074, n_14075, n_14076, n_14077, n_14082, n_14083,
       n_14084;
  wire n_14085, n_14086, n_14087, n_14088, n_14089, n_14090, n_14091,
       n_14092;
  wire n_14093, n_14098, n_14099, n_14100, n_14101, n_14102, n_14103,
       n_14104;
  wire n_14105, n_14106, n_14107, n_14108, n_14109, n_14110, n_14115,
       n_14116;
  wire n_14117, n_14118, n_14119, n_14120, n_14121, n_14122, n_14123,
       n_14124;
  wire n_14125, n_14126, n_14131, n_14132, n_14133, n_14134, n_14135,
       n_14136;
  wire n_14137, n_14138, n_14139, n_14140, n_14141, n_14142, n_14147,
       n_14148;
  wire n_14149, n_14150, n_14151, n_14152, n_14153, n_14154, n_14155,
       n_14156;
  wire n_14157, n_14158, n_14159, n_14160, n_14161, n_14162, n_14163,
       n_14164;
  wire n_14165, n_14166, n_14167, n_14168, n_14169, n_14170, n_14171,
       n_14172;
  wire n_14173, n_14174, n_14175, n_14176, n_14177, n_14178, n_14179,
       n_14180;
  wire n_14181, n_14182, n_14183, n_14184, n_14185, n_14186, n_14187,
       n_14188;
  wire n_14189, n_14190, n_14191, n_14192, n_14193, n_14194, n_14195,
       n_14196;
  wire n_14197, n_14198, n_14199, n_14200, n_14201, n_14202, n_14203,
       n_14204;
  wire n_14205, n_14206, n_14207, n_14208, n_14209, n_14210, n_14211,
       n_14212;
  wire n_14213, n_14214, n_14215, n_14216, n_14217, n_14218, n_14219,
       n_14220;
  wire n_14221, n_14222, n_14223, n_14224, n_14225, n_14230, n_14231,
       n_14232;
  wire n_14233, n_14234, n_14235, n_14236, n_14237, n_14242, n_14243,
       n_14244;
  wire n_14245, n_14246, n_14247, n_14248, n_14249, n_14254, n_14255,
       n_14256;
  wire n_14257, n_14258, n_14259, n_14260, n_14261, n_14262, n_14263,
       n_14268;
  wire n_14269, n_14270, n_14271, n_14272, n_14273, n_14274, n_14275,
       n_14280;
  wire n_14281, n_14282, n_14283, n_14288, n_14289, n_14290, n_14291,
       n_14296;
  wire n_14297, n_14298, n_14299, n_14300, n_14301, n_14302, n_14303,
       n_14304;
  wire n_14305, n_14306, n_14307, n_14308, n_14313, n_14314, n_14315,
       n_14316;
  wire n_14317, n_14318, n_14319, n_14320, n_14325, n_14326, n_14327,
       n_14328;
  wire n_14329, n_14330, n_14331, n_14332, n_14333, n_14334, n_14335,
       n_14336;
  wire n_14341, n_14342, n_14343, n_14344, n_14345, n_14346, n_14347,
       n_14348;
  wire n_14349, n_14350, n_14351, n_14352, n_14357, n_14358, n_14359,
       n_14360;
  wire n_14361, n_14362, n_14363, n_14364, n_14365, n_14366, n_14367,
       n_14368;
  wire n_14369, n_14370, n_14371, n_14372, n_14373, n_14374, n_14375,
       n_14376;
  wire n_14377, n_14378, n_14379, n_14380, n_14381, n_14382, n_14383,
       n_14384;
  wire n_14389, n_14390, n_14391, n_14392, n_14393, n_14394, n_14395,
       n_14396;
  wire n_14397, n_14398, n_14399, n_14400, n_14405, n_14406, n_14407,
       n_14408;
  wire n_14409, n_14410, n_14411, n_14412, n_14413, n_14414, n_14415,
       n_14416;
  wire n_14417, n_14418, n_14419, n_14420, n_14421, n_14422, n_14423,
       n_14424;
  wire n_14429, n_14430, n_14431, n_14432, n_14433, n_14434, n_14435,
       n_14436;
  wire n_14437, n_14438, n_14439, n_14440, n_14441, n_14442, n_14443,
       n_14444;
  wire n_14445, n_14446, n_14447, n_14448, n_14449, n_14450, n_14451,
       n_14452;
  wire n_14453, n_14454, n_14455, n_14456, n_14457, n_14458, n_14459,
       n_14460;
  wire n_14461, n_14462, n_14463, n_14464, n_14465, n_14466, n_14467,
       n_14468;
  wire n_14469, n_14470, n_14471, n_14472, n_14473, n_14474, n_14475,
       n_14476;
  wire n_14477, n_14478, n_14479, n_14480, n_14481, n_14482, n_14483,
       n_14484;
  wire n_14485, n_14486, n_14487, n_14488, n_14489, n_14494, n_14495,
       n_14496;
  wire n_14497, n_14498, n_14499, n_14500, n_14501, n_14502, n_14503,
       n_14504;
  wire n_14505, n_14506, n_14507, n_14508, n_14509, n_14510, n_14511,
       n_14512;
  wire n_14513, n_14514, n_14515, n_14516, n_14517, n_14518, n_14519,
       n_14520;
  wire n_14521, n_14522, n_14523, n_14524, n_14525, n_14526, n_14527,
       n_14528;
  wire n_14529, n_14530, n_14531, n_14532, n_14533, n_14534, n_14535,
       n_14540;
  wire n_14541, n_14542, n_14543, n_14544, n_14545, n_14546, n_14547,
       n_14548;
  wire n_14549, n_14554, n_14555, n_14556, n_14557, n_14558, n_14559,
       n_14560;
  wire n_14561, n_14566, n_14567, n_14568, n_14569, n_14570, n_14571,
       n_14572;
  wire n_14573, n_14578, n_14579, n_14580, n_14581, n_14582, n_14583,
       n_14584;
  wire n_14585, n_14586, n_14591, n_14592, n_14593, n_14594, n_14595,
       n_14596;
  wire n_14597, n_14598, n_14603, n_14604, n_14605, n_14606, n_14607,
       n_14608;
  wire n_14609, n_14610, n_14611, n_14616, n_14617, n_14618, n_14619,
       n_14620;
  wire n_14621, n_14622, n_14623, n_14624, n_14629, n_14630, n_14631,
       n_14632;
  wire n_14637, n_14638, n_14639, n_14640, n_14641, n_14646, n_14647,
       n_14648;
  wire n_14649, n_14650, n_14651, n_14652, n_14653, n_14654, n_14655,
       n_14656;
  wire n_14657, n_14658, n_14659, n_14660, n_14661, n_14662, n_14663,
       n_14664;
  wire n_14665, n_14670, n_14671, n_14672, n_14673, n_14674, n_14675,
       n_14676;
  wire n_14677, n_14678, n_14679, n_14680, n_14681, n_14682, n_14683,
       n_14684;
  wire n_14685, n_14686, n_14687, n_14688, n_14689, n_14694, n_14695,
       n_14696;
  wire n_14697, n_14698, n_14699, n_14700, n_14701, n_14702, n_14703,
       n_14704;
  wire n_14705, n_14706, n_14707, n_14708, n_14709, n_14710, n_14711,
       n_14712;
  wire n_14713, n_14714, n_14719, n_14720, n_14721, n_14722, n_14723,
       n_14724;
  wire n_14725, n_14726, n_14727, n_14728, n_14729, n_14730, n_14731,
       n_14736;
  wire n_14737, n_14738, n_14739, n_14740, n_14741, n_14742, n_14743,
       n_14744;
  wire n_14745, n_14746, n_14747, n_14752, n_14753, n_14754, n_14755,
       n_14756;
  wire n_14757, n_14758, n_14759, n_14760, n_14761, n_14762, n_14763,
       n_14764;
  wire n_14769, n_14770, n_14771, n_14772, n_14773, n_14774, n_14775,
       n_14776;
  wire n_14777, n_14778, n_14779, n_14780, n_14785, n_14786, n_14787,
       n_14788;
  wire n_14789, n_14790, n_14791, n_14792, n_14793, n_14794, n_14795,
       n_14796;
  wire n_14797, n_14798, n_14799, n_14800, n_14801, n_14802, n_14803,
       n_14804;
  wire n_14805, n_14806, n_14807, n_14808, n_14809, n_14810, n_14815,
       n_14816;
  wire n_14817, n_14818, n_14819, n_14820, n_14821, n_14822, n_14823,
       n_14824;
  wire n_14825, n_14826, n_14827, n_14828, n_14829, n_14830, n_14831,
       n_14832;
  wire n_14833, n_14834, n_14835, n_14836, n_14837, n_14838, n_14839,
       n_14840;
  wire n_14841, n_14842, n_14843, n_14844, n_14845, n_14846, n_14847,
       n_14848;
  wire n_14849, n_14850, n_14851, n_14852, n_14853, n_14858, n_14859,
       n_14860;
  wire n_14861, n_14862, n_14863, n_14864, n_14865, n_14866, n_14871,
       n_14872;
  wire n_14873, n_14874, n_14875, n_14876, n_14877, n_14878, n_14883,
       n_14884;
  wire n_14885, n_14886, n_14887, n_14888, n_14889, n_14890, n_14895,
       n_14896;
  wire n_14897, n_14898, n_14899, n_14900, n_14901, n_14902, n_14903,
       n_14904;
  wire n_14909, n_14910, n_14911, n_14912, n_14913, n_14914, n_14915,
       n_14916;
  wire n_14921, n_14922, n_14923, n_14924, n_14929, n_14930, n_14931,
       n_14932;
  wire n_14933, n_14938, n_14939, n_14940, n_14941, n_14946, n_14947,
       n_14948;
  wire n_14949, n_14950, n_14951, n_14952, n_14953, n_14954, n_14955,
       n_14956;
  wire n_14957, n_14958, n_14959, n_14960, n_14961, n_14962, n_14963,
       n_14964;
  wire n_14965, n_14966, n_14967, n_14972, n_14973, n_14974, n_14975,
       n_14976;
  wire n_14977, n_14978, n_14979, n_14980, n_14981, n_14982, n_14983,
       n_14984;
  wire n_14989, n_14990, n_14991, n_14992, n_14993, n_14994, n_14995,
       n_14996;
  wire n_14997, n_14998, n_14999, n_15000, n_15005, n_15006, n_15007,
       n_15008;
  wire n_15009, n_15010, n_15011, n_15012, n_15013, n_15014, n_15015,
       n_15016;
  wire n_15021, n_15022, n_15023, n_15024, n_15025, n_15026, n_15027,
       n_15028;
  wire n_15029, n_15030, n_15031, n_15032, n_15037, n_15038, n_15039,
       n_15040;
  wire n_15041, n_15042, n_15043, n_15044, n_15045, n_15046, n_15047,
       n_15048;
  wire n_15053, n_15054, n_15055, n_15056, n_15057, n_15058, n_15059,
       n_15060;
  wire n_15061, n_15062, n_15063, n_15064, n_15065, n_15066, n_15067,
       n_15068;
  wire n_15069, n_15070, n_15071, n_15072, n_15073, n_15074, n_15075,
       n_15076;
  wire n_15077, n_15078, n_15079, n_15080, n_15081, n_15082, n_15083,
       n_15084;
  wire n_15085, n_15086, n_15087, n_15088, n_15089, n_15090, n_15091,
       n_15092;
  wire n_15093, n_15094, n_15095, n_15096, n_15097, n_15098, n_15099,
       n_15100;
  wire n_15101, n_15102, n_15103, n_15104, n_15105, n_15106, n_15107,
       n_15108;
  wire n_15109, n_15110, n_15111, n_15112, n_15113, n_15114, n_15115,
       n_15116;
  wire n_15117, n_15118, n_15119, n_15120, n_15121, n_15122, n_15123,
       n_15124;
  wire n_15125, n_15126, n_15127, n_15128, n_15129, n_15130, n_15131,
       n_15132;
  wire n_15133, n_15134, n_15135, n_15136, n_15137, n_15138, n_15139,
       n_15140;
  wire n_15141, n_15142, n_15143, n_15144, n_15145, n_15146, n_15147,
       n_15148;
  wire n_15149, n_15150, n_15151, n_15152, n_15153, n_15154, n_15155,
       n_15156;
  wire n_15157, n_15158, n_15159, n_15160, n_15161, n_15162, n_15163,
       n_15164;
  wire n_15165, n_15166, n_15167, n_15168, n_15169, n_15170, n_15171,
       n_15172;
  wire n_15173, n_15174, n_15175, n_15176, n_15177, n_15178, n_15179,
       n_15180;
  wire n_15181, n_15182, n_15183, n_15184, n_15185, n_15186, n_15187,
       n_15188;
  wire n_15189, n_15190, n_15195, n_15196, n_15197, n_15198, n_15199,
       n_15200;
  wire n_15201, n_15202, n_15207, n_15208, n_15209, n_15210, n_15211,
       n_15212;
  wire n_15213, n_15214, n_15215, n_15216, n_15217, n_15218, n_15219,
       n_15220;
  wire n_15221, n_15222, n_15223, n_15224, n_15225, n_15226, n_15227,
       n_15228;
  wire n_15233, n_15234, n_15235, n_15236, n_15237, n_15238, n_15239,
       n_15240;
  wire n_15241, n_15242, n_15243, n_15244, n_15245, n_15246, n_15247,
       n_15248;
  wire n_15249, n_15250, n_15251, n_15252, n_15257, n_15258, n_15259,
       n_15260;
  wire n_15265, n_15266, n_15267, n_15268, n_15273, n_15274, n_15275,
       n_15276;
  wire n_15281, n_15282, n_15283, n_15284, n_15285, n_15286, n_15287,
       n_15288;
  wire n_15289, n_15290, n_15291, n_15292, n_15293, n_15294, n_15295,
       n_15300;
  wire n_15301, n_15302, n_15303, n_15304, n_15305, n_15306, n_15307,
       n_15308;
  wire n_15313, n_15314, n_15315, n_15316, n_15317, n_15318, n_15319,
       n_15320;
  wire n_15321, n_15322, n_15323, n_15324, n_15325, n_15330, n_15331,
       n_15332;
  wire n_15333, n_15334, n_15335, n_15336, n_15337, n_15338, n_15339,
       n_15340;
  wire n_15341, n_15342, n_15343, n_15344, n_15345, n_15346, n_15347,
       n_15348;
  wire n_15349, n_15350, n_15351, n_15352, n_15353, n_15354, n_15355,
       n_15356;
  wire n_15357, n_15362, n_15363, n_15364, n_15365, n_15366, n_15367,
       n_15368;
  wire n_15369, n_15370, n_15371, n_15372, n_15373, n_15378, n_15379,
       n_15380;
  wire n_15381, n_15382, n_15383, n_15384, n_15385, n_15386, n_15387,
       n_15388;
  wire n_15389, n_15390, n_15391, n_15392, n_15393, n_15394, n_15395,
       n_15396;
  wire n_15397, n_15402, n_15403, n_15404, n_15405, n_15406, n_15407,
       n_15408;
  wire n_15409, n_15410, n_15411, n_15412, n_15413, n_15414, n_15415,
       n_15416;
  wire n_15417, n_15418, n_15419, n_15420, n_15421, n_15422, n_15423,
       n_15424;
  wire n_15425, n_15426, n_15427, n_15428, n_15429, n_15430, n_15431,
       n_15432;
  wire n_15433, n_15434, n_15435, n_15436, n_15437, n_15438, n_15439,
       n_15440;
  wire n_15441, n_15442, n_15443, n_15444, n_15445, n_15446, n_15447,
       n_15448;
  wire n_15449, n_15450, n_15451, n_15452, n_15453, n_15454, n_15455,
       n_15456;
  wire n_15457, n_15458, n_15459, n_15460, n_15461, n_15462, n_15463,
       n_15464;
  wire n_15465, n_15466, n_15467, n_15468, n_15469, n_15470, n_15471,
       n_15472;
  wire n_15473, n_15478, n_15479, n_15480, n_15481, n_15482, n_15483,
       n_15484;
  wire n_15485, n_15486, n_15491, n_15492, n_15493, n_15494, n_15495,
       n_15496;
  wire n_15497, n_15498, n_15503, n_15504, n_15505, n_15506, n_15507,
       n_15508;
  wire n_15509, n_15510, n_15515, n_15516, n_15517, n_15518, n_15519,
       n_15520;
  wire n_15521, n_15522, n_15523, n_15528, n_15529, n_15530, n_15531,
       n_15532;
  wire n_15533, n_15534, n_15535, n_15540, n_15541, n_15542, n_15543,
       n_15544;
  wire n_15545, n_15546, n_15547, n_15552, n_15553, n_15554, n_15555,
       n_15560;
  wire n_15561, n_15562, n_15563, n_15564, n_15565, n_15566, n_15567,
       n_15568;
  wire n_15569, n_15570, n_15571, n_15572, n_15573, n_15574, n_15575,
       n_15576;
  wire n_15577, n_15578, n_15579, n_15580, n_15581, n_15586, n_15587,
       n_15588;
  wire n_15589, n_15590, n_15591, n_15592, n_15593, n_15594, n_15595,
       n_15596;
  wire n_15597, n_15598, n_15603, n_15604, n_15605, n_15606, n_15607,
       n_15608;
  wire n_15609, n_15610, n_15611, n_15612, n_15613, n_15614, n_15615,
       n_15616;
  wire n_15617, n_15618, n_15619, n_15620, n_15621, n_15622, n_15623,
       n_15628;
  wire n_15629, n_15630, n_15631, n_15632, n_15633, n_15634, n_15635,
       n_15636;
  wire n_15637, n_15638, n_15639, n_15640, n_15645, n_15646, n_15647,
       n_15648;
  wire n_15649, n_15650, n_15651, n_15652, n_15653, n_15654, n_15655,
       n_15656;
  wire n_15661, n_15662, n_15663, n_15664, n_15665, n_15666, n_15667,
       n_15668;
  wire n_15669, n_15670, n_15671, n_15672, n_15673, n_15678, n_15679,
       n_15680;
  wire n_15681, n_15682, n_15683, n_15684, n_15685, n_15686, n_15687,
       n_15688;
  wire n_15689, n_15694, n_15695, n_15696, n_15697, n_15698, n_15699,
       n_15700;
  wire n_15701, n_15702, n_15703, n_15704, n_15705, n_15710, n_15711,
       n_15712;
  wire n_15713, n_15714, n_15715, n_15716, n_15717, n_15718, n_15719,
       n_15720;
  wire n_15721, n_15726, n_15727, n_15728, n_15729, n_15730, n_15731,
       n_15732;
  wire n_15733, n_15734, n_15735, n_15736, n_15737, n_15738, n_15739,
       n_15740;
  wire n_15741, n_15742, n_15743, n_15744, n_15745, n_15746, n_15747,
       n_15748;
  wire n_15749, n_15750, n_15751, n_15752, n_15753, n_15754, n_15755,
       n_15756;
  wire n_15757, n_15758, n_15759, n_15760, n_15761, n_15762, n_15763,
       n_15764;
  wire n_15765, n_15766, n_15767, n_15768, n_15769, n_15770, n_15771,
       n_15772;
  wire n_15777, n_15778, n_15779, n_15780, n_15781, n_15782, n_15783,
       n_15784;
  wire n_15785, n_15790, n_15791, n_15792, n_15793, n_15794, n_15795,
       n_15796;
  wire n_15797, n_15798, n_15803, n_15804, n_15805, n_15806, n_15807,
       n_15808;
  wire n_15809, n_15810, n_15811, n_15816, n_15817, n_15818, n_15819,
       n_15820;
  wire n_15825, n_15826, n_15827, n_15828, n_15833, n_15834, n_15835,
       n_15836;
  wire n_15837, n_15842, n_15843, n_15844, n_15845, n_15850, n_15851,
       n_15852;
  wire n_15853, n_15854, n_15855, n_15856, n_15857, n_15858, n_15859,
       n_15860;
  wire n_15865, n_15866, n_15867, n_15868, n_15869, n_15870, n_15871,
       n_15872;
  wire n_15873, n_15874, n_15875, n_15876, n_15881, n_15882, n_15883,
       n_15884;
  wire n_15885, n_15886, n_15887, n_15888, n_15889, n_15890, n_15891,
       n_15892;
  wire n_15897, n_15898, n_15899, n_15900, n_15901, n_15902, n_15903,
       n_15904;
  wire n_15905, n_15906, n_15907, n_15908, n_15913, n_15914, n_15915,
       n_15916;
  wire n_15917, n_15918, n_15919, n_15920, n_15921, n_15922, n_15923,
       n_15924;
  wire n_15929, n_15930, n_15931, n_15932, n_15933, n_15934, n_15935,
       n_15936;
  wire n_15937, n_15938, n_15939, n_15940, n_15941, n_15942, n_15943,
       n_15944;
  wire n_15945, n_15946, n_15947, n_15948, n_15949, n_15950, n_15951,
       n_15952;
  wire n_15953, n_15954, n_15955, n_15956, n_15957, n_15958, n_15959,
       n_15960;
  wire n_15961, n_15962, n_15963, n_15964, n_15965, n_15966, n_15967,
       n_15968;
  wire n_15969, n_15970, n_15971, n_15972, n_15973, n_15974, n_15975,
       n_15976;
  wire n_15977, n_15978, n_15979, n_15980, n_15981, n_15982, n_15983,
       n_15984;
  wire n_15985, n_15986, n_15987, n_15988, n_15989, n_15990, n_15991,
       n_15992;
  wire n_15993, n_15994, n_15995, n_15996, n_15997, n_15998, n_15999,
       n_16000;
  wire n_16001, n_16002, n_16003, n_16004, n_16005, n_16006, n_16007,
       n_16008;
  wire n_16009, n_16010, n_16011, n_16012, n_16013, n_16014, n_16015,
       n_16016;
  wire n_16017, n_16018, n_16019, n_16020, n_16021, n_16022, n_16023,
       n_16024;
  wire n_16025, n_16026, n_16027, n_16028, n_16029, n_16030, n_16031,
       n_16032;
  wire n_16033, n_16034, n_16035, n_16036, n_16037, n_16038, n_16039,
       n_16040;
  wire n_16041, n_16042, n_16043, n_16044, n_16045, n_16046, n_16047,
       n_16048;
  wire n_16049, n_16050, n_16051, n_16052, n_16053, n_16054, n_16055,
       n_16056;
  wire n_16057, n_16058, n_16059, n_16060, n_16061, n_16062, n_16063,
       n_16064;
  wire n_16065, n_16066, n_16067, n_16068, n_16069, n_16070, n_16071,
       n_16072;
  wire n_16073, n_16074, n_16075, n_16076, n_16077, n_16078, n_16079,
       n_16080;
  wire n_16081, n_16086, n_16087, n_16088, n_16089, n_16090, n_16091,
       n_16092;
  wire n_16093, n_16098, n_16099, n_16100, n_16101, n_16102, n_16103,
       n_16104;
  wire n_16105, n_16110, n_16111, n_16112, n_16113, n_16114, n_16115,
       n_16116;
  wire n_16117, n_16118, n_16119, n_16120, n_16121, n_16122, n_16123,
       n_16124;
  wire n_16125, n_16126, n_16127, n_16128, n_16129, n_16130, n_16135,
       n_16136;
  wire n_16137, n_16138, n_16143, n_16144, n_16145, n_16146, n_16151,
       n_16152;
  wire n_16153, n_16154, n_16155, n_16156, n_16157, n_16158, n_16159,
       n_16160;
  wire n_16161, n_16162, n_16163, n_16164, n_16165, n_16166, n_16167,
       n_16168;
  wire n_16169, n_16170, n_16171, n_16172, n_16173, n_16174, n_16175,
       n_16176;
  wire n_16177, n_16178, n_16183, n_16184, n_16185, n_16186, n_16187,
       n_16188;
  wire n_16189, n_16190, n_16191, n_16192, n_16193, n_16194, n_16199,
       n_16200;
  wire n_16201, n_16202, n_16203, n_16204, n_16205, n_16206, n_16207,
       n_16208;
  wire n_16209, n_16210, n_16211, n_16212, n_16213, n_16214, n_16215,
       n_16216;
  wire n_16217, n_16218, n_16223, n_16224, n_16225, n_16226, n_16227,
       n_16228;
  wire n_16229, n_16230, n_16231, n_16232, n_16233, n_16234, n_16235,
       n_16240;
  wire n_16241, n_16242, n_16243, n_16244, n_16245, n_16246, n_16247,
       n_16248;
  wire n_16249, n_16250, n_16251, n_16256, n_16257, n_16258, n_16259,
       n_16260;
  wire n_16261, n_16262, n_16263, n_16264, n_16265, n_16266, n_16267,
       n_16272;
  wire n_16273, n_16274, n_16275, n_16276, n_16277, n_16278, n_16279,
       n_16280;
  wire n_16281, n_16282, n_16283, n_16284, n_16285, n_16286, n_16287,
       n_16288;
  wire n_16289, n_16290, n_16291, n_16292, n_16293, n_16294, n_16295,
       n_16296;
  wire n_16297, n_16298, n_16299, n_16300, n_16301, n_16302, n_16303,
       n_16304;
  wire n_16305, n_16306, n_16307, n_16308, n_16309, n_16310, n_16311,
       n_16312;
  wire n_16313, n_16314, n_16315, n_16316, n_16317, n_16318, n_16319,
       n_16320;
  wire n_16321, n_16322, n_16323, n_16324, n_16325, n_16326, n_16327,
       n_16328;
  wire n_16329, n_16330, n_16331, n_16332, n_16333, n_16334, n_16335,
       n_16336;
  wire n_16337, n_16338, n_16339, n_16340, n_16341, n_16342, n_16343,
       n_16344;
  wire n_16345, n_16346, n_16347, n_16348, n_16349, n_16350, n_16351,
       n_16352;
  wire n_16353, n_16354, n_16355, n_16360, n_16361, n_16362, n_16363,
       n_16364;
  wire n_16365, n_16366, n_16367, n_16368, n_16373, n_16374, n_16375,
       n_16376;
  wire n_16377, n_16378, n_16379, n_16380, n_16385, n_16386, n_16387,
       n_16388;
  wire n_16389, n_16390, n_16391, n_16392, n_16397, n_16398, n_16399,
       n_16400;
  wire n_16401, n_16402, n_16403, n_16404, n_16409, n_16410, n_16411,
       n_16412;
  wire n_16413, n_16414, n_16415, n_16416, n_16417, n_16418, n_16419,
       n_16420;
  wire n_16421, n_16422, n_16423, n_16424, n_16425, n_16426, n_16427,
       n_16432;
  wire n_16433, n_16434, n_16435, n_16436, n_16437, n_16438, n_16439,
       n_16440;
  wire n_16441, n_16442, n_16443, n_16444, n_16449, n_16450, n_16451,
       n_16452;
  wire n_16453, n_16454, n_16455, n_16456, n_16457, n_16458, n_16459,
       n_16460;
  wire n_16465, n_16466, n_16467, n_16468, n_16469, n_16470, n_16471,
       n_16472;
  wire n_16473, n_16474, n_16475, n_16476, n_16481, n_16482, n_16483,
       n_16484;
  wire n_16485, n_16486, n_16487, n_16488, n_16489, n_16490, n_16491,
       n_16492;
  wire n_16493, n_16498, n_16499, n_16500, n_16501, n_16502, n_16503,
       n_16504;
  wire n_16505, n_16506, n_16507, n_16508, n_16509, n_16514, n_16515,
       n_16516;
  wire n_16517, n_16518, n_16519, n_16520, n_16521, n_16522, n_16523,
       n_16524;
  wire n_16525, n_16530, n_16531, n_16532, n_16533, n_16534, n_16535,
       n_16536;
  wire n_16537, n_16538, n_16539, n_16540, n_16541, n_16546, n_16547,
       n_16548;
  wire n_16549, n_16550, n_16551, n_16552, n_16553, n_16554, n_16555,
       n_16556;
  wire n_16557, n_16562, n_16563, n_16564, n_16565, n_16566, n_16567,
       n_16568;
  wire n_16569, n_16570, n_16571, n_16572, n_16573, n_16578, n_16579,
       n_16580;
  wire n_16581, n_16582, n_16583, n_16584, n_16585, n_16586, n_16587,
       n_16588;
  wire n_16589, n_16594, n_16595, n_16596, n_16597, n_16598, n_16599,
       n_16600;
  wire n_16601, n_16602, n_16603, n_16604, n_16605, n_16606, n_16607,
       n_16608;
  wire n_16609, n_16610, n_16611, n_16612, n_16613, n_16614, n_16615,
       n_16616;
  wire n_16617, n_16618, n_16619, n_16620, n_16621, n_16622, n_16623,
       n_16624;
  wire n_16625, n_16626, n_16627, n_16628, n_16629, n_16630, n_16631,
       n_16632;
  wire n_16633, n_16634, n_16635, n_16636, n_16637, n_16638, n_16639,
       n_16640;
  wire n_16641, n_16642, n_16643, n_16644, n_16649, n_16650, n_16651,
       n_16652;
  wire n_16653, n_16654, n_16655, n_16656, n_16657, n_16658, n_16659,
       n_16660;
  wire n_16661, n_16662, n_16663, n_16664, n_16665, n_16666, n_16667,
       n_16668;
  wire n_16669, n_16674, n_16675, n_16676, n_16677, n_16678, n_16679,
       n_16680;
  wire n_16681, n_16686, n_16687, n_16688, n_16689, n_16690, n_16691,
       n_16692;
  wire n_16693, n_16694, n_16699, n_16700, n_16701, n_16702, n_16703,
       n_16704;
  wire n_16705, n_16706, n_16711, n_16712, n_16713, n_16714, n_16715,
       n_16720;
  wire n_16721, n_16722, n_16723, n_16728, n_16729, n_16730, n_16731,
       n_16732;
  wire n_16737, n_16738, n_16739, n_16740, n_16741, n_16742, n_16743,
       n_16744;
  wire n_16745, n_16746, n_16747, n_16748, n_16749, n_16750, n_16751,
       n_16752;
  wire n_16753, n_16754, n_16755, n_16756, n_16757, n_16758, n_16759,
       n_16760;
  wire n_16761, n_16762, n_16763, n_16768, n_16769, n_16770, n_16771,
       n_16772;
  wire n_16773, n_16774, n_16775, n_16776, n_16777, n_16778, n_16779,
       n_16784;
  wire n_16785, n_16786, n_16787, n_16788, n_16789, n_16790, n_16791,
       n_16792;
  wire n_16793, n_16794, n_16795, n_16800, n_16801, n_16802, n_16803,
       n_16804;
  wire n_16805, n_16806, n_16807, n_16808, n_16809, n_16810, n_16811,
       n_16812;
  wire n_16813, n_16814, n_16815, n_16816, n_16817, n_16818, n_16819,
       n_16824;
  wire n_16825, n_16826, n_16827, n_16828, n_16829, n_16830, n_16831,
       n_16832;
  wire n_16833, n_16834, n_16835, n_16836, n_16837, n_16838, n_16839,
       n_16840;
  wire n_16841, n_16842, n_16843, n_16844, n_16845, n_16846, n_16847,
       n_16848;
  wire n_16849, n_16850, n_16851, n_16852, n_16853, n_16854, n_16855,
       n_16856;
  wire n_16857, n_16858, n_16859, n_16864, n_16865, n_16866, n_16867,
       n_16868;
  wire n_16869, n_16870, n_16871, n_16872, n_16873, n_16874, n_16875,
       n_16876;
  wire n_16877, n_16878, n_16879, n_16880, n_16881, n_16882, n_16883,
       n_16884;
  wire n_16885, n_16886, n_16887, n_16888, n_16889, n_16890, n_16891,
       n_16892;
  wire n_16893, n_16894, n_16895, n_16896, n_16897, n_16898, n_16899,
       n_16900;
  wire n_16901, n_16902, n_16903, n_16904, n_16905, n_16906, n_16907,
       n_16908;
  wire n_16909, n_16910, n_16911, n_16912, n_16917, n_16918, n_16919,
       n_16920;
  wire n_16921, n_16922, n_16923, n_16924, n_16929, n_16930, n_16931,
       n_16932;
  wire n_16933, n_16934, n_16935, n_16936, n_16937, n_16942, n_16943,
       n_16944;
  wire n_16945, n_16946, n_16947, n_16948, n_16949, n_16954, n_16955,
       n_16956;
  wire n_16957, n_16958, n_16959, n_16960, n_16961, n_16962, n_16967,
       n_16968;
  wire n_16969, n_16970, n_16971, n_16972, n_16973, n_16974, n_16979,
       n_16980;
  wire n_16981, n_16982, n_16987, n_16988, n_16989, n_16990, n_16995,
       n_16996;
  wire n_16997, n_16998, n_17003, n_17004, n_17005, n_17006, n_17007,
       n_17008;
  wire n_17009, n_17010, n_17011, n_17012, n_17013, n_17014, n_17015,
       n_17016;
  wire n_17017, n_17018, n_17019, n_17024, n_17025, n_17026, n_17027,
       n_17028;
  wire n_17029, n_17030, n_17031, n_17032, n_17033, n_17034, n_17035,
       n_17036;
  wire n_17037, n_17038, n_17039, n_17040, n_17041, n_17042, n_17043,
       n_17048;
  wire n_17049, n_17050, n_17051, n_17052, n_17053, n_17054, n_17055,
       n_17056;
  wire n_17057, n_17058, n_17059, n_17060, n_17061, n_17066, n_17067,
       n_17068;
  wire n_17069, n_17070, n_17071, n_17072, n_17073, n_17074, n_17075,
       n_17076;
  wire n_17077, n_17082, n_17083, n_17084, n_17085, n_17086, n_17087,
       n_17088;
  wire n_17089, n_17090, n_17091, n_17092, n_17093, n_17094, n_17099,
       n_17100;
  wire n_17101, n_17102, n_17103, n_17104, n_17105, n_17106, n_17107,
       n_17108;
  wire n_17109, n_17110, n_17111, n_17112, n_17113, n_17114, n_17115,
       n_17116;
  wire n_17117, n_17118, n_17119, n_17120, n_17121, n_17122, n_17123,
       n_17124;
  wire n_17125, n_17126, n_17131, n_17132, n_17133, n_17134, n_17135,
       n_17136;
  wire n_17137, n_17138, n_17139, n_17140, n_17141, n_17142, n_17143,
       n_17144;
  wire n_17145, n_17146, n_17147, n_17148, n_17149, n_17150, n_17151,
       n_17152;
  wire n_17153, n_17154, n_17155, n_17156, n_17157, n_17158, n_17159,
       n_17160;
  wire n_17161, n_17162, n_17163, n_17164, n_17165, n_17166, n_17167,
       n_17168;
  wire n_17169, n_17170, n_17175, n_17176, n_17177, n_17178, n_17179,
       n_17180;
  wire n_17181, n_17182, n_17183, n_17188, n_17189, n_17190, n_17191,
       n_17192;
  wire n_17193, n_17194, n_17195, n_17200, n_17201, n_17202, n_17203,
       n_17204;
  wire n_17205, n_17206, n_17207, n_17208, n_17213, n_17214, n_17215,
       n_17216;
  wire n_17221, n_17222, n_17223, n_17224, n_17225, n_17226, n_17227,
       n_17228;
  wire n_17229, n_17230, n_17231, n_17232, n_17233, n_17234, n_17235,
       n_17236;
  wire n_17237, n_17238, n_17239, n_17240, n_17241, n_17246, n_17247,
       n_17248;
  wire n_17249, n_17250, n_17251, n_17252, n_17253, n_17254, n_17255,
       n_17256;
  wire n_17257, n_17258, n_17259, n_17260, n_17261, n_17262, n_17263,
       n_17264;
  wire n_17265, n_17270, n_17271, n_17272, n_17273, n_17274, n_17275,
       n_17276;
  wire n_17277, n_17278, n_17279, n_17280, n_17281, n_17286, n_17287,
       n_17288;
  wire n_17289, n_17290, n_17291, n_17292, n_17293, n_17294, n_17295,
       n_17296;
  wire n_17297, n_17298, n_17303, n_17304, n_17305, n_17306, n_17307,
       n_17308;
  wire n_17309, n_17310, n_17311, n_17312, n_17313, n_17314, n_17319,
       n_17320;
  wire n_17321, n_17322, n_17323, n_17324, n_17325, n_17326, n_17327,
       n_17328;
  wire n_17329, n_17330, n_17335, n_17336, n_17337, n_17338, n_17339,
       n_17340;
  wire n_17341, n_17342, n_17343, n_17344, n_17345, n_17346, n_17351,
       n_17352;
  wire n_17353, n_17354, n_17355, n_17356, n_17357, n_17358, n_17359,
       n_17360;
  wire n_17361, n_17362, n_17367, n_17368, n_17369, n_17370, n_17371,
       n_17372;
  wire n_17373, n_17374, n_17375, n_17376, n_17377, n_17378, n_17383,
       n_17384;
  wire n_17385, n_17386, n_17387, n_17388, n_17389, n_17390, n_17391,
       n_17392;
  wire n_17393, n_17394, n_17395, n_17396, n_17397, n_17402, n_17403,
       n_17404;
  wire n_17405, n_17406, n_17407, n_17408, n_17409, n_17410, n_17411,
       n_17412;
  wire n_17413, n_17414, n_17415, n_17416, n_17417, n_17418, n_17419,
       n_17420;
  wire n_17421, n_17422, n_17423, n_17424, n_17425, n_17426, n_17427,
       n_17428;
  wire n_17429, n_17430, n_17431, n_17436, n_17437, n_17438, n_17439,
       n_17440;
  wire n_17441, n_17442, n_17443, n_17448, n_17449, n_17450, n_17451,
       n_17452;
  wire n_17453, n_17454, n_17455, n_17460, n_17461, n_17462, n_17463,
       n_17464;
  wire n_17465, n_17466, n_17467, n_17472, n_17473, n_17474, n_17475,
       n_17476;
  wire n_17477, n_17478, n_17479, n_17484, n_17485, n_17486, n_17487,
       n_17488;
  wire n_17493, n_17494, n_17495, n_17496, n_17501, n_17502, n_17503,
       n_17504;
  wire n_17509, n_17510, n_17511, n_17512, n_17513, n_17514, n_17515,
       n_17516;
  wire n_17517, n_17518, n_17523, n_17524, n_17525, n_17526, n_17527,
       n_17528;
  wire n_17529, n_17530, n_17531, n_17532, n_17533, n_17534, n_17535,
       n_17536;
  wire n_17537, n_17538, n_17539, n_17540, n_17541, n_17542, n_17547,
       n_17548;
  wire n_17549, n_17550, n_17551, n_17552, n_17553, n_17554, n_17555,
       n_17556;
  wire n_17557, n_17558, n_17559, n_17560, n_17561, n_17562, n_17563,
       n_17564;
  wire n_17565, n_17566, n_17571, n_17572, n_17573, n_17574, n_17575,
       n_17576;
  wire n_17577, n_17578, n_17579, n_17580, n_17581, n_17582, n_17583,
       n_17588;
  wire n_17589, n_17590, n_17591, n_17592, n_17593, n_17594, n_17595,
       n_17596;
  wire n_17597, n_17598, n_17599, n_17600, n_17601, n_17602, n_17603,
       n_17604;
  wire n_17605, n_17606, n_17607, n_17608, n_17609, n_17610, n_17611,
       n_17612;
  wire n_17613, n_17614, n_17615, n_17620, n_17621, n_17622, n_17623,
       n_17624;
  wire n_17625, n_17626, n_17627, n_17628, n_17629, n_17630, n_17631,
       n_17636;
  wire n_17637, n_17638, n_17639, n_17640, n_17641, n_17642, n_17643,
       n_17644;
  wire n_17645, n_17646, n_17647, n_17648, n_17649, n_17650, n_17651,
       n_17652;
  wire n_17653, n_17654, n_17655, n_17656, n_17657, n_17658, n_17659,
       n_17660;
  wire n_17661, n_17662, n_17663, n_17664, n_17665, n_17666, n_17667,
       n_17668;
  wire n_17669, n_17670, n_17671, n_17672, n_17673, n_17674, n_17675,
       n_17676;
  wire n_17677, n_17678, n_17679, n_17680, n_17681, n_17682, n_17683,
       n_17684;
  wire n_17685, n_17686, n_17687, n_17688, n_17689, n_17690, n_17691,
       n_17692;
  wire n_17697, n_17698, n_17699, n_17700, n_17701, n_17702, n_17703,
       n_17704;
  wire n_17705, n_17710, n_17711, n_17712, n_17713, n_17714, n_17715,
       n_17716;
  wire n_17717, n_17722, n_17723, n_17724, n_17725, n_17726, n_17727,
       n_17728;
  wire n_17729, n_17730, n_17735, n_17736, n_17737, n_17738, n_17739,
       n_17740;
  wire n_17741, n_17742, n_17747, n_17748, n_17749, n_17750, n_17755,
       n_17756;
  wire n_17757, n_17758, n_17763, n_17764, n_17765, n_17766, n_17771,
       n_17772;
  wire n_17773, n_17774, n_17779, n_17780, n_17781, n_17782, n_17783,
       n_17784;
  wire n_17785, n_17786, n_17787, n_17788, n_17789, n_17790, n_17791,
       n_17792;
  wire n_17793, n_17794, n_17795, n_17796, n_17797, n_17798, n_17799,
       n_17800;
  wire n_17801, n_17802, n_17803, n_17804, n_17805, n_17806, n_17807,
       n_17808;
  wire n_17809, n_17810, n_17811, n_17812, n_17817, n_17818, n_17819,
       n_17820;
  wire n_17821, n_17822, n_17823, n_17824, n_17825, n_17826, n_17827,
       n_17828;
  wire n_17829, n_17830, n_17835, n_17836, n_17837, n_17838, n_17839,
       n_17840;
  wire n_17841, n_17842, n_17843, n_17844, n_17845, n_17846, n_17847,
       n_17848;
  wire n_17849, n_17850, n_17851, n_17852, n_17853, n_17854, n_17855,
       n_17856;
  wire n_17857, n_17858, n_17859, n_17860, n_17861, n_17862, n_17863,
       n_17864;
  wire n_17865, n_17866, n_17867, n_17868, n_17869, n_17870, n_17871,
       n_17872;
  wire n_17873, n_17874, n_17875, n_17876, n_17877, n_17878, n_17883,
       n_17884;
  wire n_17885, n_17886, n_17887, n_17888, n_17889, n_17890, n_17891,
       n_17892;
  wire n_17893, n_17894, n_17899, n_17900, n_17901, n_17902, n_17903,
       n_17904;
  wire n_17905, n_17906, n_17907, n_17908, n_17909, n_17910, n_17911,
       n_17912;
  wire n_17913, n_17914, n_17915, n_17916, n_17917, n_17918, n_17919,
       n_17920;
  wire n_17921, n_17922, n_17923, n_17924, n_17925, n_17926, n_17927,
       n_17928;
  wire n_17929, n_17930, n_17931, n_17932, n_17933, n_17934, n_17939,
       n_17940;
  wire n_17941, n_17942, n_17943, n_17944, n_17945, n_17946, n_17947,
       n_17952;
  wire n_17953, n_17954, n_17955, n_17956, n_17957, n_17958, n_17959,
       n_17960;
  wire n_17965, n_17966, n_17967, n_17968, n_17969, n_17970, n_17971,
       n_17972;
  wire n_17977, n_17978, n_17979, n_17980, n_17981, n_17982, n_17983,
       n_17984;
  wire n_17985, n_17986, n_17987, n_17988, n_17989, n_17990, n_17991,
       n_17992;
  wire n_17997, n_17998, n_17999, n_18000, n_18001, n_18002, n_18003,
       n_18004;
  wire n_18005, n_18006, n_18007, n_18008, n_18009, n_18014, n_18015,
       n_18016;
  wire n_18017, n_18018, n_18019, n_18020, n_18021, n_18022, n_18023,
       n_18024;
  wire n_18025, n_18026, n_18031, n_18032, n_18033, n_18034, n_18035,
       n_18036;
  wire n_18037, n_18038, n_18039, n_18040, n_18041, n_18042, n_18047,
       n_18048;
  wire n_18049, n_18050, n_18051, n_18052, n_18053, n_18054, n_18055,
       n_18056;
  wire n_18057, n_18058, n_18059, n_18064, n_18065, n_18066, n_18067,
       n_18068;
  wire n_18069, n_18070, n_18071, n_18072, n_18073, n_18074, n_18075,
       n_18080;
  wire n_18081, n_18082, n_18083, n_18084, n_18085, n_18086, n_18087,
       n_18088;
  wire n_18089, n_18090, n_18091, n_18096, n_18097, n_18098, n_18099,
       n_18100;
  wire n_18101, n_18102, n_18103, n_18104, n_18105, n_18106, n_18107,
       n_18112;
  wire n_18113, n_18114, n_18115, n_18116, n_18117, n_18118, n_18119,
       n_18120;
  wire n_18121, n_18122, n_18123, n_18128, n_18129, n_18130, n_18131,
       n_18132;
  wire n_18133, n_18134, n_18135, n_18136, n_18137, n_18138, n_18139,
       n_18144;
  wire n_18145, n_18146, n_18147, n_18148, n_18149, n_18150, n_18151,
       n_18152;
  wire n_18153, n_18154, n_18155, n_18156, n_18157, n_18158, n_18159,
       n_18160;
  wire n_18161, n_18162, n_18163, n_18164, n_18165, n_18166, n_18167,
       n_18168;
  wire n_18169, n_18170, n_18171, n_18172, n_18173, n_18174, n_18175,
       n_18176;
  wire n_18177, n_18178, n_18179, n_18180, n_18181, n_18182, n_18183,
       n_18184;
  wire n_18185, n_18186, n_18187, n_18188, n_18189, n_18190, n_18195,
       n_18196;
  wire n_18197, n_18198, n_18199, n_18200, n_18201, n_18202, n_18203,
       n_18204;
  wire n_18205, n_18206, n_18207, n_18208, n_18209, n_18210, n_18211,
       n_18212;
  wire n_18213, n_18214, n_18215, n_18220, n_18221, n_18222, n_18223,
       n_18224;
  wire n_18225, n_18226, n_18227, n_18232, n_18233, n_18234, n_18235,
       n_18240;
  wire n_18241, n_18242, n_18243, n_18248, n_18249, n_18250, n_18251,
       n_18252;
  wire n_18253, n_18254, n_18255, n_18256, n_18257, n_18258, n_18259,
       n_18260;
  wire n_18261, n_18262, n_18263, n_18264, n_18265, n_18266, n_18267,
       n_18268;
  wire n_18269, n_18270, n_18271, n_18272, n_18273, n_18274, n_18275,
       n_18276;
  wire n_18277, n_18278, n_18279, n_18280, n_18281, n_18282, n_18287,
       n_18288;
  wire n_18289, n_18290, n_18291, n_18292, n_18293, n_18294, n_18295,
       n_18296;
  wire n_18297, n_18298, n_18303, n_18304, n_18305, n_18306, n_18307,
       n_18308;
  wire n_18309, n_18310, n_18311, n_18312, n_18313, n_18314, n_18315,
       n_18320;
  wire n_18321, n_18322, n_18323, n_18324, n_18325, n_18326, n_18327,
       n_18328;
  wire n_18329, n_18330, n_18331, n_18332, n_18333, n_18334, n_18335,
       n_18336;
  wire n_18337, n_18338, n_18339, n_18340, n_18341, n_18342, n_18343,
       n_18344;
  wire n_18345, n_18346, n_18347, n_18352, n_18353, n_18354, n_18355,
       n_18356;
  wire n_18357, n_18358, n_18359, n_18360, n_18361, n_18362, n_18363,
       n_18368;
  wire n_18369, n_18370, n_18371, n_18372, n_18373, n_18374, n_18375,
       n_18376;
  wire n_18377, n_18378, n_18379, n_18384, n_18385, n_18386, n_18387,
       n_18388;
  wire n_18389, n_18390, n_18391, n_18392, n_18393, n_18394, n_18395,
       n_18396;
  wire n_18397, n_18398, n_18399, n_18400, n_18401, n_18402, n_18403,
       n_18404;
  wire n_18405, n_18406, n_18407, n_18408, n_18409, n_18410, n_18411,
       n_18412;
  wire n_18413, n_18414, n_18415, n_18416, n_18417, n_18418, n_18419,
       n_18420;
  wire n_18421, n_18422, n_18423, n_18424, n_18429, n_18430, n_18431,
       n_18432;
  wire n_18433, n_18434, n_18435, n_18436, n_18441, n_18442, n_18443,
       n_18444;
  wire n_18445, n_18446, n_18447, n_18448, n_18449, n_18450, n_18455,
       n_18456;
  wire n_18457, n_18458, n_18459, n_18460, n_18461, n_18462, n_18467,
       n_18468;
  wire n_18469, n_18470, n_18475, n_18476, n_18477, n_18478, n_18483,
       n_18484;
  wire n_18485, n_18486, n_18487, n_18488, n_18489, n_18490, n_18491,
       n_18492;
  wire n_18493, n_18494, n_18495, n_18496, n_18497, n_18498, n_18499,
       n_18500;
  wire n_18501, n_18502, n_18503, n_18504, n_18505, n_18506, n_18507,
       n_18508;
  wire n_18513, n_18514, n_18515, n_18516, n_18517, n_18518, n_18519,
       n_18520;
  wire n_18521, n_18522, n_18523, n_18524, n_18529, n_18530, n_18531,
       n_18532;
  wire n_18533, n_18534, n_18535, n_18536, n_18537, n_18538, n_18539,
       n_18540;
  wire n_18541, n_18542, n_18543, n_18544, n_18545, n_18546, n_18547,
       n_18548;
  wire n_18553, n_18554, n_18555, n_18556, n_18557, n_18558, n_18559,
       n_18560;
  wire n_18561, n_18562, n_18563, n_18564, n_18565, n_18570, n_18571,
       n_18572;
  wire n_18573, n_18574, n_18575, n_18576, n_18577, n_18578, n_18579,
       n_18580;
  wire n_18581, n_18582, n_18583, n_18584, n_18585, n_18586, n_18587,
       n_18588;
  wire n_18589, n_18594, n_18595, n_18596, n_18597, n_18598, n_18599,
       n_18600;
  wire n_18601, n_18602, n_18603, n_18604, n_18605, n_18610, n_18611,
       n_18612;
  wire n_18613, n_18614, n_18615, n_18616, n_18617, n_18618, n_18619,
       n_18620;
  wire n_18621, n_18622, n_18623, n_18624, n_18625, n_18626, n_18627,
       n_18628;
  wire n_18629, n_18630, n_18631, n_18632, n_18633, n_18634, n_18635,
       n_18636;
  wire n_18637, n_18638, n_18639, n_18640, n_18641, n_18642, n_18643,
       n_18644;
  wire n_18645, n_18646, n_18647, n_18648, n_18649, n_18650, n_18651,
       n_18652;
  wire n_18657, n_18658, n_18659, n_18660, n_18661, n_18662, n_18663,
       n_18664;
  wire n_18665, n_18666, n_18671, n_18672, n_18673, n_18674, n_18675,
       n_18676;
  wire n_18677, n_18678, n_18683, n_18684, n_18685, n_18686, n_18687,
       n_18688;
  wire n_18689, n_18690, n_18691, n_18696, n_18697, n_18698, n_18699,
       n_18700;
  wire n_18701, n_18702, n_18703, n_18704, n_18705, n_18706, n_18707,
       n_18712;
  wire n_18713, n_18714, n_18715, n_18716, n_18717, n_18718, n_18719,
       n_18720;
  wire n_18721, n_18722, n_18723, n_18728, n_18729, n_18730, n_18731,
       n_18732;
  wire n_18733, n_18734, n_18735, n_18736, n_18737, n_18738, n_18739,
       n_18744;
  wire n_18745, n_18746, n_18747, n_18748, n_18749, n_18750, n_18751,
       n_18752;
  wire n_18753, n_18754, n_18755, n_18756, n_18757, n_18758, n_18759,
       n_18760;
  wire n_18761, n_18762, n_18763, n_18768, n_18769, n_18770, n_18771,
       n_18772;
  wire n_18773, n_18774, n_18775, n_18776, n_18777, n_18778, n_18779,
       n_18784;
  wire n_18785, n_18786, n_18787, n_18788, n_18789, n_18790, n_18791,
       n_18792;
  wire n_18793, n_18794, n_18795, n_18800, n_18801, n_18802, n_18803,
       n_18804;
  wire n_18805, n_18806, n_18807, n_18808, n_18809, n_18810, n_18811,
       n_18816;
  wire n_18817, n_18818, n_18819, n_18820, n_18821, n_18822, n_18823,
       n_18824;
  wire n_18825, n_18826, n_18827, n_18832, n_18833, n_18834, n_18835,
       n_18836;
  wire n_18837, n_18838, n_18839, n_18840, n_18841, n_18842, n_18843,
       n_18848;
  wire n_18849, n_18850, n_18851, n_18852, n_18853, n_18854, n_18855,
       n_18856;
  wire n_18857, n_18858, n_18859, n_18860, n_18861, n_18862, n_18863,
       n_18864;
  wire n_18865, n_18866, n_18867, n_18868, n_18869, n_18870, n_18871,
       n_18872;
  wire n_18873, n_18874, n_18875, n_18876, n_18877, n_18878, n_18879,
       n_18880;
  wire n_18881, n_18886, n_18887, n_18888, n_18889, n_18890, n_18891,
       n_18892;
  wire n_18893, n_18894, n_18895, n_18896, n_18897, n_18898, n_18899,
       n_18900;
  wire n_18901, n_18902, n_18903, n_18904, n_18905, n_18906, n_18911,
       n_18912;
  wire n_18913, n_18914, n_18919, n_18920, n_18921, n_18922, n_18923,
       n_18924;
  wire n_18925, n_18926, n_18927, n_18928, n_18929, n_18930, n_18931,
       n_18932;
  wire n_18933, n_18934, n_18935, n_18936, n_18937, n_18938, n_18939,
       n_18940;
  wire n_18941, n_18942, n_18943, n_18944, n_18945, n_18946, n_18951,
       n_18952;
  wire n_18953, n_18954, n_18955, n_18956, n_18957, n_18958, n_18959,
       n_18960;
  wire n_18961, n_18962, n_18967, n_18968, n_18969, n_18970, n_18971,
       n_18972;
  wire n_18973, n_18974, n_18975, n_18976, n_18977, n_18978, n_18983,
       n_18984;
  wire n_18985, n_18986, n_18987, n_18988, n_18989, n_18990, n_18991,
       n_18992;
  wire n_18993, n_18994, n_18995, n_18996, n_18997, n_18998, n_18999,
       n_19000;
  wire n_19001, n_19002, n_19003, n_19004, n_19005, n_19006, n_19007,
       n_19008;
  wire n_19009, n_19010, n_19011, n_19016, n_19017, n_19018, n_19019,
       n_19020;
  wire n_19021, n_19022, n_19023, n_19024, n_19025, n_19026, n_19027,
       n_19032;
  wire n_19033, n_19034, n_19035, n_19036, n_19037, n_19038, n_19039,
       n_19040;
  wire n_19041, n_19042, n_19043, n_19048, n_19049, n_19050, n_19051,
       n_19052;
  wire n_19053, n_19054, n_19055, n_19056, n_19057, n_19058, n_19059,
       n_19064;
  wire n_19065, n_19066, n_19067, n_19068, n_19069, n_19070, n_19071,
       n_19072;
  wire n_19073, n_19074, n_19075, n_19076, n_19077, n_19078, n_19079,
       n_19080;
  wire n_19081, n_19082, n_19083, n_19084, n_19085, n_19086, n_19087,
       n_19088;
  wire n_19089, n_19090, n_19091, n_19092, n_19093, n_19094, n_19095,
       n_19096;
  wire n_19097, n_19098, n_19099, n_19100, n_19101, n_19102, n_19103,
       n_19104;
  wire n_19105, n_19106, n_19107, n_19108, n_19109, n_19110, n_19111,
       n_19112;
  wire n_19113, n_19114, n_19115, n_19120, n_19121, n_19122, n_19123,
       n_19124;
  wire n_19125, n_19126, n_19127, n_19132, n_19133, n_19134, n_19135,
       n_19136;
  wire n_19137, n_19138, n_19139, n_19140, n_19145, n_19146, n_19147,
       n_19148;
  wire n_19153, n_19154, n_19155, n_19156, n_19161, n_19162, n_19163,
       n_19164;
  wire n_19169, n_19170, n_19171, n_19172, n_19177, n_19178, n_19179,
       n_19180;
  wire n_19181, n_19182, n_19183, n_19184, n_19185, n_19186, n_19187,
       n_19188;
  wire n_19189, n_19190, n_19191, n_19192, n_19193, n_19194, n_19195,
       n_19196;
  wire n_19197, n_19198, n_19199, n_19200, n_19201, n_19202, n_19203,
       n_19204;
  wire n_19205, n_19206, n_19207, n_19208, n_19209, n_19210, n_19211,
       n_19212;
  wire n_19213, n_19214, n_19215, n_19216, n_19217, n_19218, n_19223,
       n_19224;
  wire n_19225, n_19226, n_19227, n_19228, n_19229, n_19230, n_19231,
       n_19232;
  wire n_19233, n_19234, n_19235, n_19240, n_19241, n_19242, n_19243,
       n_19244;
  wire n_19245, n_19246, n_19247, n_19248, n_19249, n_19250, n_19251,
       n_19252;
  wire n_19253, n_19254, n_19255, n_19256, n_19257, n_19258, n_19259,
       n_19264;
  wire n_19265, n_19266, n_19267, n_19268, n_19269, n_19270, n_19271,
       n_19272;
  wire n_19273, n_19274, n_19275, n_19280, n_19281, n_19282, n_19283,
       n_19284;
  wire n_19285, n_19286, n_19287, n_19288, n_19289, n_19290, n_19291,
       n_19292;
  wire n_19293, n_19294, n_19295, n_19296, n_19297, n_19298, n_19299,
       n_19300;
  wire n_19301, n_19302, n_19303, n_19304, n_19305, n_19306, n_19307,
       n_19308;
  wire n_19309, n_19310, n_19311, n_19312, n_19313, n_19314, n_19315,
       n_19316;
  wire n_19317, n_19318, n_19319, n_19320, n_19321, n_19322, n_19323,
       n_19328;
  wire n_19329, n_19330, n_19331, n_19332, n_19333, n_19334, n_19335,
       n_19336;
  wire n_19341, n_19342, n_19343, n_19344, n_19345, n_19350, n_19351,
       n_19352;
  wire n_19353, n_19354, n_19355, n_19356, n_19357, n_19358, n_19359,
       n_19360;
  wire n_19361, n_19362, n_19363, n_19364, n_19365, n_19366, n_19367,
       n_19368;
  wire n_19369, n_19374, n_19375, n_19376, n_19377, n_19378, n_19379,
       n_19380;
  wire n_19381, n_19382, n_19383, n_19384, n_19385, n_19390, n_19391,
       n_19392;
  wire n_19393, n_19394, n_19395, n_19396, n_19397, n_19398, n_19399,
       n_19400;
  wire n_19401, n_19406, n_19407, n_19408, n_19409, n_19410, n_19411,
       n_19412;
  wire n_19413, n_19414, n_19415, n_19416, n_19417, n_19422, n_19423,
       n_19424;
  wire n_19425, n_19426, n_19427, n_19428, n_19429, n_19430, n_19431,
       n_19432;
  wire n_19433, n_19438, n_19439, n_19440, n_19441, n_19442, n_19443,
       n_19444;
  wire n_19445, n_19446, n_19447, n_19448, n_19449, n_19454, n_19455,
       n_19456;
  wire n_19457, n_19458, n_19459, n_19460, n_19461, n_19462, n_19463,
       n_19464;
  wire n_19465, n_19470, n_19471, n_19472, n_19473, n_19474, n_19475,
       n_19476;
  wire n_19477, n_19478, n_19479, n_19480, n_19481, n_19486, n_19487,
       n_19488;
  wire n_19489, n_19490, n_19491, n_19492, n_19493, n_19494, n_19495,
       n_19496;
  wire n_19497, n_19498, n_19499, n_19500, n_19501, n_19502, n_19503,
       n_19504;
  wire n_19505, n_19510, n_19511, n_19512, n_19513, n_19514, n_19515,
       n_19516;
  wire n_19517, n_19518, n_19519, n_19520, n_19521, n_19522, n_19523,
       n_19524;
  wire n_19525, n_19526, n_19527, n_19528, n_19529, n_19530, n_19531,
       n_19532;
  wire n_19533, n_19534, n_19535, n_19536, n_19537, n_19538, n_19539,
       n_19540;
  wire n_19541, n_19542, n_19543, n_19544, n_19545, n_19550, n_19551,
       n_19552;
  wire n_19553, n_19554, n_19555, n_19556, n_19557, n_19562, n_19563,
       n_19564;
  wire n_19565, n_19570, n_19571, n_19572, n_19573, n_19578, n_19579,
       n_19580;
  wire n_19581, n_19586, n_19587, n_19588, n_19589, n_19590, n_19591,
       n_19592;
  wire n_19593, n_19594, n_19595, n_19600, n_19601, n_19602, n_19603,
       n_19604;
  wire n_19605, n_19606, n_19607, n_19608, n_19609, n_19610, n_19611,
       n_19612;
  wire n_19613, n_19614, n_19615, n_19616, n_19617, n_19618, n_19619,
       n_19620;
  wire n_19625, n_19626, n_19627, n_19628, n_19629, n_19630, n_19631,
       n_19632;
  wire n_19633, n_19634, n_19635, n_19636, n_19637, n_19638, n_19639,
       n_19640;
  wire n_19641, n_19642, n_19643, n_19644, n_19645, n_19646, n_19647,
       n_19648;
  wire n_19649, n_19650, n_19651, n_19652, n_19653, n_19654, n_19659,
       n_19660;
  wire n_19661, n_19662, n_19663, n_19664, n_19665, n_19666, n_19667,
       n_19668;
  wire n_19669, n_19670, n_19675, n_19676, n_19677, n_19678, n_19679,
       n_19680;
  wire n_19681, n_19682, n_19683, n_19684, n_19685, n_19686, n_19691,
       n_19692;
  wire n_19693, n_19694, n_19695, n_19696, n_19697, n_19698, n_19699,
       n_19700;
  wire n_19701, n_19702, n_19707, n_19708, n_19709, n_19710, n_19711,
       n_19712;
  wire n_19713, n_19714, n_19715, n_19716, n_19717, n_19718, n_19719,
       n_19720;
  wire n_19721, n_19722, n_19723, n_19724, n_19725, n_19726, n_19727,
       n_19728;
  wire n_19729, n_19730, n_19731, n_19732, n_19733, n_19734, n_19735,
       n_19736;
  wire n_19737, n_19738, n_19739, n_19740, n_19741, n_19742, n_19743,
       n_19744;
  wire n_19745, n_19746, n_19747, n_19748, n_19753, n_19754, n_19755,
       n_19756;
  wire n_19757, n_19758, n_19759, n_19760, n_19761, n_19766, n_19767,
       n_19768;
  wire n_19769, n_19774, n_19775, n_19776, n_19777, n_19782, n_19783,
       n_19784;
  wire n_19785, n_19790, n_19791, n_19792, n_19793, n_19794, n_19795,
       n_19796;
  wire n_19797, n_19798, n_19799, n_19800, n_19801, n_19802, n_19807,
       n_19808;
  wire n_19809, n_19810, n_19811, n_19812, n_19813, n_19814, n_19815,
       n_19816;
  wire n_19817, n_19818, n_19819, n_19820, n_19821, n_19822, n_19827,
       n_19828;
  wire n_19829, n_19830, n_19831, n_19832, n_19833, n_19834, n_19835,
       n_19836;
  wire n_19837, n_19838, n_19839, n_19840, n_19845, n_19846, n_19847,
       n_19848;
  wire n_19849, n_19850, n_19851, n_19852, n_19853, n_19854, n_19855,
       n_19856;
  wire n_19857, n_19858, n_19859, n_19860, n_19861, n_19862, n_19863,
       n_19864;
  wire n_19869, n_19870, n_19871, n_19872, n_19873, n_19874, n_19875,
       n_19876;
  wire n_19877, n_19878, n_19879, n_19880, n_19885, n_19886, n_19887,
       n_19888;
  wire n_19889, n_19890, n_19891, n_19892, n_19893, n_19894, n_19895,
       n_19896;
  wire n_19897, n_19898, n_19899, n_19900, n_19901, n_19902, n_19903,
       n_19904;
  wire n_19905, n_19906, n_19907, n_19908, n_19909, n_19910, n_19911,
       n_19912;
  wire n_19917, n_19918, n_19919, n_19920, n_19921, n_19922, n_19923,
       n_19924;
  wire n_19925, n_19926, n_19927, n_19928, n_19929, n_19930, n_19931,
       n_19932;
  wire n_19933, n_19934, n_19935, n_19936, n_19937, n_19938, n_19939,
       n_19940;
  wire n_19945, n_19946, n_19947, n_19948, n_19949, n_19954, n_19955,
       n_19956;
  wire n_19957, n_19958, n_19959, n_19960, n_19961, n_19962, n_19963,
       n_19964;
  wire n_19965, n_19966, n_19967, n_19968, n_19969, n_19970, n_19971,
       n_19976;
  wire n_19977, n_19978, n_19979, n_19980, n_19981, n_19982, n_19983,
       n_19988;
  wire n_19989, n_19990, n_19991, n_19992, n_19993, n_19994, n_19995,
       n_19996;
  wire n_19997, n_19998, n_19999, n_20000, n_20001, n_20002, n_20003,
       n_20004;
  wire n_20005, n_20006, n_20007, n_20012, n_20013, n_20014, n_20015,
       n_20016;
  wire n_20017, n_20018, n_20019, n_20020, n_20021, n_20022, n_20023,
       n_20028;
  wire n_20029, n_20030, n_20031, n_20032, n_20033, n_20034, n_20035,
       n_20036;
  wire n_20037, n_20038, n_20039, n_20044, n_20045, n_20046, n_20047,
       n_20048;
  wire n_20049, n_20050, n_20051, n_20052, n_20053, n_20054, n_20055,
       n_20060;
  wire n_20061, n_20062, n_20063, n_20064, n_20065, n_20066, n_20067,
       n_20068;
  wire n_20069, n_20070, n_20071, n_20076, n_20077, n_20078, n_20079,
       n_20080;
  wire n_20081, n_20082, n_20083, n_20084, n_20085, n_20086, n_20087,
       n_20088;
  wire n_20089, n_20090, n_20091, n_20092, n_20093, n_20094, n_20095,
       n_20100;
  wire n_20101, n_20102, n_20103, n_20104, n_20105, n_20106, n_20107,
       n_20108;
  wire n_20109, n_20110, n_20111, n_20116, n_20117, n_20118, n_20119,
       n_20120;
  wire n_20121, n_20122, n_20123, n_20124, n_20125, n_20126, n_20127,
       n_20128;
  wire n_20129, n_20130, n_20131, n_20132, n_20133, n_20134, n_20135,
       n_20136;
  wire n_20137, n_20138, n_20139, n_20140, n_20141, n_20142, n_20143,
       n_20144;
  wire n_20145, n_20146, n_20147, n_20152, n_20153, n_20154, n_20155,
       n_20160;
  wire n_20161, n_20162, n_20163, n_20168, n_20169, n_20170, n_20171,
       n_20176;
  wire n_20177, n_20178, n_20179, n_20180, n_20181, n_20182, n_20183,
       n_20184;
  wire n_20185, n_20186, n_20191, n_20192, n_20193, n_20194, n_20195,
       n_20196;
  wire n_20197, n_20198, n_20199, n_20200, n_20201, n_20202, n_20203,
       n_20204;
  wire n_20205, n_20206, n_20207, n_20208, n_20209, n_20210, n_20211,
       n_20212;
  wire n_20213, n_20214, n_20215, n_20216, n_20217, n_20218, n_20219,
       n_20220;
  wire n_20221, n_20222, n_20223, n_20224, n_20225, n_20226, n_20227,
       n_20232;
  wire n_20233, n_20234, n_20235, n_20236, n_20237, n_20238, n_20239,
       n_20240;
  wire n_20241, n_20242, n_20243, n_20248, n_20249, n_20250, n_20251,
       n_20252;
  wire n_20253, n_20254, n_20255, n_20256, n_20257, n_20258, n_20259,
       n_20264;
  wire n_20265, n_20266, n_20267, n_20268, n_20269, n_20270, n_20271,
       n_20272;
  wire n_20273, n_20274, n_20275, n_20280, n_20281, n_20282, n_20283,
       n_20284;
  wire n_20285, n_20286, n_20287, n_20288, n_20289, n_20290, n_20291,
       n_20292;
  wire n_20293, n_20294, n_20295, n_20296, n_20297, n_20298, n_20299,
       n_20304;
  wire n_20305, n_20306, n_20307, n_20308, n_20309, n_20310, n_20311,
       n_20312;
  wire n_20313, n_20314, n_20315, n_20316, n_20317, n_20318, n_20319,
       n_20320;
  wire n_20321, n_20322, n_20323, n_20324, n_20325, n_20326, n_20327,
       n_20328;
  wire n_20329, n_20330, n_20331, n_20332, n_20333, n_20334, n_20335,
       n_20340;
  wire n_20341, n_20342, n_20343, n_20348, n_20349, n_20350, n_20351,
       n_20356;
  wire n_20357, n_20358, n_20359, n_20364, n_20365, n_20366, n_20367,
       n_20368;
  wire n_20369, n_20370, n_20371, n_20372, n_20373, n_20374, n_20375,
       n_20376;
  wire n_20381, n_20382, n_20383, n_20384, n_20385, n_20386, n_20387,
       n_20388;
  wire n_20389, n_20394, n_20395, n_20396, n_20397, n_20398, n_20399,
       n_20400;
  wire n_20401, n_20402, n_20403, n_20404, n_20405, n_20406, n_20407,
       n_20408;
  wire n_20409, n_20410, n_20411, n_20412, n_20413, n_20414, n_20415,
       n_20416;
  wire n_20417, n_20418, n_20419, n_20420, n_20421, n_20426, n_20427,
       n_20428;
  wire n_20429, n_20430, n_20431, n_20432, n_20433, n_20434, n_20435,
       n_20436;
  wire n_20437, n_20442, n_20443, n_20444, n_20445, n_20446, n_20447,
       n_20448;
  wire n_20449, n_20450, n_20451, n_20452, n_20453, n_20454, n_20455,
       n_20456;
  wire n_20457, n_20458, n_20459, n_20460, n_20461, n_20462, n_20463,
       n_20464;
  wire n_20465, n_20466, n_20467, n_20468, n_20469, n_20474, n_20475,
       n_20476;
  wire n_20477, n_20478, n_20479, n_20480, n_20481, n_20482, n_20483,
       n_20484;
  wire n_20485, n_20490, n_20491, n_20492, n_20493, n_20494, n_20495,
       n_20496;
  wire n_20497, n_20498, n_20499, n_20500, n_20501, n_20502, n_20503,
       n_20504;
  wire n_20505, n_20506, n_20507, n_20508, n_20509, n_20510, n_20511,
       n_20516;
  wire n_20517, n_20518, n_20519, n_20524, n_20525, n_20526, n_20527,
       n_20528;
  wire n_20529, n_20530, n_20531, n_20532, n_20533, n_20534, n_20535,
       n_20536;
  wire n_20537, n_20538, n_20539, n_20540, n_20541, n_20546, n_20547,
       n_20548;
  wire n_20549, n_20550, n_20551, n_20552, n_20553, n_20558, n_20559,
       n_20560;
  wire n_20561, n_20562, n_20563, n_20564, n_20565, n_20566, n_20567,
       n_20568;
  wire n_20569, n_20570, n_20571, n_20572, n_20573, n_20574, n_20575,
       n_20576;
  wire n_20577, n_20582, n_20583, n_20584, n_20585, n_20586, n_20587,
       n_20588;
  wire n_20589, n_20590, n_20591, n_20592, n_20593, n_20598, n_20599,
       n_20600;
  wire n_20601, n_20602, n_20603, n_20604, n_20605, n_20606, n_20607,
       n_20608;
  wire n_20609, n_20614, n_20615, n_20616, n_20617, n_20618, n_20619,
       n_20620;
  wire n_20621, n_20622, n_20623, n_20624, n_20625, n_20630, n_20631,
       n_20632;
  wire n_20633, n_20634, n_20635, n_20636, n_20637, n_20638, n_20639,
       n_20640;
  wire n_20641, n_20642, n_20643, n_20644, n_20645, n_20646, n_20647,
       n_20648;
  wire n_20649, n_20654, n_20655, n_20656, n_20657, n_20658, n_20659,
       n_20660;
  wire n_20661, n_20662, n_20663, n_20664, n_20665, n_20670, n_20671,
       n_20672;
  wire n_20673, n_20674, n_20675, n_20676, n_20677, n_20678, n_20679,
       n_20680;
  wire n_20681, n_20682, n_20683, n_20684, n_20685, n_20686, n_20687,
       n_20688;
  wire n_20689, n_20690, n_20691, n_20692, n_20693, n_20694, n_20695,
       n_20696;
  wire n_20697, n_20698, n_20699, n_20700, n_20701, n_20702, n_20707,
       n_20708;
  wire n_20709, n_20710, n_20715, n_20716, n_20717, n_20718, n_20723,
       n_20724;
  wire n_20725, n_20726, n_20727, n_20728, n_20729, n_20730, n_20731,
       n_20732;
  wire n_20733, n_20738, n_20739, n_20740, n_20741, n_20742, n_20743,
       n_20744;
  wire n_20745, n_20746, n_20747, n_20748, n_20749, n_20750, n_20751,
       n_20752;
  wire n_20753, n_20754, n_20755, n_20756, n_20757, n_20758, n_20759,
       n_20760;
  wire n_20761, n_20762, n_20763, n_20764, n_20765, n_20770, n_20771,
       n_20772;
  wire n_20773, n_20774, n_20775, n_20776, n_20777, n_20778, n_20779,
       n_20780;
  wire n_20781, n_20786, n_20787, n_20788, n_20789, n_20790, n_20791,
       n_20792;
  wire n_20793, n_20794, n_20795, n_20796, n_20797, n_20802, n_20803,
       n_20804;
  wire n_20805, n_20806, n_20807, n_20808, n_20809, n_20810, n_20811,
       n_20812;
  wire n_20813, n_20818, n_20819, n_20820, n_20821, n_20822, n_20823,
       n_20824;
  wire n_20825, n_20826, n_20827, n_20828, n_20829, n_20830, n_20831,
       n_20832;
  wire n_20833, n_20834, n_20835, n_20836, n_20837, n_20842, n_20843,
       n_20844;
  wire n_20845, n_20846, n_20847, n_20848, n_20849, n_20850, n_20851,
       n_20852;
  wire n_20853, n_20854, n_20855, n_20856, n_20857, n_20858, n_20859,
       n_20860;
  wire n_20861, n_20862, n_20863, n_20864, n_20865, n_20866, n_20867,
       n_20868;
  wire n_20869, n_20870, n_20871, n_20872, n_20873, n_20878, n_20879,
       n_20880;
  wire n_20881, n_20886, n_20887, n_20888, n_20889, n_20894, n_20895,
       n_20896;
  wire n_20897, n_20898, n_20899, n_20900, n_20901, n_20902, n_20903,
       n_20904;
  wire n_20905, n_20906, n_20911, n_20912, n_20913, n_20914, n_20915,
       n_20916;
  wire n_20917, n_20918, n_20919, n_20924, n_20925, n_20926, n_20927,
       n_20928;
  wire n_20929, n_20930, n_20931, n_20932, n_20933, n_20934, n_20935,
       n_20936;
  wire n_20937, n_20938, n_20939, n_20940, n_20941, n_20942, n_20943,
       n_20948;
  wire n_20949, n_20950, n_20951, n_20952, n_20953, n_20954, n_20955,
       n_20956;
  wire n_20957, n_20958, n_20959, n_20964, n_20965, n_20966, n_20967,
       n_20968;
  wire n_20969, n_20970, n_20971, n_20972, n_20973, n_20974, n_20975,
       n_20976;
  wire n_20977, n_20978, n_20979, n_20980, n_20981, n_20982, n_20983,
       n_20984;
  wire n_20985, n_20986, n_20987, n_20988, n_20989, n_20990, n_20991,
       n_20996;
  wire n_20997, n_20998, n_20999, n_21000, n_21001, n_21002, n_21003,
       n_21004;
  wire n_21005, n_21006, n_21007, n_21012, n_21013, n_21014, n_21015,
       n_21016;
  wire n_21017, n_21018, n_21019, n_21020, n_21021, n_21022, n_21023,
       n_21024;
  wire n_21025, n_21026, n_21027, n_21028, n_21029, n_21030, n_21031,
       n_21036;
  wire n_21037, n_21038, n_21039, n_21040, n_21041, n_21042, n_21043,
       n_21044;
  wire n_21045, n_21046, n_21047, n_21048, n_21049, n_21050, n_21051,
       n_21056;
  wire n_21057, n_21058, n_21059, n_21060, n_21061, n_21062, n_21063,
       n_21068;
  wire n_21069, n_21070, n_21071, n_21072, n_21073, n_21074, n_21075,
       n_21076;
  wire n_21077, n_21078, n_21079, n_21080, n_21081, n_21086, n_21087,
       n_21088;
  wire n_21089, n_21090, n_21091, n_21092, n_21093, n_21094, n_21095,
       n_21096;
  wire n_21097, n_21098, n_21103, n_21104, n_21105, n_21106, n_21107,
       n_21108;
  wire n_21109, n_21110, n_21111, n_21112, n_21113, n_21114, n_21119,
       n_21120;
  wire n_21121, n_21122, n_21123, n_21124, n_21125, n_21126, n_21127,
       n_21128;
  wire n_21129, n_21130, n_21131, n_21132, n_21133, n_21134, n_21135,
       n_21136;
  wire n_21137, n_21138, n_21143, n_21144, n_21145, n_21146, n_21147,
       n_21148;
  wire n_21149, n_21150, n_21151, n_21152, n_21153, n_21154, n_21159,
       n_21160;
  wire n_21161, n_21162, n_21163, n_21164, n_21165, n_21166, n_21167,
       n_21168;
  wire n_21169, n_21170, n_21175, n_21176, n_21177, n_21178, n_21179,
       n_21180;
  wire n_21181, n_21182, n_21183, n_21184, n_21185, n_21186, n_21187,
       n_21188;
  wire n_21189, n_21190, n_21191, n_21192, n_21193, n_21194, n_21195,
       n_21196;
  wire n_21197, n_21198, n_21199, n_21200, n_21201, n_21202, n_21203,
       n_21204;
  wire n_21205, n_21206, n_21207, n_21212, n_21213, n_21214, n_21215,
       n_21216;
  wire n_21217, n_21218, n_21219, n_21220, n_21221, n_21222, n_21223,
       n_21224;
  wire n_21225, n_21226, n_21227, n_21228, n_21229, n_21230, n_21231,
       n_21236;
  wire n_21237, n_21238, n_21239, n_21240, n_21241, n_21242, n_21243,
       n_21244;
  wire n_21245, n_21246, n_21247, n_21252, n_21253, n_21254, n_21255,
       n_21256;
  wire n_21257, n_21258, n_21259, n_21260, n_21261, n_21262, n_21263,
       n_21268;
  wire n_21269, n_21270, n_21271, n_21272, n_21273, n_21274, n_21275,
       n_21276;
  wire n_21277, n_21278, n_21279, n_21284, n_21285, n_21286, n_21287,
       n_21288;
  wire n_21289, n_21290, n_21291, n_21292, n_21293, n_21294, n_21295,
       n_21296;
  wire n_21301, n_21302, n_21303, n_21304, n_21305, n_21306, n_21307,
       n_21308;
  wire n_21309, n_21310, n_21311, n_21312, n_21313, n_21318, n_21319,
       n_21320;
  wire n_21321, n_21322, n_21323, n_21324, n_21325, n_21326, n_21327,
       n_21328;
  wire n_21329, n_21334, n_21335, n_21336, n_21337, n_21338, n_21339,
       n_21340;
  wire n_21341, n_21342, n_21343, n_21344, n_21345, n_21346, n_21347,
       n_21348;
  wire n_21349, n_21350, n_21351, n_21352, n_21353, n_21354, n_21355,
       n_21356;
  wire n_21357, n_21358, n_21359, n_21360, n_21361, n_21362, n_21363,
       n_21368;
  wire n_21369, n_21370, n_21371, n_21376, n_21377, n_21378, n_21379,
       n_21380;
  wire n_21381, n_21382, n_21383, n_21384, n_21385, n_21386, n_21387,
       n_21388;
  wire n_21389, n_21390, n_21395, n_21396, n_21397, n_21398, n_21399,
       n_21400;
  wire n_21401, n_21402, n_21403, n_21408, n_21409, n_21410, n_21411,
       n_21412;
  wire n_21413, n_21414, n_21415, n_21416, n_21417, n_21418, n_21419,
       n_21424;
  wire n_21425, n_21426, n_21427, n_21428, n_21429, n_21430, n_21431,
       n_21432;
  wire n_21433, n_21434, n_21435, n_21440, n_21441, n_21442, n_21443,
       n_21444;
  wire n_21445, n_21446, n_21447, n_21448, n_21449, n_21450, n_21451,
       n_21452;
  wire n_21453, n_21454, n_21455, n_21456, n_21457, n_21458, n_21459,
       n_21460;
  wire n_21461, n_21462, n_21463, n_21464, n_21465, n_21466, n_21467,
       n_21472;
  wire n_21473, n_21474, n_21475, n_21476, n_21477, n_21478, n_21479,
       n_21480;
  wire n_21481, n_21482, n_21483, n_21488, n_21489, n_21490, n_21491,
       n_21492;
  wire n_21493, n_21494, n_21495, n_21496, n_21497, n_21498, n_21499,
       n_21500;
  wire n_21501, n_21502, n_21503, n_21504, n_21505, n_21506, n_21507,
       n_21512;
  wire n_21513, n_21514, n_21515, n_21516, n_21517, n_21518, n_21519,
       n_21520;
  wire n_21521, n_21522, n_21523, n_21524, n_21525, n_21526, n_21527,
       n_21528;
  wire n_21533, n_21534, n_21535, n_21536, n_21537, n_21538, n_21539,
       n_21540;
  wire n_21545, n_21546, n_21547, n_21548, n_21549, n_21550, n_21551,
       n_21552;
  wire n_21553, n_21554, n_21555, n_21556, n_21557, n_21558, n_21559,
       n_21564;
  wire n_21565, n_21566, n_21567, n_21568, n_21569, n_21570, n_21571,
       n_21572;
  wire n_21573, n_21574, n_21575, n_21576, n_21581, n_21582, n_21583,
       n_21584;
  wire n_21585, n_21586, n_21587, n_21588, n_21589, n_21590, n_21591,
       n_21592;
  wire n_21593, n_21594, n_21595, n_21596, n_21597, n_21598, n_21599,
       n_21600;
  wire n_21605, n_21606, n_21607, n_21608, n_21609, n_21610, n_21611,
       n_21612;
  wire n_21613, n_21614, n_21615, n_21616, n_21621, n_21622, n_21623,
       n_21624;
  wire n_21625, n_21626, n_21627, n_21628, n_21629, n_21630, n_21631,
       n_21632;
  wire n_21637, n_21638, n_21639, n_21640, n_21641, n_21642, n_21643,
       n_21644;
  wire n_21645, n_21646, n_21647, n_21648, n_21649, n_21650, n_21651,
       n_21652;
  wire n_21653, n_21654, n_21655, n_21656, n_21657, n_21658, n_21659,
       n_21660;
  wire n_21661, n_21662, n_21663, n_21664, n_21665, n_21666, n_21667,
       n_21668;
  wire n_21669, n_21670, n_21671, n_21672, n_21673, n_21674, n_21675,
       n_21676;
  wire n_21677, n_21678, n_21679, n_21680, n_21681, n_21682, n_21683,
       n_21684;
  wire n_21685, n_21686, n_21687, n_21688, n_21689, n_21690, n_21691,
       n_21692;
  wire n_21693, n_21698, n_21699, n_21700, n_21701, n_21702, n_21703,
       n_21704;
  wire n_21705, n_21706, n_21707, n_21708, n_21709, n_21714, n_21715,
       n_21716;
  wire n_21717, n_21718, n_21719, n_21720, n_21721, n_21722, n_21723,
       n_21724;
  wire n_21725, n_21730, n_21731, n_21732, n_21733, n_21734, n_21735,
       n_21736;
  wire n_21737, n_21738, n_21739, n_21740, n_21741, n_21742, n_21747,
       n_21748;
  wire n_21749, n_21750, n_21751, n_21752, n_21753, n_21754, n_21755,
       n_21756;
  wire n_21757, n_21758, n_21759, n_21764, n_21765, n_21766, n_21767,
       n_21768;
  wire n_21769, n_21770, n_21771, n_21772, n_21773, n_21774, n_21775,
       n_21780;
  wire n_21781, n_21782, n_21783, n_21784, n_21785, n_21786, n_21787,
       n_21788;
  wire n_21789, n_21790, n_21791, n_21792, n_21793, n_21794, n_21795,
       n_21796;
  wire n_21797, n_21798, n_21799, n_21800, n_21801, n_21802, n_21803,
       n_21804;
  wire n_21805, n_21806, n_21807, n_21808, n_21809, n_21814, n_21815,
       n_21816;
  wire n_21817, n_21822, n_21823, n_21824, n_21825, n_21830, n_21831,
       n_21832;
  wire n_21833, n_21834, n_21835, n_21836, n_21837, n_21838, n_21839,
       n_21840;
  wire n_21841, n_21842, n_21843, n_21844, n_21849, n_21850, n_21851,
       n_21852;
  wire n_21853, n_21854, n_21855, n_21856, n_21861, n_21862, n_21863,
       n_21864;
  wire n_21865, n_21866, n_21867, n_21868, n_21869, n_21870, n_21871,
       n_21872;
  wire n_21877, n_21878, n_21879, n_21880, n_21881, n_21882, n_21883,
       n_21884;
  wire n_21885, n_21886, n_21887, n_21888, n_21889, n_21890, n_21891,
       n_21892;
  wire n_21893, n_21894, n_21895, n_21896, n_21897, n_21898, n_21899,
       n_21900;
  wire n_21901, n_21902, n_21903, n_21904, n_21905, n_21906, n_21907,
       n_21908;
  wire n_21909, n_21910, n_21911, n_21912, n_21917, n_21918, n_21919,
       n_21920;
  wire n_21921, n_21922, n_21923, n_21924, n_21925, n_21926, n_21927,
       n_21928;
  wire n_21929, n_21930, n_21931, n_21932, n_21933, n_21934, n_21935,
       n_21936;
  wire n_21941, n_21942, n_21943, n_21944, n_21949, n_21950, n_21951,
       n_21952;
  wire n_21957, n_21958, n_21959, n_21960, n_21961, n_21962, n_21963,
       n_21964;
  wire n_21965, n_21966, n_21967, n_21968, n_21973, n_21974, n_21975,
       n_21976;
  wire n_21977, n_21978, n_21979, n_21980, n_21981, n_21982, n_21983,
       n_21984;
  wire n_21989, n_21990, n_21991, n_21992, n_21993, n_21994, n_21995,
       n_21996;
  wire n_21997, n_21998, n_21999, n_22000, n_22001, n_22002, n_22003,
       n_22004;
  wire n_22005, n_22006, n_22007, n_22008, n_22009, n_22010, n_22015,
       n_22016;
  wire n_22017, n_22018, n_22019, n_22020, n_22021, n_22022, n_22023,
       n_22024;
  wire n_22025, n_22026, n_22027, n_22028, n_22029, n_22030, n_22031,
       n_22032;
  wire n_22033, n_22034, n_22035, n_22036, n_22037, n_22038, n_22039,
       n_22040;
  wire n_22041, n_22042, n_22047, n_22048, n_22049, n_22050, n_22051,
       n_22052;
  wire n_22053, n_22054, n_22055, n_22056, n_22057, n_22058, n_22059,
       n_22060;
  wire n_22061, n_22062, n_22063, n_22064, n_22065, n_22066, n_22067,
       n_22068;
  wire n_22069, n_22070, n_22071, n_22072, n_22073, n_22074, n_22075,
       n_22076;
  wire n_22077, n_22078, n_22079, n_22084, n_22085, n_22086, n_22087,
       n_22088;
  wire n_22089, n_22090, n_22091, n_22092, n_22093, n_22094, n_22095,
       n_22096;
  wire n_22097, n_22098, n_22099, n_22100, n_22101, n_22102, n_22103,
       n_22104;
  wire n_22105, n_22106, n_22107, n_22108, n_22109, n_22110, n_22115,
       n_22116;
  wire n_22117, n_22118, n_22119, n_22120, n_22121, n_22122, n_22123,
       n_22124;
  wire n_22125, n_22126, n_22131, n_22132, n_22133, n_22134, n_22135,
       n_22136;
  wire n_22137, n_22138, n_22139, n_22140, n_22141, n_22142, n_22147,
       n_22148;
  wire n_22149, n_22150, n_22151, n_22152, n_22153, n_22154, n_22155,
       n_22156;
  wire n_22157, n_22158, n_22163, n_22164, n_22165, n_22166, n_22167,
       n_22168;
  wire n_22169, n_22170, n_22171, n_22172, n_22173, n_22174, n_22175,
       n_22176;
  wire n_22177, n_22178, n_22179, n_22180, n_22181, n_22182, n_22183,
       n_22184;
  wire n_22185, n_22186, n_22187, n_22188, n_22189, n_22190, n_22191,
       n_22192;
  wire n_22193, n_22194, n_22195, n_22196, n_22197, n_22198, n_22199,
       n_22200;
  wire n_22201, n_22202, n_22207, n_22208, n_22209, n_22210, n_22215,
       n_22216;
  wire n_22217, n_22218, n_22223, n_22224, n_22225, n_22226, n_22231,
       n_22232;
  wire n_22233, n_22234, n_22235, n_22236, n_22237, n_22238, n_22239,
       n_22240;
  wire n_22241, n_22242, n_22243, n_22244, n_22245, n_22246, n_22247,
       n_22248;
  wire n_22249, n_22250, n_22251, n_22252, n_22253, n_22254, n_22255,
       n_22256;
  wire n_22257, n_22258, n_22259, n_22260, n_22261, n_22262, n_22263,
       n_22264;
  wire n_22265, n_22266, n_22267, n_22268, n_22269, n_22270, n_22271,
       n_22272;
  wire n_22273, n_22274, n_22275, n_22276, n_22277, n_22278, n_22279,
       n_22280;
  wire n_22281, n_22282, n_22283, n_22284, n_22285, n_22286, n_22287,
       n_22288;
  wire n_22289, n_22290, n_22295, n_22296, n_22297, n_22298, n_22299,
       n_22300;
  wire n_22301, n_22302, n_22303, n_22304, n_22305, n_22306, n_22307,
       n_22308;
  wire n_22309, n_22310, n_22311, n_22312, n_22313, n_22314, n_22315,
       n_22320;
  wire n_22321, n_22322, n_22323, n_22328, n_22329, n_22330, n_22331,
       n_22336;
  wire n_22337, n_22338, n_22339, n_22344, n_22345, n_22346, n_22347,
       n_22348;
  wire n_22349, n_22350, n_22351, n_22352, n_22353, n_22354, n_22355,
       n_22356;
  wire n_22357, n_22358, n_22359, n_22360, n_22365, n_22366, n_22367,
       n_22368;
  wire n_22369, n_22370, n_22371, n_22372, n_22373, n_22378, n_22379,
       n_22380;
  wire n_22381, n_22382, n_22383, n_22384, n_22385, n_22386, n_22387,
       n_22388;
  wire n_22389, n_22390, n_22391, n_22392, n_22393, n_22394, n_22395,
       n_22396;
  wire n_22397, n_22398, n_22399, n_22400, n_22401, n_22402, n_22403,
       n_22404;
  wire n_22405, n_22406, n_22407, n_22408, n_22409, n_22410, n_22411,
       n_22412;
  wire n_22413, n_22414, n_22415, n_22416, n_22417, n_22418, n_22419,
       n_22420;
  wire n_22421, n_22422, n_22423, n_22424, n_22425, n_22426, n_22427,
       n_22428;
  wire n_22429, n_22430, n_22431, n_22432, n_22433, n_22434, n_22435,
       n_22436;
  wire n_22437, n_22438, n_22439, n_22440, n_22441, n_22442, n_22447,
       n_22448;
  wire n_22449, n_22450, n_22455, n_22456, n_22457, n_22458, n_22463,
       n_22464;
  wire n_22465, n_22466, n_22467, n_22468, n_22469, n_22470, n_22471,
       n_22472;
  wire n_22477, n_22478, n_22479, n_22480, n_22481, n_22482, n_22483,
       n_22484;
  wire n_22485, n_22486, n_22487, n_22488, n_22489, n_22490, n_22491,
       n_22492;
  wire n_22493, n_22494, n_22495, n_22496, n_22497, n_22498, n_22499,
       n_22500;
  wire n_22501, n_22502, n_22503, n_22504, n_22509, n_22510, n_22511,
       n_22512;
  wire n_22513, n_22514, n_22515, n_22516, n_22517, n_22518, n_22519,
       n_22520;
  wire n_22521, n_22522, n_22523, n_22524, n_22525, n_22526, n_22527,
       n_22528;
  wire n_22529, n_22530, n_22531, n_22532, n_22533, n_22534, n_22535,
       n_22536;
  wire n_22537, n_22542, n_22543, n_22544, n_22545, n_22550, n_22551,
       n_22552;
  wire n_22553, n_22558, n_22559, n_22560, n_22561, n_22562, n_22563,
       n_22564;
  wire n_22565, n_22566, n_22567, n_22568, n_22569, n_22570, n_22575,
       n_22576;
  wire n_22577, n_22578, n_22579, n_22580, n_22581, n_22582, n_22583,
       n_22584;
  wire n_22585, n_22586, n_22587, n_22588, n_22589, n_22590, n_22591,
       n_22592;
  wire n_22593, n_22594, n_22595, n_22596, n_22597, n_22598, n_22599,
       n_22600;
  wire n_22601, n_22602, n_22603, n_22604, n_22605, n_22606, n_22607,
       n_22608;
  wire n_22613, n_22614, n_22615, n_22616, n_22617, n_22618, n_22619,
       n_22620;
  wire n_22621, n_22622, n_22623, n_22624, n_22625, n_22626, n_22627,
       n_22628;
  wire n_22629, n_22630, n_22631, n_22632, n_22633, n_22634, n_22635,
       n_22636;
  wire n_22637, n_22638, n_22639, n_22640, n_22641, n_22642, n_22643,
       n_22648;
  wire n_22649, n_22650, n_22651, n_22656, n_22657, n_22658, n_22659,
       n_22664;
  wire n_22665, n_22666, n_22667, n_22668, n_22673, n_22674, n_22675,
       n_22676;
  wire n_22677, n_22678, n_22679, n_22680, n_22681, n_22682, n_22683,
       n_22684;
  wire n_22685, n_22686, n_22687, n_22688, n_22689, n_22690, n_22691,
       n_22692;
  wire n_22693, n_22698, n_22699, n_22700, n_22701, n_22702, n_22703,
       n_22704;
  wire n_22705, n_22706, n_22707, n_22708, n_22709, n_22710, n_22711,
       n_22712;
  wire n_22713, n_22714, n_22715, n_22716, n_22717, n_22718, n_22719,
       n_22720;
  wire n_22721, n_22722, n_22723, n_22724, n_22725, n_22726, n_22727,
       n_22728;
  wire n_22729, n_22730, n_22731, n_22732, n_22733, n_22734, n_22735,
       n_22736;
  wire n_22737, n_22738, n_22739, n_22740, n_22741, n_22742, n_22743,
       n_22744;
  wire n_22745, n_22746, n_22747, n_22748, n_22753, n_22754, n_22755,
       n_22756;
  wire n_22761, n_22762, n_22763, n_22764, n_22769, n_22770, n_22771,
       n_22772;
  wire n_22773, n_22774, n_22775, n_22776, n_22777, n_22778, n_22779,
       n_22780;
  wire n_22781, n_22782, n_22783, n_22784, n_22785, n_22786, n_22787,
       n_22788;
  wire n_22789, n_22790, n_22791, n_22792, n_22793, n_22794, n_22795,
       n_22796;
  wire n_22797, n_22798, n_22799, n_22800, n_22801, n_22802, n_22803,
       n_22804;
  wire n_22805, n_22806, n_22807, n_22808, n_22809, n_22810, n_22811,
       n_22812;
  wire n_22813, n_22814, n_22815, n_22816, n_22817, n_22818, n_22819,
       n_22820;
  wire n_22821, n_22822, n_22823, n_22824, n_22825, n_22826, n_22827,
       n_22828;
  wire n_22829, n_22830, n_22831, n_22836, n_22837, n_22838, n_22839,
       n_22844;
  wire n_22845, n_22846, n_22847, n_22848, n_22849, n_22850, n_22851,
       n_22852;
  wire n_22853, n_22854, n_22855, n_22856, n_22857, n_22858, n_22859,
       n_22860;
  wire n_22861, n_22862, n_22867, n_22868, n_22869, n_22870, n_22871,
       n_22872;
  wire n_22873, n_22874, n_22875, n_22876, n_22877, n_22878, n_22879,
       n_22880;
  wire n_22881, n_22882, n_22883, n_22884, n_22885, n_22886, n_22891,
       n_22892;
  wire n_22893, n_22894, n_22895, n_22896, n_22897, n_22898, n_22899,
       n_22900;
  wire n_22901, n_22902, n_22903, n_22904, n_22905, n_22906, n_22907,
       n_22908;
  wire n_22909, n_22910, n_22911, n_22912, n_22913, n_22914, n_22915,
       n_22916;
  wire n_22917, n_22918, n_22919, n_22920, n_22921, n_22926, n_22927,
       n_22928;
  wire n_22929, n_22934, n_22935, n_22936, n_22937, n_22942, n_22943,
       n_22944;
  wire n_22945, n_22946, n_22947, n_22948, n_22949, n_22950, n_22951,
       n_22952;
  wire n_22953, n_22954, n_22955, n_22956, n_22957, n_22958, n_22959,
       n_22960;
  wire n_22961, n_22962, n_22963, n_22964, n_22965, n_22966, n_22967,
       n_22968;
  wire n_22969, n_22970, n_22971, n_22972, n_22973, n_22974, n_22975,
       n_22976;
  wire n_22977, n_22982, n_22983, n_22984, n_22985, n_22986, n_22987,
       n_22988;
  wire n_22989, n_22990, n_22991, n_22992, n_22993, n_22994, n_22995,
       n_22996;
  wire n_22997, n_22998, n_22999, n_23000, n_23001, n_23002, n_23003,
       n_23004;
  wire n_23005, n_23006, n_23007, n_23008, n_23013, n_23014, n_23015,
       n_23016;
  wire n_23021, n_23022, n_23023, n_23024, n_23025, n_23026, n_23027,
       n_23028;
  wire n_23029, n_23030, n_23035, n_23036, n_23037, n_23038, n_23039,
       n_23040;
  wire n_23041, n_23042, n_23043, n_23044, n_23045, n_23046, n_23047,
       n_23048;
  wire n_23049, n_23050, n_23051, n_23052, n_23053, n_23054, n_23055,
       n_23056;
  wire n_23057, n_23058, n_23059, n_23060, n_23061, n_23062, n_23063,
       n_23064;
  wire n_23065, n_23066, n_23067, n_23068, n_23069, n_23070, n_23071,
       n_23072;
  wire n_23073, n_23074, n_23075, n_23076, n_23077, n_23078, n_23079,
       n_23080;
  wire n_23081, n_23082, n_23083, n_23088, n_23089, n_23090, n_23091,
       n_23092;
  wire n_23093, n_23094, n_23095, n_23100, n_23101, n_23102, n_23103,
       n_23104;
  wire n_23105, n_23106, n_23107, n_23108, n_23109, n_23110, n_23111,
       n_23116;
  wire n_23117, n_23118, n_23119, n_23120, n_23121, n_23122, n_23123,
       n_23124;
  wire n_23125, n_23126, n_23127, n_23128, n_23129, n_23130, n_23131,
       n_23132;
  wire n_23133, n_23134, n_23135, n_23136, n_23137, n_23138, n_23139,
       n_23140;
  wire n_23141, n_23142, n_23143, n_23144, n_23145, n_23146, n_23151,
       n_23152;
  wire n_23153, n_23154, n_23155, n_23156, n_23157, n_23158, n_23159,
       n_23160;
  wire n_23165, n_23166, n_23167, n_23168, n_23169, n_23170, n_23171,
       n_23172;
  wire n_23173, n_23174, n_23175, n_23176, n_23181, n_23182, n_23183,
       n_23184;
  wire n_23185, n_23186, n_23187, n_23188, n_23189, n_23190, n_23191,
       n_23192;
  wire n_23193, n_23194, n_23195, n_23196, n_23197, n_23198, n_23199,
       n_23200;
  wire n_23201, n_23202, n_23203, n_23204, n_23205, n_23206, n_23207,
       n_23208;
  wire n_23209, n_23210, n_23211, n_23212, n_23213, n_23214, n_23215,
       n_23216;
  wire n_23217, n_23218, n_23219, n_23220, n_23225, n_23226, n_23227,
       n_23228;
  wire n_23229, n_23230, n_23231, n_23232, n_23233, n_23234, n_23235,
       n_23236;
  wire n_23237, n_23238, n_23239, n_23240, n_23241, n_23242, n_23243,
       n_23244;
  wire n_23245, n_23246, n_23247, n_23248, n_23249, n_23250, n_23251,
       n_23252;
  wire n_23253, n_23254, n_23255, n_23256, n_23257, n_23258, n_23259,
       n_23260;
  wire n_23261, n_23262, n_23263, n_23264, n_23265, n_23266, n_23267,
       n_23268;
  wire n_23269, n_23270, n_23271, n_23272, n_23273, n_23278, n_23279,
       n_23280;
  wire n_23281, n_23282, n_23283, n_23284, n_23285, n_23286, n_23287,
       n_23288;
  wire n_23289, n_23290, n_23291, n_23292, n_23293, n_23294, n_23295,
       n_23296;
  wire n_23301, n_23302, n_23303, n_23304, n_23305, n_23306, n_23307,
       n_23308;
  wire n_23309, n_23310, n_23311, n_23312, n_23313, n_23314, n_23315,
       n_23316;
  wire n_23317, n_23318, n_23319, n_23320, n_23321, n_23322, n_23323,
       n_23324;
  wire n_23325, n_23326, n_23327, n_23328, n_23329, n_23330, n_23331,
       n_23336;
  wire n_23337, n_23338, n_23339, n_23340, n_23341, n_23342, n_23343,
       n_23344;
  wire n_23345, n_23346, n_23347, n_23348, n_23349, n_23350, n_23351,
       n_23352;
  wire n_23353, n_23354, n_23355, n_23356, n_23357, n_23358, n_23363,
       n_23364;
  wire n_23365, n_23366, n_23367, n_23368, n_23369, n_23370, n_23371,
       n_23372;
  wire n_23373, n_23374, n_23375, n_23376, n_23377, n_23378, n_23379,
       n_23380;
  wire n_23381, n_23382, n_23383, n_23384, n_23385, n_23386, n_23387,
       n_23388;
  wire n_23389, n_23390, n_23391, n_23392, n_23393, n_23394, n_23395,
       n_23396;
  wire n_23397, n_23398, n_23399, n_23400, n_23401, n_23402, n_23403,
       n_23404;
  wire n_23405, n_23406, n_23407, n_23408, n_23409, n_23410, n_23411,
       n_23412;
  wire n_23413, n_23414, n_23415, n_23416, n_23417, n_23418, n_23419,
       n_23420;
  wire n_23421, n_23422, n_23423, n_23424, n_23425, n_23426, n_23427,
       n_23428;
  wire n_23429, n_23430, n_23431, n_23432, n_23437, n_23438, n_23439,
       n_23440;
  wire n_23441, n_23442, n_23443, n_23444, n_23445, n_23446, n_23447,
       n_23448;
  wire n_23449, n_23450, n_23451, n_23452, n_23453, n_23454, n_23455,
       n_23456;
  wire n_23457, n_23458, n_23459, n_23460, n_23461, n_23462, n_23463,
       n_23464;
  wire n_23465, n_23466, n_23467, n_23468, n_23469, n_23470, n_23471,
       n_23472;
  wire n_23473, n_23478, n_23479, n_23480, n_23481, n_23482, n_23483,
       n_23484;
  wire n_23485, n_23486, n_23487, n_23488, n_23489, n_23490, n_23491,
       n_23492;
  wire n_23493, n_23494, n_23495, n_23496, n_23497, n_23498, n_23499,
       n_23500;
  wire n_23501, n_23502, n_23503, n_23504, n_23505, n_23506, n_23507,
       n_23508;
  wire n_23509, n_23510, n_23511, n_23512, n_23513, n_23514, n_23515,
       n_23516;
  wire n_23517, n_23518, n_23519, n_23520, n_23521, n_23522, n_23523,
       n_23524;
  wire n_23525, n_23526, n_23527, n_23528, n_23529, n_23530, n_23531,
       n_23532;
  wire n_23533, n_23534, n_23535, n_23536, n_23537, n_23538, n_23539,
       n_23540;
  wire n_23541, n_23542, n_23543, n_23544, n_23545, n_23546, n_23547,
       n_23548;
  wire n_23549, n_23550, n_23551, n_23552, n_23553, n_23554, n_23555,
       n_23556;
  wire n_23557, n_23558, n_23559, n_23560, n_23561, n_23562, n_23563,
       n_23564;
  wire n_23565, n_23566, n_23567, n_23568, n_23569, n_23570;
  and g1 (n257, \a[0] , \b[0] );
  not g2 (n_4, n257);
  and g3 (n258, \a[2] , n_4);
  not g4 (n_5, \a[2] );
  and g5 (n259, n_5, n_4);
  not g6 (n_6, n258);
  not g7 (n_7, n259);
  and g8 (\f[0] , n_6, n_7);
  not g9 (n_8, \a[0] );
  and g10 (n261, n_8, \a[1] );
  and g11 (n262, \b[0] , n261);
  not g12 (n_10, \a[1] );
  and g13 (n263, n_10, \a[2] );
  and g14 (n264, \a[1] , n_5);
  not g15 (n_11, n263);
  not g16 (n_12, n264);
  and g17 (n265, n_11, n_12);
  and g18 (n266, \a[0] , n265);
  and g19 (n267, \b[1] , n266);
  not g20 (n_14, n262);
  not g21 (n_15, n267);
  and g22 (n268, n_14, n_15);
  not g23 (n_16, n265);
  and g24 (n269, \a[0] , n_16);
  not g25 (n_17, \b[1] );
  and g26 (n270, \b[0] , n_17);
  not g27 (n_18, \b[0] );
  and g28 (n271, n_18, \b[1] );
  not g29 (n_19, n270);
  not g30 (n_20, n271);
  and g31 (n272, n_19, n_20);
  not g32 (n_21, n272);
  and g33 (n273, n269, n_21);
  not g34 (n_22, n273);
  and g35 (n274, n268, n_22);
  not g36 (n_23, n274);
  and g37 (n275, \a[2] , n_23);
  not g38 (n_24, n275);
  and g39 (n276, \a[2] , n_24);
  and g40 (n277, n_23, n_24);
  not g41 (n_25, n276);
  not g42 (n_26, n277);
  and g43 (n278, n_25, n_26);
  not g44 (n_27, n278);
  and g45 (n279, n258, n_27);
  and g46 (n280, n_6, n278);
  not g47 (n_28, n279);
  not g48 (n_29, n280);
  and g49 (\f[1] , n_28, n_29);
  and g50 (n282, \b[2] , n266);
  and g51 (n283, n_8, n_16);
  and g52 (n284, n_10, n283);
  and g53 (n285, \b[0] , n284);
  and g54 (n286, \b[1] , n261);
  not g60 (n_34, \b[2] );
  and g61 (n289, \b[0] , n_34);
  and g62 (n290, \b[1] , n289);
  and g63 (n291, \b[1] , n_34);
  and g64 (n292, n_17, \b[2] );
  not g65 (n_35, n291);
  not g66 (n_36, n292);
  and g67 (n293, n_35, n_36);
  and g68 (n294, \b[0] , \b[1] );
  not g69 (n_37, n294);
  and g70 (n295, n293, n_37);
  not g71 (n_38, n290);
  not g72 (n_39, n295);
  and g73 (n296, n_38, n_39);
  and g74 (n297, n269, n296);
  not g77 (n_41, n298);
  and g78 (n299, \a[2] , n_41);
  not g79 (n_42, n299);
  and g80 (n300, \a[2] , n_42);
  and g81 (n301, n_41, n_42);
  not g82 (n_43, n300);
  not g83 (n_44, n301);
  and g84 (n302, n_43, n_44);
  not g85 (n_45, n302);
  and g86 (n303, n279, n_45);
  and g87 (n304, n_28, n302);
  not g88 (n_46, n303);
  not g89 (n_47, n304);
  and g90 (\f[2] , n_46, n_47);
  and g91 (n306, \b[3] , n266);
  and g92 (n307, \b[1] , n284);
  and g93 (n308, \b[2] , n261);
  and g99 (n311, \b[1] , \b[2] );
  not g100 (n_52, n311);
  and g101 (n312, n_38, n_52);
  not g102 (n_53, \b[3] );
  and g103 (n313, n_34, n_53);
  and g104 (n314, \b[2] , \b[3] );
  not g105 (n_54, n313);
  not g106 (n_55, n314);
  and g107 (n315, n_54, n_55);
  not g108 (n_56, n312);
  and g109 (n316, n_56, n315);
  not g110 (n_57, n315);
  and g111 (n317, n312, n_57);
  not g112 (n_58, n316);
  not g113 (n_59, n317);
  and g114 (n318, n_58, n_59);
  and g115 (n319, n269, n318);
  not g118 (n_61, n320);
  and g119 (n321, \a[2] , n_61);
  not g120 (n_62, n321);
  and g121 (n322, \a[2] , n_62);
  and g122 (n323, n_61, n_62);
  not g123 (n_63, n322);
  not g124 (n_64, n323);
  and g125 (n324, n_63, n_64);
  not g126 (n_66, \a[3] );
  and g127 (n325, \a[2] , n_66);
  and g128 (n326, n_5, \a[3] );
  not g129 (n_67, n325);
  not g130 (n_68, n326);
  and g131 (n327, n_67, n_68);
  not g132 (n_69, n327);
  and g133 (n328, \b[0] , n_69);
  not g134 (n_70, n324);
  and g135 (n329, n_70, n328);
  not g136 (n_71, n328);
  and g137 (n330, n324, n_71);
  not g138 (n_72, n329);
  not g139 (n_73, n330);
  and g140 (n331, n_72, n_73);
  and g141 (n332, n303, n331);
  not g142 (n_74, n331);
  and g143 (n333, n_46, n_74);
  not g144 (n_75, n332);
  not g145 (n_76, n333);
  and g146 (\f[3] , n_75, n_76);
  and g147 (n335, \b[4] , n266);
  and g148 (n336, \b[2] , n284);
  and g149 (n337, \b[3] , n261);
  and g155 (n340, n_55, n_58);
  not g156 (n_81, \b[4] );
  and g157 (n341, n_53, n_81);
  and g158 (n342, \b[3] , \b[4] );
  not g159 (n_82, n341);
  not g160 (n_83, n342);
  and g161 (n343, n_82, n_83);
  not g162 (n_84, n340);
  and g163 (n344, n_84, n343);
  not g164 (n_85, n343);
  and g165 (n345, n340, n_85);
  not g166 (n_86, n344);
  not g167 (n_87, n345);
  and g168 (n346, n_86, n_87);
  and g169 (n347, n269, n346);
  not g172 (n_89, n348);
  and g173 (n349, \a[2] , n_89);
  not g174 (n_90, n349);
  and g175 (n350, \a[2] , n_90);
  and g176 (n351, n_89, n_90);
  not g177 (n_91, n350);
  not g178 (n_92, n351);
  and g179 (n352, n_91, n_92);
  and g180 (n353, \a[5] , n_71);
  and g181 (n354, n_66, \a[4] );
  not g182 (n_95, \a[4] );
  and g183 (n355, \a[3] , n_95);
  not g184 (n_96, n354);
  not g185 (n_97, n355);
  and g186 (n356, n_96, n_97);
  not g187 (n_98, n356);
  and g188 (n357, n327, n_98);
  and g189 (n358, \b[0] , n357);
  and g190 (n359, n_95, \a[5] );
  not g191 (n_99, \a[5] );
  and g192 (n360, \a[4] , n_99);
  not g193 (n_100, n359);
  not g194 (n_101, n360);
  and g195 (n361, n_100, n_101);
  and g196 (n362, n_69, n361);
  and g197 (n363, \b[1] , n362);
  not g198 (n_102, n358);
  not g199 (n_103, n363);
  and g200 (n364, n_102, n_103);
  not g201 (n_104, n361);
  and g202 (n365, n_69, n_104);
  and g203 (n366, n_21, n365);
  not g204 (n_105, n366);
  and g205 (n367, n364, n_105);
  not g206 (n_106, n367);
  and g207 (n368, \a[5] , n_106);
  not g208 (n_107, n368);
  and g209 (n369, \a[5] , n_107);
  and g210 (n370, n_106, n_107);
  not g211 (n_108, n369);
  not g212 (n_109, n370);
  and g213 (n371, n_108, n_109);
  not g214 (n_110, n371);
  and g215 (n372, n353, n_110);
  not g216 (n_111, n353);
  and g217 (n373, n_111, n371);
  not g218 (n_112, n372);
  not g219 (n_113, n373);
  and g220 (n374, n_112, n_113);
  not g221 (n_114, n352);
  and g222 (n375, n_114, n374);
  not g223 (n_115, n375);
  and g224 (n376, n374, n_115);
  and g225 (n377, n_114, n_115);
  not g226 (n_116, n376);
  not g227 (n_117, n377);
  and g228 (n378, n_116, n_117);
  and g229 (n379, n_72, n_75);
  not g230 (n_118, n378);
  not g231 (n_119, n379);
  and g232 (n380, n_118, n_119);
  and g233 (n381, n378, n379);
  not g234 (n_120, n380);
  not g235 (n_121, n381);
  and g236 (\f[4] , n_120, n_121);
  and g237 (n383, \b[5] , n266);
  and g238 (n384, \b[3] , n284);
  and g239 (n385, \b[4] , n261);
  and g245 (n388, n_83, n_86);
  not g246 (n_126, \b[5] );
  and g247 (n389, n_81, n_126);
  and g248 (n390, \b[4] , \b[5] );
  not g249 (n_127, n389);
  not g250 (n_128, n390);
  and g251 (n391, n_127, n_128);
  not g252 (n_129, n388);
  and g253 (n392, n_129, n391);
  not g254 (n_130, n391);
  and g255 (n393, n388, n_130);
  not g256 (n_131, n392);
  not g257 (n_132, n393);
  and g258 (n394, n_131, n_132);
  and g259 (n395, n269, n394);
  not g262 (n_134, n396);
  and g263 (n397, \a[2] , n_134);
  not g264 (n_135, n397);
  and g265 (n398, \a[2] , n_135);
  and g266 (n399, n_134, n_135);
  not g267 (n_136, n398);
  not g268 (n_137, n399);
  and g269 (n400, n_136, n_137);
  and g270 (n401, \b[2] , n362);
  and g271 (n402, n327, n_104);
  and g272 (n403, n356, n402);
  and g273 (n404, \b[0] , n403);
  and g274 (n405, \b[1] , n357);
  not g275 (n_138, n404);
  not g276 (n_139, n405);
  and g277 (n406, n_138, n_139);
  not g278 (n_140, n401);
  and g279 (n407, n_140, n406);
  not g280 (n_141, n365);
  and g281 (n408, n_141, n407);
  not g282 (n_142, n296);
  and g283 (n409, n_142, n407);
  not g284 (n_143, n408);
  not g285 (n_144, n409);
  and g286 (n410, n_143, n_144);
  not g287 (n_145, n410);
  and g288 (n411, \a[5] , n_145);
  and g289 (n412, n_99, n410);
  not g290 (n_146, n411);
  not g291 (n_147, n412);
  and g292 (n413, n_146, n_147);
  not g293 (n_148, n413);
  and g294 (n414, n372, n_148);
  and g295 (n415, n_112, n413);
  not g296 (n_149, n414);
  not g297 (n_150, n415);
  and g298 (n416, n_149, n_150);
  not g299 (n_151, n400);
  and g300 (n417, n_151, n416);
  not g301 (n_152, n417);
  and g302 (n418, n416, n_152);
  and g303 (n419, n_151, n_152);
  not g304 (n_153, n418);
  not g305 (n_154, n419);
  and g306 (n420, n_153, n_154);
  and g307 (n421, n_115, n_120);
  not g308 (n_155, n420);
  not g309 (n_156, n421);
  and g310 (n422, n_155, n_156);
  and g311 (n423, n420, n421);
  not g312 (n_157, n422);
  not g313 (n_158, n423);
  and g314 (\f[5] , n_157, n_158);
  and g315 (n425, n_152, n_157);
  not g316 (n_160, \a[6] );
  and g317 (n426, \a[5] , n_160);
  and g318 (n427, n_99, \a[6] );
  not g319 (n_161, n426);
  not g320 (n_162, n427);
  and g321 (n428, n_161, n_162);
  not g322 (n_163, n428);
  and g323 (n429, \b[0] , n_163);
  and g324 (n430, n414, n429);
  not g325 (n_164, n430);
  and g326 (n431, n414, n_164);
  and g327 (n432, n429, n_164);
  not g328 (n_165, n431);
  not g329 (n_166, n432);
  and g330 (n433, n_165, n_166);
  and g331 (n434, \b[3] , n362);
  and g332 (n435, \b[1] , n403);
  and g333 (n436, \b[2] , n357);
  and g339 (n439, n318, n365);
  not g342 (n_171, n440);
  and g343 (n441, \a[5] , n_171);
  not g344 (n_172, n441);
  and g345 (n442, \a[5] , n_172);
  and g346 (n443, n_171, n_172);
  not g347 (n_173, n442);
  not g348 (n_174, n443);
  and g349 (n444, n_173, n_174);
  not g350 (n_175, n433);
  and g351 (n445, n_175, n444);
  not g352 (n_176, n444);
  and g353 (n446, n433, n_176);
  not g354 (n_177, n445);
  not g355 (n_178, n446);
  and g356 (n447, n_177, n_178);
  and g357 (n448, \b[6] , n266);
  and g358 (n449, \b[4] , n284);
  and g359 (n450, \b[5] , n261);
  and g365 (n453, n_128, n_131);
  not g366 (n_183, \b[6] );
  and g367 (n454, n_126, n_183);
  and g368 (n455, \b[5] , \b[6] );
  not g369 (n_184, n454);
  not g370 (n_185, n455);
  and g371 (n456, n_184, n_185);
  not g372 (n_186, n453);
  and g373 (n457, n_186, n456);
  not g374 (n_187, n456);
  and g375 (n458, n453, n_187);
  not g376 (n_188, n457);
  not g377 (n_189, n458);
  and g378 (n459, n_188, n_189);
  and g379 (n460, n269, n459);
  not g382 (n_191, n461);
  and g383 (n462, \a[2] , n_191);
  not g384 (n_192, n462);
  and g385 (n463, \a[2] , n_192);
  and g386 (n464, n_191, n_192);
  not g387 (n_193, n463);
  not g388 (n_194, n464);
  and g389 (n465, n_193, n_194);
  not g390 (n_195, n447);
  not g391 (n_196, n465);
  and g392 (n466, n_195, n_196);
  and g393 (n467, n447, n465);
  not g394 (n_197, n466);
  not g395 (n_198, n467);
  and g396 (n468, n_197, n_198);
  not g397 (n_199, n425);
  and g398 (n469, n_199, n468);
  not g399 (n_200, n468);
  and g400 (n470, n425, n_200);
  not g401 (n_201, n469);
  not g402 (n_202, n470);
  and g403 (\f[6] , n_201, n_202);
  and g404 (n472, n_197, n_201);
  and g405 (n473, \b[7] , n266);
  and g406 (n474, \b[5] , n284);
  and g407 (n475, \b[6] , n261);
  and g413 (n478, n_185, n_188);
  not g414 (n_207, \b[7] );
  and g415 (n479, n_183, n_207);
  and g416 (n480, \b[6] , \b[7] );
  not g417 (n_208, n479);
  not g418 (n_209, n480);
  and g419 (n481, n_208, n_209);
  not g420 (n_210, n478);
  and g421 (n482, n_210, n481);
  not g422 (n_211, n481);
  and g423 (n483, n478, n_211);
  not g424 (n_212, n482);
  not g425 (n_213, n483);
  and g426 (n484, n_212, n_213);
  and g427 (n485, n269, n484);
  not g430 (n_215, n486);
  and g431 (n487, \a[2] , n_215);
  not g432 (n_216, n487);
  and g433 (n488, \a[2] , n_216);
  and g434 (n489, n_215, n_216);
  not g435 (n_217, n488);
  not g436 (n_218, n489);
  and g437 (n490, n_217, n_218);
  and g438 (n491, \b[4] , n362);
  and g439 (n492, \b[2] , n403);
  and g440 (n493, \b[3] , n357);
  and g446 (n496, n346, n365);
  not g449 (n_223, n497);
  and g450 (n498, \a[5] , n_223);
  not g451 (n_224, n498);
  and g452 (n499, \a[5] , n_224);
  and g453 (n500, n_223, n_224);
  not g454 (n_225, n499);
  not g455 (n_226, n500);
  and g456 (n501, n_225, n_226);
  not g457 (n_228, n429);
  and g458 (n502, \a[8] , n_228);
  and g459 (n503, n_160, \a[7] );
  not g460 (n_230, \a[7] );
  and g461 (n504, \a[6] , n_230);
  not g462 (n_231, n503);
  not g463 (n_232, n504);
  and g464 (n505, n_231, n_232);
  not g465 (n_233, n505);
  and g466 (n506, n428, n_233);
  and g467 (n507, \b[0] , n506);
  and g468 (n508, n_230, \a[8] );
  not g469 (n_234, \a[8] );
  and g470 (n509, \a[7] , n_234);
  not g471 (n_235, n508);
  not g472 (n_236, n509);
  and g473 (n510, n_235, n_236);
  and g474 (n511, n_163, n510);
  and g475 (n512, \b[1] , n511);
  not g476 (n_237, n507);
  not g477 (n_238, n512);
  and g478 (n513, n_237, n_238);
  not g479 (n_239, n510);
  and g480 (n514, n_163, n_239);
  and g481 (n515, n_21, n514);
  not g482 (n_240, n515);
  and g483 (n516, n513, n_240);
  not g484 (n_241, n516);
  and g485 (n517, \a[8] , n_241);
  not g486 (n_242, n517);
  and g487 (n518, \a[8] , n_242);
  and g488 (n519, n_241, n_242);
  not g489 (n_243, n518);
  not g490 (n_244, n519);
  and g491 (n520, n_243, n_244);
  not g492 (n_245, n520);
  and g493 (n521, n502, n_245);
  not g494 (n_246, n502);
  and g495 (n522, n_246, n520);
  not g496 (n_247, n521);
  not g497 (n_248, n522);
  and g498 (n523, n_247, n_248);
  not g499 (n_249, n501);
  and g500 (n524, n_249, n523);
  not g501 (n_250, n524);
  and g502 (n525, n523, n_250);
  and g503 (n526, n_249, n_250);
  not g504 (n_251, n525);
  not g505 (n_252, n526);
  and g506 (n527, n_251, n_252);
  and g507 (n528, n_175, n_176);
  not g508 (n_253, n528);
  and g509 (n529, n_164, n_253);
  not g510 (n_254, n527);
  not g511 (n_255, n529);
  and g512 (n530, n_254, n_255);
  and g513 (n531, n527, n529);
  not g514 (n_256, n530);
  not g515 (n_257, n531);
  and g516 (n532, n_256, n_257);
  not g517 (n_258, n490);
  and g518 (n533, n_258, n532);
  not g519 (n_259, n532);
  and g520 (n534, n490, n_259);
  not g521 (n_260, n533);
  not g522 (n_261, n534);
  and g523 (n535, n_260, n_261);
  not g524 (n_262, n472);
  and g525 (n536, n_262, n535);
  not g526 (n_263, n535);
  and g527 (n537, n472, n_263);
  not g528 (n_264, n536);
  not g529 (n_265, n537);
  and g530 (\f[7] , n_264, n_265);
  and g531 (n539, \b[2] , n511);
  and g532 (n540, n428, n_239);
  and g533 (n541, n505, n540);
  and g534 (n542, \b[0] , n541);
  and g535 (n543, \b[1] , n506);
  and g541 (n546, n296, n514);
  not g544 (n_270, n547);
  and g545 (n548, \a[8] , n_270);
  not g546 (n_271, n548);
  and g547 (n549, \a[8] , n_271);
  and g548 (n550, n_270, n_271);
  not g549 (n_272, n549);
  not g550 (n_273, n550);
  and g551 (n551, n_272, n_273);
  and g552 (n552, n_247, n551);
  not g553 (n_274, n551);
  and g554 (n553, n521, n_274);
  not g555 (n_275, n552);
  not g556 (n_276, n553);
  and g557 (n554, n_275, n_276);
  and g558 (n555, \b[5] , n362);
  and g559 (n556, \b[3] , n403);
  and g560 (n557, \b[4] , n357);
  and g566 (n560, n365, n394);
  not g569 (n_281, n561);
  and g570 (n562, \a[5] , n_281);
  not g571 (n_282, n562);
  and g572 (n563, \a[5] , n_282);
  and g573 (n564, n_281, n_282);
  not g574 (n_283, n563);
  not g575 (n_284, n564);
  and g576 (n565, n_283, n_284);
  not g577 (n_285, n565);
  and g578 (n566, n554, n_285);
  not g579 (n_286, n566);
  and g580 (n567, n554, n_286);
  and g581 (n568, n_285, n_286);
  not g582 (n_287, n567);
  not g583 (n_288, n568);
  and g584 (n569, n_287, n_288);
  and g585 (n570, n_250, n_256);
  and g586 (n571, n569, n570);
  not g587 (n_289, n569);
  not g588 (n_290, n570);
  and g589 (n572, n_289, n_290);
  not g590 (n_291, n571);
  not g591 (n_292, n572);
  and g592 (n573, n_291, n_292);
  and g593 (n574, \b[8] , n266);
  and g594 (n575, \b[6] , n284);
  and g595 (n576, \b[7] , n261);
  and g601 (n579, n_209, n_212);
  not g602 (n_297, \b[8] );
  and g603 (n580, n_207, n_297);
  and g604 (n581, \b[7] , \b[8] );
  not g605 (n_298, n580);
  not g606 (n_299, n581);
  and g607 (n582, n_298, n_299);
  not g608 (n_300, n579);
  and g609 (n583, n_300, n582);
  not g610 (n_301, n582);
  and g611 (n584, n579, n_301);
  not g612 (n_302, n583);
  not g613 (n_303, n584);
  and g614 (n585, n_302, n_303);
  and g615 (n586, n269, n585);
  not g618 (n_305, n587);
  and g619 (n588, \a[2] , n_305);
  not g620 (n_306, n588);
  and g621 (n589, \a[2] , n_306);
  and g622 (n590, n_305, n_306);
  not g623 (n_307, n589);
  not g624 (n_308, n590);
  and g625 (n591, n_307, n_308);
  not g626 (n_309, n591);
  and g627 (n592, n573, n_309);
  not g628 (n_310, n592);
  and g629 (n593, n573, n_310);
  and g630 (n594, n_309, n_310);
  not g631 (n_311, n593);
  not g632 (n_312, n594);
  and g633 (n595, n_311, n_312);
  and g634 (n596, n_260, n_264);
  not g635 (n_313, n595);
  not g636 (n_314, n596);
  and g637 (n597, n_313, n_314);
  and g638 (n598, n595, n596);
  not g639 (n_315, n597);
  not g640 (n_316, n598);
  and g641 (\f[8] , n_315, n_316);
  and g642 (n600, \b[6] , n362);
  and g643 (n601, \b[4] , n403);
  and g644 (n602, \b[5] , n357);
  and g650 (n605, n365, n459);
  not g653 (n_321, n606);
  and g654 (n607, \a[5] , n_321);
  not g655 (n_322, n607);
  and g656 (n608, \a[5] , n_322);
  and g657 (n609, n_321, n_322);
  not g658 (n_323, n608);
  not g659 (n_324, n609);
  and g660 (n610, n_323, n_324);
  not g661 (n_326, \a[9] );
  and g662 (n611, \a[8] , n_326);
  and g663 (n612, n_234, \a[9] );
  not g664 (n_327, n611);
  not g665 (n_328, n612);
  and g666 (n613, n_327, n_328);
  not g667 (n_329, n613);
  and g668 (n614, \b[0] , n_329);
  and g669 (n615, n_276, n614);
  not g670 (n_330, n614);
  and g671 (n616, n553, n_330);
  not g672 (n_331, n615);
  not g673 (n_332, n616);
  and g674 (n617, n_331, n_332);
  and g675 (n618, \b[3] , n511);
  and g676 (n619, \b[1] , n541);
  and g677 (n620, \b[2] , n506);
  and g683 (n623, n318, n514);
  not g686 (n_337, n624);
  and g687 (n625, \a[8] , n_337);
  not g688 (n_338, n625);
  and g689 (n626, \a[8] , n_338);
  and g690 (n627, n_337, n_338);
  not g691 (n_339, n626);
  not g692 (n_340, n627);
  and g693 (n628, n_339, n_340);
  not g694 (n_341, n617);
  not g695 (n_342, n628);
  and g696 (n629, n_341, n_342);
  and g697 (n630, n617, n628);
  not g698 (n_343, n629);
  not g699 (n_344, n630);
  and g700 (n631, n_343, n_344);
  not g701 (n_345, n610);
  and g702 (n632, n_345, n631);
  not g703 (n_346, n632);
  and g704 (n633, n631, n_346);
  and g705 (n634, n_345, n_346);
  not g706 (n_347, n633);
  not g707 (n_348, n634);
  and g708 (n635, n_347, n_348);
  and g709 (n636, n_286, n_292);
  and g710 (n637, n635, n636);
  not g711 (n_349, n635);
  not g712 (n_350, n636);
  and g713 (n638, n_349, n_350);
  not g714 (n_351, n637);
  not g715 (n_352, n638);
  and g716 (n639, n_351, n_352);
  and g717 (n640, \b[9] , n266);
  and g718 (n641, \b[7] , n284);
  and g719 (n642, \b[8] , n261);
  and g725 (n645, n_299, n_302);
  not g726 (n_357, \b[9] );
  and g727 (n646, n_297, n_357);
  and g728 (n647, \b[8] , \b[9] );
  not g729 (n_358, n646);
  not g730 (n_359, n647);
  and g731 (n648, n_358, n_359);
  not g732 (n_360, n645);
  and g733 (n649, n_360, n648);
  not g734 (n_361, n648);
  and g735 (n650, n645, n_361);
  not g736 (n_362, n649);
  not g737 (n_363, n650);
  and g738 (n651, n_362, n_363);
  and g739 (n652, n269, n651);
  not g742 (n_365, n653);
  and g743 (n654, \a[2] , n_365);
  not g744 (n_366, n654);
  and g745 (n655, \a[2] , n_366);
  and g746 (n656, n_365, n_366);
  not g747 (n_367, n655);
  not g748 (n_368, n656);
  and g749 (n657, n_367, n_368);
  not g750 (n_369, n657);
  and g751 (n658, n639, n_369);
  not g752 (n_370, n658);
  and g753 (n659, n639, n_370);
  and g754 (n660, n_369, n_370);
  not g755 (n_371, n659);
  not g756 (n_372, n660);
  and g757 (n661, n_371, n_372);
  and g758 (n662, n_310, n_315);
  not g759 (n_373, n661);
  not g760 (n_374, n662);
  and g761 (n663, n_373, n_374);
  and g762 (n664, n661, n662);
  not g763 (n_375, n663);
  not g764 (n_376, n664);
  and g765 (\f[9] , n_375, n_376);
  and g766 (n666, n_370, n_375);
  and g767 (n667, \b[7] , n362);
  and g768 (n668, \b[5] , n403);
  and g769 (n669, \b[6] , n357);
  and g775 (n672, n365, n484);
  not g778 (n_381, n673);
  and g779 (n674, \a[5] , n_381);
  not g780 (n_382, n674);
  and g781 (n675, \a[5] , n_382);
  and g782 (n676, n_381, n_382);
  not g783 (n_383, n675);
  not g784 (n_384, n676);
  and g785 (n677, n_383, n_384);
  and g786 (n678, n553, n614);
  not g787 (n_385, n678);
  and g788 (n679, n_343, n_385);
  and g789 (n680, \b[4] , n511);
  and g790 (n681, \b[2] , n541);
  and g791 (n682, \b[3] , n506);
  and g797 (n685, n346, n514);
  not g800 (n_390, n686);
  and g801 (n687, \a[8] , n_390);
  not g802 (n_391, n687);
  and g803 (n688, \a[8] , n_391);
  and g804 (n689, n_390, n_391);
  not g805 (n_392, n688);
  not g806 (n_393, n689);
  and g807 (n690, n_392, n_393);
  and g808 (n691, \a[11] , n_330);
  and g809 (n692, n_326, \a[10] );
  not g810 (n_396, \a[10] );
  and g811 (n693, \a[9] , n_396);
  not g812 (n_397, n692);
  not g813 (n_398, n693);
  and g814 (n694, n_397, n_398);
  not g815 (n_399, n694);
  and g816 (n695, n613, n_399);
  and g817 (n696, \b[0] , n695);
  and g818 (n697, n_396, \a[11] );
  not g819 (n_400, \a[11] );
  and g820 (n698, \a[10] , n_400);
  not g821 (n_401, n697);
  not g822 (n_402, n698);
  and g823 (n699, n_401, n_402);
  and g824 (n700, n_329, n699);
  and g825 (n701, \b[1] , n700);
  not g826 (n_403, n696);
  not g827 (n_404, n701);
  and g828 (n702, n_403, n_404);
  not g829 (n_405, n699);
  and g830 (n703, n_329, n_405);
  and g831 (n704, n_21, n703);
  not g832 (n_406, n704);
  and g833 (n705, n702, n_406);
  not g834 (n_407, n705);
  and g835 (n706, \a[11] , n_407);
  not g836 (n_408, n706);
  and g837 (n707, \a[11] , n_408);
  and g838 (n708, n_407, n_408);
  not g839 (n_409, n707);
  not g840 (n_410, n708);
  and g841 (n709, n_409, n_410);
  not g842 (n_411, n709);
  and g843 (n710, n691, n_411);
  not g844 (n_412, n691);
  and g845 (n711, n_412, n709);
  not g846 (n_413, n710);
  not g847 (n_414, n711);
  and g848 (n712, n_413, n_414);
  not g849 (n_415, n712);
  and g850 (n713, n690, n_415);
  not g851 (n_416, n690);
  and g852 (n714, n_416, n712);
  not g853 (n_417, n713);
  not g854 (n_418, n714);
  and g855 (n715, n_417, n_418);
  not g856 (n_419, n679);
  and g857 (n716, n_419, n715);
  not g858 (n_420, n715);
  and g859 (n717, n679, n_420);
  not g860 (n_421, n716);
  not g861 (n_422, n717);
  and g862 (n718, n_421, n_422);
  not g863 (n_423, n677);
  and g864 (n719, n_423, n718);
  not g865 (n_424, n719);
  and g866 (n720, n718, n_424);
  and g867 (n721, n_423, n_424);
  not g868 (n_425, n720);
  not g869 (n_426, n721);
  and g870 (n722, n_425, n_426);
  and g871 (n723, n_346, n_352);
  and g872 (n724, n722, n723);
  not g873 (n_427, n722);
  not g874 (n_428, n723);
  and g875 (n725, n_427, n_428);
  not g876 (n_429, n724);
  not g877 (n_430, n725);
  and g878 (n726, n_429, n_430);
  and g879 (n727, \b[10] , n266);
  and g880 (n728, \b[8] , n284);
  and g881 (n729, \b[9] , n261);
  and g887 (n732, n_359, n_362);
  not g888 (n_435, \b[10] );
  and g889 (n733, n_357, n_435);
  and g890 (n734, \b[9] , \b[10] );
  not g891 (n_436, n733);
  not g892 (n_437, n734);
  and g893 (n735, n_436, n_437);
  not g894 (n_438, n732);
  and g895 (n736, n_438, n735);
  not g896 (n_439, n735);
  and g897 (n737, n732, n_439);
  not g898 (n_440, n736);
  not g899 (n_441, n737);
  and g900 (n738, n_440, n_441);
  and g901 (n739, n269, n738);
  not g904 (n_443, n740);
  and g905 (n741, \a[2] , n_443);
  not g906 (n_444, n741);
  and g907 (n742, \a[2] , n_444);
  and g908 (n743, n_443, n_444);
  not g909 (n_445, n742);
  not g910 (n_446, n743);
  and g911 (n744, n_445, n_446);
  not g912 (n_447, n726);
  and g913 (n745, n_447, n744);
  not g914 (n_448, n744);
  and g915 (n746, n726, n_448);
  not g916 (n_449, n745);
  not g917 (n_450, n746);
  and g918 (n747, n_449, n_450);
  not g919 (n_451, n666);
  and g920 (n748, n_451, n747);
  not g921 (n_452, n747);
  and g922 (n749, n666, n_452);
  not g923 (n_453, n748);
  not g924 (n_454, n749);
  and g925 (\f[10] , n_453, n_454);
  and g926 (n751, n_450, n_453);
  and g927 (n752, n_424, n_430);
  and g928 (n753, \b[8] , n362);
  and g929 (n754, \b[6] , n403);
  and g930 (n755, \b[7] , n357);
  and g936 (n758, n365, n585);
  not g939 (n_459, n759);
  and g940 (n760, \a[5] , n_459);
  not g941 (n_460, n760);
  and g942 (n761, \a[5] , n_460);
  and g943 (n762, n_459, n_460);
  not g944 (n_461, n761);
  not g945 (n_462, n762);
  and g946 (n763, n_461, n_462);
  and g947 (n764, n_418, n_421);
  and g948 (n765, \b[2] , n700);
  and g949 (n766, n613, n_405);
  and g950 (n767, n694, n766);
  and g951 (n768, \b[0] , n767);
  and g952 (n769, \b[1] , n695);
  and g958 (n772, n296, n703);
  not g961 (n_467, n773);
  and g962 (n774, \a[11] , n_467);
  not g963 (n_468, n774);
  and g964 (n775, \a[11] , n_468);
  and g965 (n776, n_467, n_468);
  not g966 (n_469, n775);
  not g967 (n_470, n776);
  and g968 (n777, n_469, n_470);
  and g969 (n778, n_413, n777);
  not g970 (n_471, n777);
  and g971 (n779, n710, n_471);
  not g972 (n_472, n778);
  not g973 (n_473, n779);
  and g974 (n780, n_472, n_473);
  and g975 (n781, \b[5] , n511);
  and g976 (n782, \b[3] , n541);
  and g977 (n783, \b[4] , n506);
  and g983 (n786, n394, n514);
  not g986 (n_478, n787);
  and g987 (n788, \a[8] , n_478);
  not g988 (n_479, n788);
  and g989 (n789, \a[8] , n_479);
  and g990 (n790, n_478, n_479);
  not g991 (n_480, n789);
  not g992 (n_481, n790);
  and g993 (n791, n_480, n_481);
  not g994 (n_482, n791);
  and g995 (n792, n780, n_482);
  not g996 (n_483, n792);
  and g997 (n793, n780, n_483);
  and g998 (n794, n_482, n_483);
  not g999 (n_484, n793);
  not g1000 (n_485, n794);
  and g1001 (n795, n_484, n_485);
  not g1002 (n_486, n764);
  not g1003 (n_487, n795);
  and g1004 (n796, n_486, n_487);
  and g1005 (n797, n764, n795);
  not g1006 (n_488, n796);
  not g1007 (n_489, n797);
  and g1008 (n798, n_488, n_489);
  not g1009 (n_490, n763);
  and g1010 (n799, n_490, n798);
  not g1011 (n_491, n799);
  and g1012 (n800, n_490, n_491);
  and g1013 (n801, n798, n_491);
  not g1014 (n_492, n800);
  not g1015 (n_493, n801);
  and g1016 (n802, n_492, n_493);
  not g1017 (n_494, n752);
  not g1018 (n_495, n802);
  and g1019 (n803, n_494, n_495);
  not g1020 (n_496, n803);
  and g1021 (n804, n_494, n_496);
  and g1022 (n805, n_495, n_496);
  not g1023 (n_497, n804);
  not g1024 (n_498, n805);
  and g1025 (n806, n_497, n_498);
  and g1026 (n807, \b[11] , n266);
  and g1027 (n808, \b[9] , n284);
  and g1028 (n809, \b[10] , n261);
  and g1034 (n812, n_437, n_440);
  not g1035 (n_503, \b[11] );
  and g1036 (n813, n_435, n_503);
  and g1037 (n814, \b[10] , \b[11] );
  not g1038 (n_504, n813);
  not g1039 (n_505, n814);
  and g1040 (n815, n_504, n_505);
  not g1041 (n_506, n812);
  and g1042 (n816, n_506, n815);
  not g1043 (n_507, n815);
  and g1044 (n817, n812, n_507);
  not g1045 (n_508, n816);
  not g1046 (n_509, n817);
  and g1047 (n818, n_508, n_509);
  and g1048 (n819, n269, n818);
  not g1051 (n_511, n820);
  and g1052 (n821, \a[2] , n_511);
  not g1053 (n_512, n821);
  and g1054 (n822, \a[2] , n_512);
  and g1055 (n823, n_511, n_512);
  not g1056 (n_513, n822);
  not g1057 (n_514, n823);
  and g1058 (n824, n_513, n_514);
  not g1059 (n_515, n806);
  and g1060 (n825, n_515, n824);
  not g1061 (n_516, n824);
  and g1062 (n826, n806, n_516);
  not g1063 (n_517, n825);
  not g1064 (n_518, n826);
  and g1065 (n827, n_517, n_518);
  not g1066 (n_519, n751);
  not g1067 (n_520, n827);
  and g1068 (n828, n_519, n_520);
  and g1069 (n829, n751, n827);
  not g1070 (n_521, n828);
  not g1071 (n_522, n829);
  and g1072 (\f[11] , n_521, n_522);
  and g1073 (n831, \b[12] , n266);
  and g1074 (n832, \b[10] , n284);
  and g1075 (n833, \b[11] , n261);
  and g1081 (n836, n_505, n_508);
  not g1082 (n_527, \b[12] );
  and g1083 (n837, n_503, n_527);
  and g1084 (n838, \b[11] , \b[12] );
  not g1085 (n_528, n837);
  not g1086 (n_529, n838);
  and g1087 (n839, n_528, n_529);
  not g1088 (n_530, n836);
  and g1089 (n840, n_530, n839);
  not g1090 (n_531, n839);
  and g1091 (n841, n836, n_531);
  not g1092 (n_532, n840);
  not g1093 (n_533, n841);
  and g1094 (n842, n_532, n_533);
  and g1095 (n843, n269, n842);
  not g1098 (n_535, n844);
  and g1099 (n845, \a[2] , n_535);
  not g1100 (n_536, n845);
  and g1101 (n846, \a[2] , n_536);
  and g1102 (n847, n_535, n_536);
  not g1103 (n_537, n846);
  not g1104 (n_538, n847);
  and g1105 (n848, n_537, n_538);
  and g1106 (n849, \b[6] , n511);
  and g1107 (n850, \b[4] , n541);
  and g1108 (n851, \b[5] , n506);
  and g1114 (n854, n459, n514);
  not g1117 (n_543, n855);
  and g1118 (n856, \a[8] , n_543);
  not g1119 (n_544, n856);
  and g1120 (n857, \a[8] , n_544);
  and g1121 (n858, n_543, n_544);
  not g1122 (n_545, n857);
  not g1123 (n_546, n858);
  and g1124 (n859, n_545, n_546);
  not g1125 (n_548, \a[12] );
  and g1126 (n860, \a[11] , n_548);
  and g1127 (n861, n_400, \a[12] );
  not g1128 (n_549, n860);
  not g1129 (n_550, n861);
  and g1130 (n862, n_549, n_550);
  not g1131 (n_551, n862);
  and g1132 (n863, \b[0] , n_551);
  and g1133 (n864, n_473, n863);
  not g1134 (n_552, n863);
  and g1135 (n865, n779, n_552);
  not g1136 (n_553, n864);
  not g1137 (n_554, n865);
  and g1138 (n866, n_553, n_554);
  and g1139 (n867, \b[3] , n700);
  and g1140 (n868, \b[1] , n767);
  and g1141 (n869, \b[2] , n695);
  and g1147 (n872, n318, n703);
  not g1150 (n_559, n873);
  and g1151 (n874, \a[11] , n_559);
  not g1152 (n_560, n874);
  and g1153 (n875, \a[11] , n_560);
  and g1154 (n876, n_559, n_560);
  not g1155 (n_561, n875);
  not g1156 (n_562, n876);
  and g1157 (n877, n_561, n_562);
  not g1158 (n_563, n866);
  not g1159 (n_564, n877);
  and g1160 (n878, n_563, n_564);
  and g1161 (n879, n866, n877);
  not g1162 (n_565, n878);
  not g1163 (n_566, n879);
  and g1164 (n880, n_565, n_566);
  not g1165 (n_567, n859);
  and g1166 (n881, n_567, n880);
  not g1167 (n_568, n881);
  and g1168 (n882, n880, n_568);
  and g1169 (n883, n_567, n_568);
  not g1170 (n_569, n882);
  not g1171 (n_570, n883);
  and g1172 (n884, n_569, n_570);
  and g1173 (n885, n_483, n_488);
  and g1174 (n886, n884, n885);
  not g1175 (n_571, n884);
  not g1176 (n_572, n885);
  and g1177 (n887, n_571, n_572);
  not g1178 (n_573, n886);
  not g1179 (n_574, n887);
  and g1180 (n888, n_573, n_574);
  and g1181 (n889, \b[9] , n362);
  and g1182 (n890, \b[7] , n403);
  and g1183 (n891, \b[8] , n357);
  and g1189 (n894, n365, n651);
  not g1192 (n_579, n895);
  and g1193 (n896, \a[5] , n_579);
  not g1194 (n_580, n896);
  and g1195 (n897, \a[5] , n_580);
  and g1196 (n898, n_579, n_580);
  not g1197 (n_581, n897);
  not g1198 (n_582, n898);
  and g1199 (n899, n_581, n_582);
  not g1200 (n_583, n888);
  and g1201 (n900, n_583, n899);
  not g1202 (n_584, n899);
  and g1203 (n901, n888, n_584);
  not g1204 (n_585, n900);
  not g1205 (n_586, n901);
  and g1206 (n902, n_585, n_586);
  and g1207 (n903, n_491, n_496);
  not g1208 (n_587, n903);
  and g1209 (n904, n902, n_587);
  not g1210 (n_588, n902);
  and g1211 (n905, n_588, n903);
  not g1212 (n_589, n904);
  not g1213 (n_590, n905);
  and g1214 (n906, n_589, n_590);
  not g1215 (n_591, n848);
  and g1216 (n907, n_591, n906);
  not g1217 (n_592, n907);
  and g1218 (n908, n906, n_592);
  and g1219 (n909, n_591, n_592);
  not g1220 (n_593, n908);
  not g1221 (n_594, n909);
  and g1222 (n910, n_593, n_594);
  and g1223 (n911, n_515, n_516);
  not g1224 (n_595, n911);
  and g1225 (n912, n_521, n_595);
  not g1226 (n_596, n910);
  not g1227 (n_597, n912);
  and g1228 (n913, n_596, n_597);
  and g1229 (n914, n910, n912);
  not g1230 (n_598, n913);
  not g1231 (n_599, n914);
  and g1232 (\f[12] , n_598, n_599);
  and g1233 (n916, n_592, n_598);
  and g1234 (n917, n_586, n_589);
  and g1235 (n918, \b[7] , n511);
  and g1236 (n919, \b[5] , n541);
  and g1237 (n920, \b[6] , n506);
  and g1243 (n923, n484, n514);
  not g1246 (n_604, n924);
  and g1247 (n925, \a[8] , n_604);
  not g1248 (n_605, n925);
  and g1249 (n926, \a[8] , n_605);
  and g1250 (n927, n_604, n_605);
  not g1251 (n_606, n926);
  not g1252 (n_607, n927);
  and g1253 (n928, n_606, n_607);
  and g1254 (n929, n779, n863);
  not g1255 (n_608, n929);
  and g1256 (n930, n_565, n_608);
  and g1257 (n931, \b[4] , n700);
  and g1258 (n932, \b[2] , n767);
  and g1259 (n933, \b[3] , n695);
  and g1265 (n936, n346, n703);
  not g1268 (n_613, n937);
  and g1269 (n938, \a[11] , n_613);
  not g1270 (n_614, n938);
  and g1271 (n939, \a[11] , n_614);
  and g1272 (n940, n_613, n_614);
  not g1273 (n_615, n939);
  not g1274 (n_616, n940);
  and g1275 (n941, n_615, n_616);
  and g1276 (n942, \a[14] , n_552);
  and g1277 (n943, n_548, \a[13] );
  not g1278 (n_619, \a[13] );
  and g1279 (n944, \a[12] , n_619);
  not g1280 (n_620, n943);
  not g1281 (n_621, n944);
  and g1282 (n945, n_620, n_621);
  not g1283 (n_622, n945);
  and g1284 (n946, n862, n_622);
  and g1285 (n947, \b[0] , n946);
  and g1286 (n948, n_619, \a[14] );
  not g1287 (n_623, \a[14] );
  and g1288 (n949, \a[13] , n_623);
  not g1289 (n_624, n948);
  not g1290 (n_625, n949);
  and g1291 (n950, n_624, n_625);
  and g1292 (n951, n_551, n950);
  and g1293 (n952, \b[1] , n951);
  not g1294 (n_626, n947);
  not g1295 (n_627, n952);
  and g1296 (n953, n_626, n_627);
  not g1297 (n_628, n950);
  and g1298 (n954, n_551, n_628);
  and g1299 (n955, n_21, n954);
  not g1300 (n_629, n955);
  and g1301 (n956, n953, n_629);
  not g1302 (n_630, n956);
  and g1303 (n957, \a[14] , n_630);
  not g1304 (n_631, n957);
  and g1305 (n958, \a[14] , n_631);
  and g1306 (n959, n_630, n_631);
  not g1307 (n_632, n958);
  not g1308 (n_633, n959);
  and g1309 (n960, n_632, n_633);
  not g1310 (n_634, n960);
  and g1311 (n961, n942, n_634);
  not g1312 (n_635, n942);
  and g1313 (n962, n_635, n960);
  not g1314 (n_636, n961);
  not g1315 (n_637, n962);
  and g1316 (n963, n_636, n_637);
  not g1317 (n_638, n963);
  and g1318 (n964, n941, n_638);
  not g1319 (n_639, n941);
  and g1320 (n965, n_639, n963);
  not g1321 (n_640, n964);
  not g1322 (n_641, n965);
  and g1323 (n966, n_640, n_641);
  not g1324 (n_642, n930);
  and g1325 (n967, n_642, n966);
  not g1326 (n_643, n966);
  and g1327 (n968, n930, n_643);
  not g1328 (n_644, n967);
  not g1329 (n_645, n968);
  and g1330 (n969, n_644, n_645);
  not g1331 (n_646, n928);
  and g1332 (n970, n_646, n969);
  not g1333 (n_647, n970);
  and g1334 (n971, n969, n_647);
  and g1335 (n972, n_646, n_647);
  not g1336 (n_648, n971);
  not g1337 (n_649, n972);
  and g1338 (n973, n_648, n_649);
  and g1339 (n974, n_568, n_574);
  and g1340 (n975, n973, n974);
  not g1341 (n_650, n973);
  not g1342 (n_651, n974);
  and g1343 (n976, n_650, n_651);
  not g1344 (n_652, n975);
  not g1345 (n_653, n976);
  and g1346 (n977, n_652, n_653);
  and g1347 (n978, \b[10] , n362);
  and g1348 (n979, \b[8] , n403);
  and g1349 (n980, \b[9] , n357);
  and g1355 (n983, n365, n738);
  not g1358 (n_658, n984);
  and g1359 (n985, \a[5] , n_658);
  not g1360 (n_659, n985);
  and g1361 (n986, \a[5] , n_659);
  and g1362 (n987, n_658, n_659);
  not g1363 (n_660, n986);
  not g1364 (n_661, n987);
  and g1365 (n988, n_660, n_661);
  not g1366 (n_662, n988);
  and g1367 (n989, n977, n_662);
  not g1368 (n_663, n977);
  and g1369 (n990, n_663, n988);
  not g1370 (n_664, n917);
  not g1371 (n_665, n990);
  and g1372 (n991, n_664, n_665);
  not g1373 (n_666, n989);
  and g1374 (n992, n_666, n991);
  not g1375 (n_667, n992);
  and g1376 (n993, n_664, n_667);
  and g1377 (n994, n_666, n_667);
  and g1378 (n995, n_665, n994);
  not g1379 (n_668, n993);
  not g1380 (n_669, n995);
  and g1381 (n996, n_668, n_669);
  and g1382 (n997, \b[13] , n266);
  and g1383 (n998, \b[11] , n284);
  and g1384 (n999, \b[12] , n261);
  and g1390 (n1002, n_529, n_532);
  not g1391 (n_674, \b[13] );
  and g1392 (n1003, n_527, n_674);
  and g1393 (n1004, \b[12] , \b[13] );
  not g1394 (n_675, n1003);
  not g1395 (n_676, n1004);
  and g1396 (n1005, n_675, n_676);
  not g1397 (n_677, n1002);
  and g1398 (n1006, n_677, n1005);
  not g1399 (n_678, n1005);
  and g1400 (n1007, n1002, n_678);
  not g1401 (n_679, n1006);
  not g1402 (n_680, n1007);
  and g1403 (n1008, n_679, n_680);
  and g1404 (n1009, n269, n1008);
  not g1407 (n_682, n1010);
  and g1408 (n1011, \a[2] , n_682);
  not g1409 (n_683, n1011);
  and g1410 (n1012, \a[2] , n_683);
  and g1411 (n1013, n_682, n_683);
  not g1412 (n_684, n1012);
  not g1413 (n_685, n1013);
  and g1414 (n1014, n_684, n_685);
  not g1415 (n_686, n996);
  and g1416 (n1015, n_686, n1014);
  not g1417 (n_687, n1014);
  and g1418 (n1016, n996, n_687);
  not g1419 (n_688, n1015);
  not g1420 (n_689, n1016);
  and g1421 (n1017, n_688, n_689);
  not g1422 (n_690, n916);
  not g1423 (n_691, n1017);
  and g1424 (n1018, n_690, n_691);
  and g1425 (n1019, n916, n1017);
  not g1426 (n_692, n1018);
  not g1427 (n_693, n1019);
  and g1428 (\f[13] , n_692, n_693);
  and g1429 (n1021, n_686, n_687);
  not g1430 (n_694, n1021);
  and g1431 (n1022, n_692, n_694);
  and g1432 (n1023, \b[14] , n266);
  and g1433 (n1024, \b[12] , n284);
  and g1434 (n1025, \b[13] , n261);
  and g1440 (n1028, n_676, n_679);
  not g1441 (n_699, \b[14] );
  and g1442 (n1029, n_674, n_699);
  and g1443 (n1030, \b[13] , \b[14] );
  not g1444 (n_700, n1029);
  not g1445 (n_701, n1030);
  and g1446 (n1031, n_700, n_701);
  not g1447 (n_702, n1028);
  and g1448 (n1032, n_702, n1031);
  not g1449 (n_703, n1031);
  and g1450 (n1033, n1028, n_703);
  not g1451 (n_704, n1032);
  not g1452 (n_705, n1033);
  and g1453 (n1034, n_704, n_705);
  and g1454 (n1035, n269, n1034);
  not g1457 (n_707, n1036);
  and g1458 (n1037, \a[2] , n_707);
  not g1459 (n_708, n1037);
  and g1460 (n1038, \a[2] , n_708);
  and g1461 (n1039, n_707, n_708);
  not g1462 (n_709, n1038);
  not g1463 (n_710, n1039);
  and g1464 (n1040, n_709, n_710);
  and g1465 (n1041, \b[11] , n362);
  and g1466 (n1042, \b[9] , n403);
  and g1467 (n1043, \b[10] , n357);
  and g1473 (n1046, n365, n818);
  not g1476 (n_715, n1047);
  and g1477 (n1048, \a[5] , n_715);
  not g1478 (n_716, n1048);
  and g1479 (n1049, \a[5] , n_716);
  and g1480 (n1050, n_715, n_716);
  not g1481 (n_717, n1049);
  not g1482 (n_718, n1050);
  and g1483 (n1051, n_717, n_718);
  and g1484 (n1052, n_647, n_653);
  and g1485 (n1053, n_641, n_644);
  and g1486 (n1054, \b[2] , n951);
  and g1487 (n1055, n862, n_628);
  and g1488 (n1056, n945, n1055);
  and g1489 (n1057, \b[0] , n1056);
  and g1490 (n1058, \b[1] , n946);
  and g1496 (n1061, n296, n954);
  not g1499 (n_723, n1062);
  and g1500 (n1063, \a[14] , n_723);
  not g1501 (n_724, n1063);
  and g1502 (n1064, \a[14] , n_724);
  and g1503 (n1065, n_723, n_724);
  not g1504 (n_725, n1064);
  not g1505 (n_726, n1065);
  and g1506 (n1066, n_725, n_726);
  and g1507 (n1067, n_636, n1066);
  not g1508 (n_727, n1066);
  and g1509 (n1068, n961, n_727);
  not g1510 (n_728, n1067);
  not g1511 (n_729, n1068);
  and g1512 (n1069, n_728, n_729);
  and g1513 (n1070, \b[5] , n700);
  and g1514 (n1071, \b[3] , n767);
  and g1515 (n1072, \b[4] , n695);
  and g1521 (n1075, n394, n703);
  not g1524 (n_734, n1076);
  and g1525 (n1077, \a[11] , n_734);
  not g1526 (n_735, n1077);
  and g1527 (n1078, \a[11] , n_735);
  and g1528 (n1079, n_734, n_735);
  not g1529 (n_736, n1078);
  not g1530 (n_737, n1079);
  and g1531 (n1080, n_736, n_737);
  not g1532 (n_738, n1080);
  and g1533 (n1081, n1069, n_738);
  not g1534 (n_739, n1069);
  and g1535 (n1082, n_739, n1080);
  not g1536 (n_740, n1053);
  not g1537 (n_741, n1082);
  and g1538 (n1083, n_740, n_741);
  not g1539 (n_742, n1081);
  and g1540 (n1084, n_742, n1083);
  not g1541 (n_743, n1084);
  and g1542 (n1085, n_740, n_743);
  and g1543 (n1086, n_742, n_743);
  and g1544 (n1087, n_741, n1086);
  not g1545 (n_744, n1085);
  not g1546 (n_745, n1087);
  and g1547 (n1088, n_744, n_745);
  and g1548 (n1089, \b[8] , n511);
  and g1549 (n1090, \b[6] , n541);
  and g1550 (n1091, \b[7] , n506);
  and g1556 (n1094, n514, n585);
  not g1559 (n_750, n1095);
  and g1560 (n1096, \a[8] , n_750);
  not g1561 (n_751, n1096);
  and g1562 (n1097, \a[8] , n_751);
  and g1563 (n1098, n_750, n_751);
  not g1564 (n_752, n1097);
  not g1565 (n_753, n1098);
  and g1566 (n1099, n_752, n_753);
  and g1567 (n1100, n1088, n1099);
  not g1568 (n_754, n1088);
  not g1569 (n_755, n1099);
  and g1570 (n1101, n_754, n_755);
  not g1571 (n_756, n1100);
  not g1572 (n_757, n1101);
  and g1573 (n1102, n_756, n_757);
  not g1574 (n_758, n1052);
  and g1575 (n1103, n_758, n1102);
  not g1576 (n_759, n1102);
  and g1577 (n1104, n1052, n_759);
  not g1578 (n_760, n1103);
  not g1579 (n_761, n1104);
  and g1580 (n1105, n_760, n_761);
  not g1581 (n_762, n1105);
  and g1582 (n1106, n1051, n_762);
  not g1583 (n_763, n1051);
  and g1584 (n1107, n_763, n1105);
  not g1585 (n_764, n1106);
  not g1586 (n_765, n1107);
  and g1587 (n1108, n_764, n_765);
  not g1588 (n_766, n994);
  and g1589 (n1109, n_766, n1108);
  not g1590 (n_767, n1108);
  and g1591 (n1110, n994, n_767);
  not g1592 (n_768, n1109);
  not g1593 (n_769, n1110);
  and g1594 (n1111, n_768, n_769);
  and g1595 (n1112, n1040, n1111);
  not g1596 (n_770, n1040);
  not g1597 (n_771, n1111);
  and g1598 (n1113, n_770, n_771);
  not g1599 (n_772, n1112);
  not g1600 (n_773, n1113);
  and g1601 (n1114, n_772, n_773);
  not g1602 (n_774, n1022);
  not g1603 (n_775, n1114);
  and g1604 (n1115, n_774, n_775);
  and g1605 (n1116, n1022, n1114);
  not g1606 (n_776, n1115);
  not g1607 (n_777, n1116);
  and g1608 (\f[14] , n_776, n_777);
  and g1609 (n1118, n_770, n1111);
  not g1610 (n_778, n1118);
  and g1611 (n1119, n_776, n_778);
  and g1612 (n1120, \b[15] , n266);
  and g1613 (n1121, \b[13] , n284);
  and g1614 (n1122, \b[14] , n261);
  and g1620 (n1125, n_701, n_704);
  not g1621 (n_783, \b[15] );
  and g1622 (n1126, n_699, n_783);
  and g1623 (n1127, \b[14] , \b[15] );
  not g1624 (n_784, n1126);
  not g1625 (n_785, n1127);
  and g1626 (n1128, n_784, n_785);
  not g1627 (n_786, n1125);
  and g1628 (n1129, n_786, n1128);
  not g1629 (n_787, n1128);
  and g1630 (n1130, n1125, n_787);
  not g1631 (n_788, n1129);
  not g1632 (n_789, n1130);
  and g1633 (n1131, n_788, n_789);
  and g1634 (n1132, n269, n1131);
  not g1637 (n_791, n1133);
  and g1638 (n1134, \a[2] , n_791);
  not g1639 (n_792, n1134);
  and g1640 (n1135, \a[2] , n_792);
  and g1641 (n1136, n_791, n_792);
  not g1642 (n_793, n1135);
  not g1643 (n_794, n1136);
  and g1644 (n1137, n_793, n_794);
  and g1645 (n1138, n_765, n_768);
  and g1646 (n1139, \b[12] , n362);
  and g1647 (n1140, \b[10] , n403);
  and g1648 (n1141, \b[11] , n357);
  and g1654 (n1144, n365, n842);
  not g1657 (n_799, n1145);
  and g1658 (n1146, \a[5] , n_799);
  not g1659 (n_800, n1146);
  and g1660 (n1147, \a[5] , n_800);
  and g1661 (n1148, n_799, n_800);
  not g1662 (n_801, n1147);
  not g1663 (n_802, n1148);
  and g1664 (n1149, n_801, n_802);
  and g1665 (n1150, n_757, n_760);
  and g1666 (n1151, \b[9] , n511);
  and g1667 (n1152, \b[7] , n541);
  and g1668 (n1153, \b[8] , n506);
  and g1674 (n1156, n514, n651);
  not g1677 (n_807, n1157);
  and g1678 (n1158, \a[8] , n_807);
  not g1679 (n_808, n1158);
  and g1680 (n1159, \a[8] , n_808);
  and g1681 (n1160, n_807, n_808);
  not g1682 (n_809, n1159);
  not g1683 (n_810, n1160);
  and g1684 (n1161, n_809, n_810);
  and g1685 (n1162, \b[6] , n700);
  and g1686 (n1163, \b[4] , n767);
  and g1687 (n1164, \b[5] , n695);
  and g1693 (n1167, n459, n703);
  not g1696 (n_815, n1168);
  and g1697 (n1169, \a[11] , n_815);
  not g1698 (n_816, n1169);
  and g1699 (n1170, \a[11] , n_816);
  and g1700 (n1171, n_815, n_816);
  not g1701 (n_817, n1170);
  not g1702 (n_818, n1171);
  and g1703 (n1172, n_817, n_818);
  not g1704 (n_820, \a[15] );
  and g1705 (n1173, \a[14] , n_820);
  and g1706 (n1174, n_623, \a[15] );
  not g1707 (n_821, n1173);
  not g1708 (n_822, n1174);
  and g1709 (n1175, n_821, n_822);
  not g1710 (n_823, n1175);
  and g1711 (n1176, \b[0] , n_823);
  and g1712 (n1177, n_729, n1176);
  not g1713 (n_824, n1176);
  and g1714 (n1178, n1068, n_824);
  not g1715 (n_825, n1177);
  not g1716 (n_826, n1178);
  and g1717 (n1179, n_825, n_826);
  and g1718 (n1180, \b[3] , n951);
  and g1719 (n1181, \b[1] , n1056);
  and g1720 (n1182, \b[2] , n946);
  and g1726 (n1185, n318, n954);
  not g1729 (n_831, n1186);
  and g1730 (n1187, \a[14] , n_831);
  not g1731 (n_832, n1187);
  and g1732 (n1188, \a[14] , n_832);
  and g1733 (n1189, n_831, n_832);
  not g1734 (n_833, n1188);
  not g1735 (n_834, n1189);
  and g1736 (n1190, n_833, n_834);
  not g1737 (n_835, n1179);
  not g1738 (n_836, n1190);
  and g1739 (n1191, n_835, n_836);
  and g1740 (n1192, n1179, n1190);
  not g1741 (n_837, n1191);
  not g1742 (n_838, n1192);
  and g1743 (n1193, n_837, n_838);
  not g1744 (n_839, n1172);
  and g1745 (n1194, n_839, n1193);
  not g1746 (n_840, n1194);
  and g1747 (n1195, n1193, n_840);
  and g1748 (n1196, n_839, n_840);
  not g1749 (n_841, n1195);
  not g1750 (n_842, n1196);
  and g1751 (n1197, n_841, n_842);
  not g1752 (n_843, n1086);
  not g1753 (n_844, n1197);
  and g1754 (n1198, n_843, n_844);
  and g1755 (n1199, n1086, n1197);
  not g1756 (n_845, n1198);
  not g1757 (n_846, n1199);
  and g1758 (n1200, n_845, n_846);
  not g1759 (n_847, n1161);
  and g1760 (n1201, n_847, n1200);
  not g1761 (n_848, n1201);
  and g1762 (n1202, n_847, n_848);
  and g1763 (n1203, n1200, n_848);
  not g1764 (n_849, n1202);
  not g1765 (n_850, n1203);
  and g1766 (n1204, n_849, n_850);
  not g1767 (n_851, n1150);
  not g1768 (n_852, n1204);
  and g1769 (n1205, n_851, n_852);
  and g1770 (n1206, n1150, n_850);
  and g1771 (n1207, n_849, n1206);
  not g1772 (n_853, n1205);
  not g1773 (n_854, n1207);
  and g1774 (n1208, n_853, n_854);
  not g1775 (n_855, n1149);
  and g1776 (n1209, n_855, n1208);
  not g1777 (n_856, n1209);
  and g1778 (n1210, n_855, n_856);
  and g1779 (n1211, n1208, n_856);
  not g1780 (n_857, n1210);
  not g1781 (n_858, n1211);
  and g1782 (n1212, n_857, n_858);
  not g1783 (n_859, n1138);
  not g1784 (n_860, n1212);
  and g1785 (n1213, n_859, n_860);
  and g1786 (n1214, n1138, n_858);
  and g1787 (n1215, n_857, n1214);
  not g1788 (n_861, n1213);
  not g1789 (n_862, n1215);
  and g1790 (n1216, n_861, n_862);
  not g1791 (n_863, n1137);
  and g1792 (n1217, n_863, n1216);
  not g1793 (n_864, n1217);
  and g1794 (n1218, n_863, n_864);
  and g1795 (n1219, n1216, n_864);
  not g1796 (n_865, n1218);
  not g1797 (n_866, n1219);
  and g1798 (n1220, n_865, n_866);
  not g1799 (n_867, n1119);
  not g1800 (n_868, n1220);
  and g1801 (n1221, n_867, n_868);
  and g1802 (n1222, n1119, n_866);
  and g1803 (n1223, n_865, n1222);
  not g1804 (n_869, n1221);
  not g1805 (n_870, n1223);
  and g1806 (\f[15] , n_869, n_870);
  and g1807 (n1225, n_864, n_869);
  and g1808 (n1226, \b[16] , n266);
  and g1809 (n1227, \b[14] , n284);
  and g1810 (n1228, \b[15] , n261);
  and g1816 (n1231, n_785, n_788);
  not g1817 (n_875, \b[16] );
  and g1818 (n1232, n_783, n_875);
  and g1819 (n1233, \b[15] , \b[16] );
  not g1820 (n_876, n1232);
  not g1821 (n_877, n1233);
  and g1822 (n1234, n_876, n_877);
  not g1823 (n_878, n1231);
  and g1824 (n1235, n_878, n1234);
  not g1825 (n_879, n1234);
  and g1826 (n1236, n1231, n_879);
  not g1827 (n_880, n1235);
  not g1828 (n_881, n1236);
  and g1829 (n1237, n_880, n_881);
  and g1830 (n1238, n269, n1237);
  not g1833 (n_883, n1239);
  and g1834 (n1240, \a[2] , n_883);
  not g1835 (n_884, n1240);
  and g1836 (n1241, \a[2] , n_884);
  and g1837 (n1242, n_883, n_884);
  not g1838 (n_885, n1241);
  not g1839 (n_886, n1242);
  and g1840 (n1243, n_885, n_886);
  and g1841 (n1244, n_856, n_861);
  and g1842 (n1245, \b[13] , n362);
  and g1843 (n1246, \b[11] , n403);
  and g1844 (n1247, \b[12] , n357);
  and g1850 (n1250, n365, n1008);
  not g1853 (n_891, n1251);
  and g1854 (n1252, \a[5] , n_891);
  not g1855 (n_892, n1252);
  and g1856 (n1253, \a[5] , n_892);
  and g1857 (n1254, n_891, n_892);
  not g1858 (n_893, n1253);
  not g1859 (n_894, n1254);
  and g1860 (n1255, n_893, n_894);
  and g1861 (n1256, n_848, n_853);
  and g1862 (n1257, \b[10] , n511);
  and g1863 (n1258, \b[8] , n541);
  and g1864 (n1259, \b[9] , n506);
  and g1870 (n1262, n514, n738);
  not g1873 (n_899, n1263);
  and g1874 (n1264, \a[8] , n_899);
  not g1875 (n_900, n1264);
  and g1876 (n1265, \a[8] , n_900);
  and g1877 (n1266, n_899, n_900);
  not g1878 (n_901, n1265);
  not g1879 (n_902, n1266);
  and g1880 (n1267, n_901, n_902);
  and g1881 (n1268, n_840, n_845);
  and g1882 (n1269, \b[7] , n700);
  and g1883 (n1270, \b[5] , n767);
  and g1884 (n1271, \b[6] , n695);
  and g1890 (n1274, n484, n703);
  not g1893 (n_907, n1275);
  and g1894 (n1276, \a[11] , n_907);
  not g1895 (n_908, n1276);
  and g1896 (n1277, \a[11] , n_908);
  and g1897 (n1278, n_907, n_908);
  not g1898 (n_909, n1277);
  not g1899 (n_910, n1278);
  and g1900 (n1279, n_909, n_910);
  and g1901 (n1280, n1068, n1176);
  not g1902 (n_911, n1280);
  and g1903 (n1281, n_837, n_911);
  and g1904 (n1282, \b[4] , n951);
  and g1905 (n1283, \b[2] , n1056);
  and g1906 (n1284, \b[3] , n946);
  and g1912 (n1287, n346, n954);
  not g1915 (n_916, n1288);
  and g1916 (n1289, \a[14] , n_916);
  not g1917 (n_917, n1289);
  and g1918 (n1290, \a[14] , n_917);
  and g1919 (n1291, n_916, n_917);
  not g1920 (n_918, n1290);
  not g1921 (n_919, n1291);
  and g1922 (n1292, n_918, n_919);
  and g1923 (n1293, \a[17] , n_824);
  and g1924 (n1294, n_820, \a[16] );
  not g1925 (n_922, \a[16] );
  and g1926 (n1295, \a[15] , n_922);
  not g1927 (n_923, n1294);
  not g1928 (n_924, n1295);
  and g1929 (n1296, n_923, n_924);
  not g1930 (n_925, n1296);
  and g1931 (n1297, n1175, n_925);
  and g1932 (n1298, \b[0] , n1297);
  and g1933 (n1299, n_922, \a[17] );
  not g1934 (n_926, \a[17] );
  and g1935 (n1300, \a[16] , n_926);
  not g1936 (n_927, n1299);
  not g1937 (n_928, n1300);
  and g1938 (n1301, n_927, n_928);
  and g1939 (n1302, n_823, n1301);
  and g1940 (n1303, \b[1] , n1302);
  not g1941 (n_929, n1298);
  not g1942 (n_930, n1303);
  and g1943 (n1304, n_929, n_930);
  not g1944 (n_931, n1301);
  and g1945 (n1305, n_823, n_931);
  and g1946 (n1306, n_21, n1305);
  not g1947 (n_932, n1306);
  and g1948 (n1307, n1304, n_932);
  not g1949 (n_933, n1307);
  and g1950 (n1308, \a[17] , n_933);
  not g1951 (n_934, n1308);
  and g1952 (n1309, \a[17] , n_934);
  and g1953 (n1310, n_933, n_934);
  not g1954 (n_935, n1309);
  not g1955 (n_936, n1310);
  and g1956 (n1311, n_935, n_936);
  not g1957 (n_937, n1311);
  and g1958 (n1312, n1293, n_937);
  not g1959 (n_938, n1293);
  and g1960 (n1313, n_938, n1311);
  not g1961 (n_939, n1312);
  not g1962 (n_940, n1313);
  and g1963 (n1314, n_939, n_940);
  not g1964 (n_941, n1314);
  and g1965 (n1315, n1292, n_941);
  not g1966 (n_942, n1292);
  and g1967 (n1316, n_942, n1314);
  not g1968 (n_943, n1315);
  not g1969 (n_944, n1316);
  and g1970 (n1317, n_943, n_944);
  not g1971 (n_945, n1281);
  and g1972 (n1318, n_945, n1317);
  not g1973 (n_946, n1317);
  and g1974 (n1319, n1281, n_946);
  not g1975 (n_947, n1318);
  not g1976 (n_948, n1319);
  and g1977 (n1320, n_947, n_948);
  not g1978 (n_949, n1320);
  and g1979 (n1321, n1279, n_949);
  not g1980 (n_950, n1279);
  and g1981 (n1322, n_950, n1320);
  not g1982 (n_951, n1321);
  not g1983 (n_952, n1322);
  and g1984 (n1323, n_951, n_952);
  not g1985 (n_953, n1268);
  and g1986 (n1324, n_953, n1323);
  not g1987 (n_954, n1323);
  and g1988 (n1325, n1268, n_954);
  not g1989 (n_955, n1324);
  not g1990 (n_956, n1325);
  and g1991 (n1326, n_955, n_956);
  not g1992 (n_957, n1326);
  and g1993 (n1327, n1267, n_957);
  not g1994 (n_958, n1267);
  and g1995 (n1328, n_958, n1326);
  not g1996 (n_959, n1327);
  not g1997 (n_960, n1328);
  and g1998 (n1329, n_959, n_960);
  not g1999 (n_961, n1256);
  and g2000 (n1330, n_961, n1329);
  not g2001 (n_962, n1329);
  and g2002 (n1331, n1256, n_962);
  not g2003 (n_963, n1330);
  not g2004 (n_964, n1331);
  and g2005 (n1332, n_963, n_964);
  not g2006 (n_965, n1332);
  and g2007 (n1333, n1255, n_965);
  not g2008 (n_966, n1255);
  and g2009 (n1334, n_966, n1332);
  not g2010 (n_967, n1333);
  not g2011 (n_968, n1334);
  and g2012 (n1335, n_967, n_968);
  not g2013 (n_969, n1244);
  and g2014 (n1336, n_969, n1335);
  not g2015 (n_970, n1335);
  and g2016 (n1337, n1244, n_970);
  not g2017 (n_971, n1336);
  not g2018 (n_972, n1337);
  and g2019 (n1338, n_971, n_972);
  and g2020 (n1339, n1243, n1338);
  not g2021 (n_973, n1243);
  not g2022 (n_974, n1338);
  and g2023 (n1340, n_973, n_974);
  not g2024 (n_975, n1339);
  not g2025 (n_976, n1340);
  and g2026 (n1341, n_975, n_976);
  not g2027 (n_977, n1225);
  not g2028 (n_978, n1341);
  and g2029 (n1342, n_977, n_978);
  and g2030 (n1343, n1225, n1341);
  not g2031 (n_979, n1342);
  not g2032 (n_980, n1343);
  and g2033 (\f[16] , n_979, n_980);
  and g2034 (n1345, \b[17] , n266);
  and g2035 (n1346, \b[15] , n284);
  and g2036 (n1347, \b[16] , n261);
  and g2042 (n1350, n_877, n_880);
  not g2043 (n_985, \b[17] );
  and g2044 (n1351, n_875, n_985);
  and g2045 (n1352, \b[16] , \b[17] );
  not g2046 (n_986, n1351);
  not g2047 (n_987, n1352);
  and g2048 (n1353, n_986, n_987);
  not g2049 (n_988, n1350);
  and g2050 (n1354, n_988, n1353);
  not g2051 (n_989, n1353);
  and g2052 (n1355, n1350, n_989);
  not g2053 (n_990, n1354);
  not g2054 (n_991, n1355);
  and g2055 (n1356, n_990, n_991);
  and g2056 (n1357, n269, n1356);
  not g2059 (n_993, n1358);
  and g2060 (n1359, \a[2] , n_993);
  not g2061 (n_994, n1359);
  and g2062 (n1360, \a[2] , n_994);
  and g2063 (n1361, n_993, n_994);
  not g2064 (n_995, n1360);
  not g2065 (n_996, n1361);
  and g2066 (n1362, n_995, n_996);
  and g2067 (n1363, n_968, n_971);
  and g2068 (n1364, \b[14] , n362);
  and g2069 (n1365, \b[12] , n403);
  and g2070 (n1366, \b[13] , n357);
  and g2076 (n1369, n365, n1034);
  not g2079 (n_1001, n1370);
  and g2080 (n1371, \a[5] , n_1001);
  not g2081 (n_1002, n1371);
  and g2082 (n1372, \a[5] , n_1002);
  and g2083 (n1373, n_1001, n_1002);
  not g2084 (n_1003, n1372);
  not g2085 (n_1004, n1373);
  and g2086 (n1374, n_1003, n_1004);
  and g2087 (n1375, n_960, n_963);
  and g2088 (n1376, \b[11] , n511);
  and g2089 (n1377, \b[9] , n541);
  and g2090 (n1378, \b[10] , n506);
  and g2096 (n1381, n514, n818);
  not g2099 (n_1009, n1382);
  and g2100 (n1383, \a[8] , n_1009);
  not g2101 (n_1010, n1383);
  and g2102 (n1384, \a[8] , n_1010);
  and g2103 (n1385, n_1009, n_1010);
  not g2104 (n_1011, n1384);
  not g2105 (n_1012, n1385);
  and g2106 (n1386, n_1011, n_1012);
  and g2107 (n1387, n_952, n_955);
  and g2108 (n1388, n_944, n_947);
  and g2109 (n1389, \b[2] , n1302);
  and g2110 (n1390, n1175, n_931);
  and g2111 (n1391, n1296, n1390);
  and g2112 (n1392, \b[0] , n1391);
  and g2113 (n1393, \b[1] , n1297);
  and g2119 (n1396, n296, n1305);
  not g2122 (n_1017, n1397);
  and g2123 (n1398, \a[17] , n_1017);
  not g2124 (n_1018, n1398);
  and g2125 (n1399, \a[17] , n_1018);
  and g2126 (n1400, n_1017, n_1018);
  not g2127 (n_1019, n1399);
  not g2128 (n_1020, n1400);
  and g2129 (n1401, n_1019, n_1020);
  and g2130 (n1402, n_939, n1401);
  not g2131 (n_1021, n1401);
  and g2132 (n1403, n1312, n_1021);
  not g2133 (n_1022, n1402);
  not g2134 (n_1023, n1403);
  and g2135 (n1404, n_1022, n_1023);
  and g2136 (n1405, \b[5] , n951);
  and g2137 (n1406, \b[3] , n1056);
  and g2138 (n1407, \b[4] , n946);
  and g2144 (n1410, n394, n954);
  not g2147 (n_1028, n1411);
  and g2148 (n1412, \a[14] , n_1028);
  not g2149 (n_1029, n1412);
  and g2150 (n1413, \a[14] , n_1029);
  and g2151 (n1414, n_1028, n_1029);
  not g2152 (n_1030, n1413);
  not g2153 (n_1031, n1414);
  and g2154 (n1415, n_1030, n_1031);
  not g2155 (n_1032, n1415);
  and g2156 (n1416, n1404, n_1032);
  not g2157 (n_1033, n1404);
  and g2158 (n1417, n_1033, n1415);
  not g2159 (n_1034, n1388);
  not g2160 (n_1035, n1417);
  and g2161 (n1418, n_1034, n_1035);
  not g2162 (n_1036, n1416);
  and g2163 (n1419, n_1036, n1418);
  not g2164 (n_1037, n1419);
  and g2165 (n1420, n_1034, n_1037);
  and g2166 (n1421, n_1036, n_1037);
  and g2167 (n1422, n_1035, n1421);
  not g2168 (n_1038, n1420);
  not g2169 (n_1039, n1422);
  and g2170 (n1423, n_1038, n_1039);
  and g2171 (n1424, \b[8] , n700);
  and g2172 (n1425, \b[6] , n767);
  and g2173 (n1426, \b[7] , n695);
  and g2179 (n1429, n585, n703);
  not g2182 (n_1044, n1430);
  and g2183 (n1431, \a[11] , n_1044);
  not g2184 (n_1045, n1431);
  and g2185 (n1432, \a[11] , n_1045);
  and g2186 (n1433, n_1044, n_1045);
  not g2187 (n_1046, n1432);
  not g2188 (n_1047, n1433);
  and g2189 (n1434, n_1046, n_1047);
  and g2190 (n1435, n1423, n1434);
  not g2191 (n_1048, n1423);
  not g2192 (n_1049, n1434);
  and g2193 (n1436, n_1048, n_1049);
  not g2194 (n_1050, n1435);
  not g2195 (n_1051, n1436);
  and g2196 (n1437, n_1050, n_1051);
  not g2197 (n_1052, n1387);
  and g2198 (n1438, n_1052, n1437);
  not g2199 (n_1053, n1437);
  and g2200 (n1439, n1387, n_1053);
  not g2201 (n_1054, n1438);
  not g2202 (n_1055, n1439);
  and g2203 (n1440, n_1054, n_1055);
  not g2204 (n_1056, n1440);
  and g2205 (n1441, n1386, n_1056);
  not g2206 (n_1057, n1386);
  and g2207 (n1442, n_1057, n1440);
  not g2208 (n_1058, n1441);
  not g2209 (n_1059, n1442);
  and g2210 (n1443, n_1058, n_1059);
  not g2211 (n_1060, n1375);
  and g2212 (n1444, n_1060, n1443);
  not g2213 (n_1061, n1443);
  and g2214 (n1445, n1375, n_1061);
  not g2215 (n_1062, n1444);
  not g2216 (n_1063, n1445);
  and g2217 (n1446, n_1062, n_1063);
  not g2218 (n_1064, n1446);
  and g2219 (n1447, n1374, n_1064);
  not g2220 (n_1065, n1374);
  and g2221 (n1448, n_1065, n1446);
  not g2222 (n_1066, n1447);
  not g2223 (n_1067, n1448);
  and g2224 (n1449, n_1066, n_1067);
  not g2225 (n_1068, n1363);
  and g2226 (n1450, n_1068, n1449);
  not g2227 (n_1069, n1449);
  and g2228 (n1451, n1363, n_1069);
  not g2229 (n_1070, n1450);
  not g2230 (n_1071, n1451);
  and g2231 (n1452, n_1070, n_1071);
  not g2232 (n_1072, n1362);
  and g2233 (n1453, n_1072, n1452);
  not g2234 (n_1073, n1453);
  and g2235 (n1454, n1452, n_1073);
  and g2236 (n1455, n_1072, n_1073);
  not g2237 (n_1074, n1454);
  not g2238 (n_1075, n1455);
  and g2239 (n1456, n_1074, n_1075);
  and g2240 (n1457, n_973, n1338);
  not g2241 (n_1076, n1457);
  and g2242 (n1458, n_979, n_1076);
  not g2243 (n_1077, n1456);
  not g2244 (n_1078, n1458);
  and g2245 (n1459, n_1077, n_1078);
  and g2246 (n1460, n1456, n1458);
  not g2247 (n_1079, n1459);
  not g2248 (n_1080, n1460);
  and g2249 (\f[17] , n_1079, n_1080);
  and g2250 (n1462, n_1067, n_1070);
  and g2251 (n1463, \b[15] , n362);
  and g2252 (n1464, \b[13] , n403);
  and g2253 (n1465, \b[14] , n357);
  and g2259 (n1468, n365, n1131);
  not g2262 (n_1085, n1469);
  and g2263 (n1470, \a[5] , n_1085);
  not g2264 (n_1086, n1470);
  and g2265 (n1471, \a[5] , n_1086);
  and g2266 (n1472, n_1085, n_1086);
  not g2267 (n_1087, n1471);
  not g2268 (n_1088, n1472);
  and g2269 (n1473, n_1087, n_1088);
  and g2270 (n1474, n_1059, n_1062);
  and g2271 (n1475, \b[12] , n511);
  and g2272 (n1476, \b[10] , n541);
  and g2273 (n1477, \b[11] , n506);
  and g2279 (n1480, n514, n842);
  not g2282 (n_1093, n1481);
  and g2283 (n1482, \a[8] , n_1093);
  not g2284 (n_1094, n1482);
  and g2285 (n1483, \a[8] , n_1094);
  and g2286 (n1484, n_1093, n_1094);
  not g2287 (n_1095, n1483);
  not g2288 (n_1096, n1484);
  and g2289 (n1485, n_1095, n_1096);
  and g2290 (n1486, n_1051, n_1054);
  and g2291 (n1487, \b[6] , n951);
  and g2292 (n1488, \b[4] , n1056);
  and g2293 (n1489, \b[5] , n946);
  and g2299 (n1492, n459, n954);
  not g2302 (n_1101, n1493);
  and g2303 (n1494, \a[14] , n_1101);
  not g2304 (n_1102, n1494);
  and g2305 (n1495, \a[14] , n_1102);
  and g2306 (n1496, n_1101, n_1102);
  not g2307 (n_1103, n1495);
  not g2308 (n_1104, n1496);
  and g2309 (n1497, n_1103, n_1104);
  not g2310 (n_1106, \a[18] );
  and g2311 (n1498, \a[17] , n_1106);
  and g2312 (n1499, n_926, \a[18] );
  not g2313 (n_1107, n1498);
  not g2314 (n_1108, n1499);
  and g2315 (n1500, n_1107, n_1108);
  not g2316 (n_1109, n1500);
  and g2317 (n1501, \b[0] , n_1109);
  and g2318 (n1502, n_1023, n1501);
  not g2319 (n_1110, n1501);
  and g2320 (n1503, n1403, n_1110);
  not g2321 (n_1111, n1502);
  not g2322 (n_1112, n1503);
  and g2323 (n1504, n_1111, n_1112);
  and g2324 (n1505, \b[3] , n1302);
  and g2325 (n1506, \b[1] , n1391);
  and g2326 (n1507, \b[2] , n1297);
  and g2332 (n1510, n318, n1305);
  not g2335 (n_1117, n1511);
  and g2336 (n1512, \a[17] , n_1117);
  not g2337 (n_1118, n1512);
  and g2338 (n1513, \a[17] , n_1118);
  and g2339 (n1514, n_1117, n_1118);
  not g2340 (n_1119, n1513);
  not g2341 (n_1120, n1514);
  and g2342 (n1515, n_1119, n_1120);
  not g2343 (n_1121, n1504);
  not g2344 (n_1122, n1515);
  and g2345 (n1516, n_1121, n_1122);
  and g2346 (n1517, n1504, n1515);
  not g2347 (n_1123, n1516);
  not g2348 (n_1124, n1517);
  and g2349 (n1518, n_1123, n_1124);
  not g2350 (n_1125, n1497);
  and g2351 (n1519, n_1125, n1518);
  not g2352 (n_1126, n1519);
  and g2353 (n1520, n1518, n_1126);
  and g2354 (n1521, n_1125, n_1126);
  not g2355 (n_1127, n1520);
  not g2356 (n_1128, n1521);
  and g2357 (n1522, n_1127, n_1128);
  not g2358 (n_1129, n1421);
  and g2359 (n1523, n_1129, n1522);
  not g2360 (n_1130, n1522);
  and g2361 (n1524, n1421, n_1130);
  not g2362 (n_1131, n1523);
  not g2363 (n_1132, n1524);
  and g2364 (n1525, n_1131, n_1132);
  and g2365 (n1526, \b[9] , n700);
  and g2366 (n1527, \b[7] , n767);
  and g2367 (n1528, \b[8] , n695);
  and g2373 (n1531, n651, n703);
  not g2376 (n_1137, n1532);
  and g2377 (n1533, \a[11] , n_1137);
  not g2378 (n_1138, n1533);
  and g2379 (n1534, \a[11] , n_1138);
  and g2380 (n1535, n_1137, n_1138);
  not g2381 (n_1139, n1534);
  not g2382 (n_1140, n1535);
  and g2383 (n1536, n_1139, n_1140);
  not g2384 (n_1141, n1525);
  not g2385 (n_1142, n1536);
  and g2386 (n1537, n_1141, n_1142);
  and g2387 (n1538, n1525, n1536);
  not g2388 (n_1143, n1537);
  not g2389 (n_1144, n1538);
  and g2390 (n1539, n_1143, n_1144);
  not g2391 (n_1145, n1486);
  and g2392 (n1540, n_1145, n1539);
  not g2393 (n_1146, n1539);
  and g2394 (n1541, n1486, n_1146);
  not g2395 (n_1147, n1540);
  not g2396 (n_1148, n1541);
  and g2397 (n1542, n_1147, n_1148);
  not g2398 (n_1149, n1542);
  and g2399 (n1543, n1485, n_1149);
  not g2400 (n_1150, n1485);
  and g2401 (n1544, n_1150, n1542);
  not g2402 (n_1151, n1543);
  not g2403 (n_1152, n1544);
  and g2404 (n1545, n_1151, n_1152);
  not g2405 (n_1153, n1474);
  and g2406 (n1546, n_1153, n1545);
  not g2407 (n_1154, n1545);
  and g2408 (n1547, n1474, n_1154);
  not g2409 (n_1155, n1546);
  not g2410 (n_1156, n1547);
  and g2411 (n1548, n_1155, n_1156);
  not g2412 (n_1157, n1473);
  and g2413 (n1549, n_1157, n1548);
  not g2414 (n_1158, n1548);
  and g2415 (n1550, n1473, n_1158);
  not g2416 (n_1159, n1549);
  not g2417 (n_1160, n1550);
  and g2418 (n1551, n_1159, n_1160);
  not g2419 (n_1161, n1462);
  and g2420 (n1552, n_1161, n1551);
  not g2421 (n_1162, n1551);
  and g2422 (n1553, n1462, n_1162);
  not g2423 (n_1163, n1552);
  not g2424 (n_1164, n1553);
  and g2425 (n1554, n_1163, n_1164);
  and g2426 (n1555, \b[18] , n266);
  and g2427 (n1556, \b[16] , n284);
  and g2428 (n1557, \b[17] , n261);
  and g2434 (n1560, n_987, n_990);
  not g2435 (n_1169, \b[18] );
  and g2436 (n1561, n_985, n_1169);
  and g2437 (n1562, \b[17] , \b[18] );
  not g2438 (n_1170, n1561);
  not g2439 (n_1171, n1562);
  and g2440 (n1563, n_1170, n_1171);
  not g2441 (n_1172, n1560);
  and g2442 (n1564, n_1172, n1563);
  not g2443 (n_1173, n1563);
  and g2444 (n1565, n1560, n_1173);
  not g2445 (n_1174, n1564);
  not g2446 (n_1175, n1565);
  and g2447 (n1566, n_1174, n_1175);
  and g2448 (n1567, n269, n1566);
  not g2451 (n_1177, n1568);
  and g2452 (n1569, \a[2] , n_1177);
  not g2453 (n_1178, n1569);
  and g2454 (n1570, \a[2] , n_1178);
  and g2455 (n1571, n_1177, n_1178);
  not g2456 (n_1179, n1570);
  not g2457 (n_1180, n1571);
  and g2458 (n1572, n_1179, n_1180);
  not g2459 (n_1181, n1572);
  and g2460 (n1573, n1554, n_1181);
  not g2461 (n_1182, n1573);
  and g2462 (n1574, n1554, n_1182);
  and g2463 (n1575, n_1181, n_1182);
  not g2464 (n_1183, n1574);
  not g2465 (n_1184, n1575);
  and g2466 (n1576, n_1183, n_1184);
  and g2467 (n1577, n_1073, n_1079);
  not g2468 (n_1185, n1576);
  not g2469 (n_1186, n1577);
  and g2470 (n1578, n_1185, n_1186);
  and g2471 (n1579, n1576, n1577);
  not g2472 (n_1187, n1578);
  not g2473 (n_1188, n1579);
  and g2474 (\f[18] , n_1187, n_1188);
  and g2475 (n1581, \b[16] , n362);
  and g2476 (n1582, \b[14] , n403);
  and g2477 (n1583, \b[15] , n357);
  and g2483 (n1586, n365, n1237);
  not g2486 (n_1193, n1587);
  and g2487 (n1588, \a[5] , n_1193);
  not g2488 (n_1194, n1588);
  and g2489 (n1589, \a[5] , n_1194);
  and g2490 (n1590, n_1193, n_1194);
  not g2491 (n_1195, n1589);
  not g2492 (n_1196, n1590);
  and g2493 (n1591, n_1195, n_1196);
  and g2494 (n1592, n_1129, n_1130);
  not g2495 (n_1197, n1592);
  and g2496 (n1593, n_1126, n_1197);
  and g2497 (n1594, \b[7] , n951);
  and g2498 (n1595, \b[5] , n1056);
  and g2499 (n1596, \b[6] , n946);
  and g2505 (n1599, n484, n954);
  not g2508 (n_1202, n1600);
  and g2509 (n1601, \a[14] , n_1202);
  not g2510 (n_1203, n1601);
  and g2511 (n1602, \a[14] , n_1203);
  and g2512 (n1603, n_1202, n_1203);
  not g2513 (n_1204, n1602);
  not g2514 (n_1205, n1603);
  and g2515 (n1604, n_1204, n_1205);
  and g2516 (n1605, n1403, n1501);
  not g2517 (n_1206, n1605);
  and g2518 (n1606, n_1123, n_1206);
  and g2519 (n1607, \b[4] , n1302);
  and g2520 (n1608, \b[2] , n1391);
  and g2521 (n1609, \b[3] , n1297);
  and g2527 (n1612, n346, n1305);
  not g2530 (n_1211, n1613);
  and g2531 (n1614, \a[17] , n_1211);
  not g2532 (n_1212, n1614);
  and g2533 (n1615, \a[17] , n_1212);
  and g2534 (n1616, n_1211, n_1212);
  not g2535 (n_1213, n1615);
  not g2536 (n_1214, n1616);
  and g2537 (n1617, n_1213, n_1214);
  and g2538 (n1618, \a[20] , n_1110);
  and g2539 (n1619, n_1106, \a[19] );
  not g2540 (n_1217, \a[19] );
  and g2541 (n1620, \a[18] , n_1217);
  not g2542 (n_1218, n1619);
  not g2543 (n_1219, n1620);
  and g2544 (n1621, n_1218, n_1219);
  not g2545 (n_1220, n1621);
  and g2546 (n1622, n1500, n_1220);
  and g2547 (n1623, \b[0] , n1622);
  and g2548 (n1624, n_1217, \a[20] );
  not g2549 (n_1221, \a[20] );
  and g2550 (n1625, \a[19] , n_1221);
  not g2551 (n_1222, n1624);
  not g2552 (n_1223, n1625);
  and g2553 (n1626, n_1222, n_1223);
  and g2554 (n1627, n_1109, n1626);
  and g2555 (n1628, \b[1] , n1627);
  not g2556 (n_1224, n1623);
  not g2557 (n_1225, n1628);
  and g2558 (n1629, n_1224, n_1225);
  not g2559 (n_1226, n1626);
  and g2560 (n1630, n_1109, n_1226);
  and g2561 (n1631, n_21, n1630);
  not g2562 (n_1227, n1631);
  and g2563 (n1632, n1629, n_1227);
  not g2564 (n_1228, n1632);
  and g2565 (n1633, \a[20] , n_1228);
  not g2566 (n_1229, n1633);
  and g2567 (n1634, \a[20] , n_1229);
  and g2568 (n1635, n_1228, n_1229);
  not g2569 (n_1230, n1634);
  not g2570 (n_1231, n1635);
  and g2571 (n1636, n_1230, n_1231);
  not g2572 (n_1232, n1636);
  and g2573 (n1637, n1618, n_1232);
  not g2574 (n_1233, n1618);
  and g2575 (n1638, n_1233, n1636);
  not g2576 (n_1234, n1637);
  not g2577 (n_1235, n1638);
  and g2578 (n1639, n_1234, n_1235);
  and g2579 (n1640, n1617, n1639);
  not g2580 (n_1236, n1617);
  not g2581 (n_1237, n1639);
  and g2582 (n1641, n_1236, n_1237);
  not g2583 (n_1238, n1640);
  not g2584 (n_1239, n1641);
  and g2585 (n1642, n_1238, n_1239);
  not g2586 (n_1240, n1606);
  not g2587 (n_1241, n1642);
  and g2588 (n1643, n_1240, n_1241);
  and g2589 (n1644, n1606, n1642);
  not g2590 (n_1242, n1643);
  not g2591 (n_1243, n1644);
  and g2592 (n1645, n_1242, n_1243);
  not g2593 (n_1244, n1604);
  and g2594 (n1646, n_1244, n1645);
  not g2595 (n_1245, n1645);
  and g2596 (n1647, n1604, n_1245);
  not g2597 (n_1246, n1646);
  not g2598 (n_1247, n1647);
  and g2599 (n1648, n_1246, n_1247);
  not g2600 (n_1248, n1593);
  and g2601 (n1649, n_1248, n1648);
  not g2602 (n_1249, n1648);
  and g2603 (n1650, n1593, n_1249);
  not g2604 (n_1250, n1649);
  not g2605 (n_1251, n1650);
  and g2606 (n1651, n_1250, n_1251);
  and g2607 (n1652, \b[10] , n700);
  and g2608 (n1653, \b[8] , n767);
  and g2609 (n1654, \b[9] , n695);
  and g2615 (n1657, n703, n738);
  not g2618 (n_1256, n1658);
  and g2619 (n1659, \a[11] , n_1256);
  not g2620 (n_1257, n1659);
  and g2621 (n1660, \a[11] , n_1257);
  and g2622 (n1661, n_1256, n_1257);
  not g2623 (n_1258, n1660);
  not g2624 (n_1259, n1661);
  and g2625 (n1662, n_1258, n_1259);
  not g2626 (n_1260, n1662);
  and g2627 (n1663, n1651, n_1260);
  not g2628 (n_1261, n1663);
  and g2629 (n1664, n1651, n_1261);
  and g2630 (n1665, n_1260, n_1261);
  not g2631 (n_1262, n1664);
  not g2632 (n_1263, n1665);
  and g2633 (n1666, n_1262, n_1263);
  and g2634 (n1667, n_1143, n_1147);
  and g2635 (n1668, n1666, n1667);
  not g2636 (n_1264, n1666);
  not g2637 (n_1265, n1667);
  and g2638 (n1669, n_1264, n_1265);
  not g2639 (n_1266, n1668);
  not g2640 (n_1267, n1669);
  and g2641 (n1670, n_1266, n_1267);
  and g2642 (n1671, \b[13] , n511);
  and g2643 (n1672, \b[11] , n541);
  and g2644 (n1673, \b[12] , n506);
  and g2650 (n1676, n514, n1008);
  not g2653 (n_1272, n1677);
  and g2654 (n1678, \a[8] , n_1272);
  not g2655 (n_1273, n1678);
  and g2656 (n1679, \a[8] , n_1273);
  and g2657 (n1680, n_1272, n_1273);
  not g2658 (n_1274, n1679);
  not g2659 (n_1275, n1680);
  and g2660 (n1681, n_1274, n_1275);
  not g2661 (n_1276, n1670);
  and g2662 (n1682, n_1276, n1681);
  not g2663 (n_1277, n1681);
  and g2664 (n1683, n1670, n_1277);
  not g2665 (n_1278, n1682);
  not g2666 (n_1279, n1683);
  and g2667 (n1684, n_1278, n_1279);
  and g2668 (n1685, n_1152, n_1155);
  not g2669 (n_1280, n1685);
  and g2670 (n1686, n1684, n_1280);
  not g2671 (n_1281, n1684);
  and g2672 (n1687, n_1281, n1685);
  not g2673 (n_1282, n1686);
  not g2674 (n_1283, n1687);
  and g2675 (n1688, n_1282, n_1283);
  not g2676 (n_1284, n1591);
  and g2677 (n1689, n_1284, n1688);
  not g2678 (n_1285, n1689);
  and g2679 (n1690, n1688, n_1285);
  and g2680 (n1691, n_1284, n_1285);
  not g2681 (n_1286, n1690);
  not g2682 (n_1287, n1691);
  and g2683 (n1692, n_1286, n_1287);
  and g2684 (n1693, n_1159, n_1163);
  and g2685 (n1694, n1692, n1693);
  not g2686 (n_1288, n1692);
  not g2687 (n_1289, n1693);
  and g2688 (n1695, n_1288, n_1289);
  not g2689 (n_1290, n1694);
  not g2690 (n_1291, n1695);
  and g2691 (n1696, n_1290, n_1291);
  and g2692 (n1697, \b[19] , n266);
  and g2693 (n1698, \b[17] , n284);
  and g2694 (n1699, \b[18] , n261);
  and g2700 (n1702, n_1171, n_1174);
  not g2701 (n_1296, \b[19] );
  and g2702 (n1703, n_1169, n_1296);
  and g2703 (n1704, \b[18] , \b[19] );
  not g2704 (n_1297, n1703);
  not g2705 (n_1298, n1704);
  and g2706 (n1705, n_1297, n_1298);
  not g2707 (n_1299, n1702);
  and g2708 (n1706, n_1299, n1705);
  not g2709 (n_1300, n1705);
  and g2710 (n1707, n1702, n_1300);
  not g2711 (n_1301, n1706);
  not g2712 (n_1302, n1707);
  and g2713 (n1708, n_1301, n_1302);
  and g2714 (n1709, n269, n1708);
  not g2717 (n_1304, n1710);
  and g2718 (n1711, \a[2] , n_1304);
  not g2719 (n_1305, n1711);
  and g2720 (n1712, \a[2] , n_1305);
  and g2721 (n1713, n_1304, n_1305);
  not g2722 (n_1306, n1712);
  not g2723 (n_1307, n1713);
  and g2724 (n1714, n_1306, n_1307);
  not g2725 (n_1308, n1714);
  and g2726 (n1715, n1696, n_1308);
  not g2727 (n_1309, n1715);
  and g2728 (n1716, n1696, n_1309);
  and g2729 (n1717, n_1308, n_1309);
  not g2730 (n_1310, n1716);
  not g2731 (n_1311, n1717);
  and g2732 (n1718, n_1310, n_1311);
  and g2733 (n1719, n_1182, n_1187);
  not g2734 (n_1312, n1718);
  not g2735 (n_1313, n1719);
  and g2736 (n1720, n_1312, n_1313);
  and g2737 (n1721, n1718, n1719);
  not g2738 (n_1314, n1720);
  not g2739 (n_1315, n1721);
  and g2740 (\f[19] , n_1314, n_1315);
  and g2741 (n1723, n_1285, n_1291);
  and g2742 (n1724, \b[17] , n362);
  and g2743 (n1725, \b[15] , n403);
  and g2744 (n1726, \b[16] , n357);
  and g2750 (n1729, n365, n1356);
  not g2753 (n_1320, n1730);
  and g2754 (n1731, \a[5] , n_1320);
  not g2755 (n_1321, n1731);
  and g2756 (n1732, \a[5] , n_1321);
  and g2757 (n1733, n_1320, n_1321);
  not g2758 (n_1322, n1732);
  not g2759 (n_1323, n1733);
  and g2760 (n1734, n_1322, n_1323);
  and g2761 (n1735, \b[14] , n511);
  and g2762 (n1736, \b[12] , n541);
  and g2763 (n1737, \b[13] , n506);
  and g2769 (n1740, n514, n1034);
  not g2772 (n_1328, n1741);
  and g2773 (n1742, \a[8] , n_1328);
  not g2774 (n_1329, n1742);
  and g2775 (n1743, \a[8] , n_1329);
  and g2776 (n1744, n_1328, n_1329);
  not g2777 (n_1330, n1743);
  not g2778 (n_1331, n1744);
  and g2779 (n1745, n_1330, n_1331);
  and g2780 (n1746, n_1261, n_1267);
  and g2781 (n1747, \b[11] , n700);
  and g2782 (n1748, \b[9] , n767);
  and g2783 (n1749, \b[10] , n695);
  and g2789 (n1752, n703, n818);
  not g2792 (n_1336, n1753);
  and g2793 (n1754, \a[11] , n_1336);
  not g2794 (n_1337, n1754);
  and g2795 (n1755, \a[11] , n_1337);
  and g2796 (n1756, n_1336, n_1337);
  not g2797 (n_1338, n1755);
  not g2798 (n_1339, n1756);
  and g2799 (n1757, n_1338, n_1339);
  and g2800 (n1758, n_1246, n_1250);
  and g2801 (n1759, n_1236, n1639);
  not g2802 (n_1340, n1759);
  and g2803 (n1760, n_1242, n_1340);
  and g2804 (n1761, \b[2] , n1627);
  and g2805 (n1762, n1500, n_1226);
  and g2806 (n1763, n1621, n1762);
  and g2807 (n1764, \b[0] , n1763);
  and g2808 (n1765, \b[1] , n1622);
  and g2814 (n1768, n296, n1630);
  not g2817 (n_1345, n1769);
  and g2818 (n1770, \a[20] , n_1345);
  not g2819 (n_1346, n1770);
  and g2820 (n1771, \a[20] , n_1346);
  and g2821 (n1772, n_1345, n_1346);
  not g2822 (n_1347, n1771);
  not g2823 (n_1348, n1772);
  and g2824 (n1773, n_1347, n_1348);
  and g2825 (n1774, n_1234, n1773);
  not g2826 (n_1349, n1773);
  and g2827 (n1775, n1637, n_1349);
  not g2828 (n_1350, n1774);
  not g2829 (n_1351, n1775);
  and g2830 (n1776, n_1350, n_1351);
  and g2831 (n1777, \b[5] , n1302);
  and g2832 (n1778, \b[3] , n1391);
  and g2833 (n1779, \b[4] , n1297);
  and g2839 (n1782, n394, n1305);
  not g2842 (n_1356, n1783);
  and g2843 (n1784, \a[17] , n_1356);
  not g2844 (n_1357, n1784);
  and g2845 (n1785, \a[17] , n_1357);
  and g2846 (n1786, n_1356, n_1357);
  not g2847 (n_1358, n1785);
  not g2848 (n_1359, n1786);
  and g2849 (n1787, n_1358, n_1359);
  not g2850 (n_1360, n1787);
  and g2851 (n1788, n1776, n_1360);
  not g2852 (n_1361, n1776);
  and g2853 (n1789, n_1361, n1787);
  not g2854 (n_1362, n1760);
  not g2855 (n_1363, n1789);
  and g2856 (n1790, n_1362, n_1363);
  not g2857 (n_1364, n1788);
  and g2858 (n1791, n_1364, n1790);
  not g2859 (n_1365, n1791);
  and g2860 (n1792, n_1362, n_1365);
  and g2861 (n1793, n_1364, n_1365);
  and g2862 (n1794, n_1363, n1793);
  not g2863 (n_1366, n1792);
  not g2864 (n_1367, n1794);
  and g2865 (n1795, n_1366, n_1367);
  and g2866 (n1796, \b[8] , n951);
  and g2867 (n1797, \b[6] , n1056);
  and g2868 (n1798, \b[7] , n946);
  and g2874 (n1801, n585, n954);
  not g2877 (n_1372, n1802);
  and g2878 (n1803, \a[14] , n_1372);
  not g2879 (n_1373, n1803);
  and g2880 (n1804, \a[14] , n_1373);
  and g2881 (n1805, n_1372, n_1373);
  not g2882 (n_1374, n1804);
  not g2883 (n_1375, n1805);
  and g2884 (n1806, n_1374, n_1375);
  and g2885 (n1807, n1795, n1806);
  not g2886 (n_1376, n1795);
  not g2887 (n_1377, n1806);
  and g2888 (n1808, n_1376, n_1377);
  not g2889 (n_1378, n1807);
  not g2890 (n_1379, n1808);
  and g2891 (n1809, n_1378, n_1379);
  not g2892 (n_1380, n1758);
  and g2893 (n1810, n_1380, n1809);
  not g2894 (n_1381, n1809);
  and g2895 (n1811, n1758, n_1381);
  not g2896 (n_1382, n1810);
  not g2897 (n_1383, n1811);
  and g2898 (n1812, n_1382, n_1383);
  not g2899 (n_1384, n1812);
  and g2900 (n1813, n1757, n_1384);
  not g2901 (n_1385, n1757);
  and g2902 (n1814, n_1385, n1812);
  not g2903 (n_1386, n1813);
  not g2904 (n_1387, n1814);
  and g2905 (n1815, n_1386, n_1387);
  not g2906 (n_1388, n1746);
  and g2907 (n1816, n_1388, n1815);
  not g2908 (n_1389, n1815);
  and g2909 (n1817, n1746, n_1389);
  not g2910 (n_1390, n1816);
  not g2911 (n_1391, n1817);
  and g2912 (n1818, n_1390, n_1391);
  not g2913 (n_1392, n1745);
  and g2914 (n1819, n_1392, n1818);
  not g2915 (n_1393, n1819);
  and g2916 (n1820, n1818, n_1393);
  and g2917 (n1821, n_1392, n_1393);
  not g2918 (n_1394, n1820);
  not g2919 (n_1395, n1821);
  and g2920 (n1822, n_1394, n_1395);
  and g2921 (n1823, n_1279, n_1282);
  not g2922 (n_1396, n1822);
  not g2923 (n_1397, n1823);
  and g2924 (n1824, n_1396, n_1397);
  and g2925 (n1825, n1822, n1823);
  not g2926 (n_1398, n1824);
  not g2927 (n_1399, n1825);
  and g2928 (n1826, n_1398, n_1399);
  not g2929 (n_1400, n1734);
  and g2930 (n1827, n_1400, n1826);
  not g2931 (n_1401, n1827);
  and g2932 (n1828, n_1400, n_1401);
  and g2933 (n1829, n1826, n_1401);
  not g2934 (n_1402, n1828);
  not g2935 (n_1403, n1829);
  and g2936 (n1830, n_1402, n_1403);
  not g2937 (n_1404, n1723);
  not g2938 (n_1405, n1830);
  and g2939 (n1831, n_1404, n_1405);
  not g2940 (n_1406, n1831);
  and g2941 (n1832, n_1404, n_1406);
  and g2942 (n1833, n_1405, n_1406);
  not g2943 (n_1407, n1832);
  not g2944 (n_1408, n1833);
  and g2945 (n1834, n_1407, n_1408);
  and g2946 (n1835, \b[20] , n266);
  and g2947 (n1836, \b[18] , n284);
  and g2948 (n1837, \b[19] , n261);
  and g2954 (n1840, n_1298, n_1301);
  not g2955 (n_1413, \b[20] );
  and g2956 (n1841, n_1296, n_1413);
  and g2957 (n1842, \b[19] , \b[20] );
  not g2958 (n_1414, n1841);
  not g2959 (n_1415, n1842);
  and g2960 (n1843, n_1414, n_1415);
  not g2961 (n_1416, n1840);
  and g2962 (n1844, n_1416, n1843);
  not g2963 (n_1417, n1843);
  and g2964 (n1845, n1840, n_1417);
  not g2965 (n_1418, n1844);
  not g2966 (n_1419, n1845);
  and g2967 (n1846, n_1418, n_1419);
  and g2968 (n1847, n269, n1846);
  not g2971 (n_1421, n1848);
  and g2972 (n1849, \a[2] , n_1421);
  not g2973 (n_1422, n1849);
  and g2974 (n1850, \a[2] , n_1422);
  and g2975 (n1851, n_1421, n_1422);
  not g2976 (n_1423, n1850);
  not g2977 (n_1424, n1851);
  and g2978 (n1852, n_1423, n_1424);
  not g2979 (n_1425, n1834);
  not g2980 (n_1426, n1852);
  and g2981 (n1853, n_1425, n_1426);
  not g2982 (n_1427, n1853);
  and g2983 (n1854, n_1425, n_1427);
  and g2984 (n1855, n_1426, n_1427);
  not g2985 (n_1428, n1854);
  not g2986 (n_1429, n1855);
  and g2987 (n1856, n_1428, n_1429);
  and g2988 (n1857, n_1309, n_1314);
  not g2989 (n_1430, n1856);
  not g2990 (n_1431, n1857);
  and g2991 (n1858, n_1430, n_1431);
  and g2992 (n1859, n1856, n1857);
  not g2993 (n_1432, n1858);
  not g2994 (n_1433, n1859);
  and g2995 (\f[20] , n_1432, n_1433);
  and g2996 (n1861, n_1393, n_1398);
  and g2997 (n1862, \b[15] , n511);
  and g2998 (n1863, \b[13] , n541);
  and g2999 (n1864, \b[14] , n506);
  and g3005 (n1867, n514, n1131);
  not g3008 (n_1438, n1868);
  and g3009 (n1869, \a[8] , n_1438);
  not g3010 (n_1439, n1869);
  and g3011 (n1870, \a[8] , n_1439);
  and g3012 (n1871, n_1438, n_1439);
  not g3013 (n_1440, n1870);
  not g3014 (n_1441, n1871);
  and g3015 (n1872, n_1440, n_1441);
  and g3016 (n1873, n_1387, n_1390);
  and g3017 (n1874, \b[12] , n700);
  and g3018 (n1875, \b[10] , n767);
  and g3019 (n1876, \b[11] , n695);
  and g3025 (n1879, n703, n842);
  not g3028 (n_1446, n1880);
  and g3029 (n1881, \a[11] , n_1446);
  not g3030 (n_1447, n1881);
  and g3031 (n1882, \a[11] , n_1447);
  and g3032 (n1883, n_1446, n_1447);
  not g3033 (n_1448, n1882);
  not g3034 (n_1449, n1883);
  and g3035 (n1884, n_1448, n_1449);
  and g3036 (n1885, n_1379, n_1382);
  and g3037 (n1886, \b[6] , n1302);
  and g3038 (n1887, \b[4] , n1391);
  and g3039 (n1888, \b[5] , n1297);
  and g3045 (n1891, n459, n1305);
  not g3048 (n_1454, n1892);
  and g3049 (n1893, \a[17] , n_1454);
  not g3050 (n_1455, n1893);
  and g3051 (n1894, \a[17] , n_1455);
  and g3052 (n1895, n_1454, n_1455);
  not g3053 (n_1456, n1894);
  not g3054 (n_1457, n1895);
  and g3055 (n1896, n_1456, n_1457);
  not g3056 (n_1459, \a[21] );
  and g3057 (n1897, \a[20] , n_1459);
  and g3058 (n1898, n_1221, \a[21] );
  not g3059 (n_1460, n1897);
  not g3060 (n_1461, n1898);
  and g3061 (n1899, n_1460, n_1461);
  not g3062 (n_1462, n1899);
  and g3063 (n1900, \b[0] , n_1462);
  and g3064 (n1901, n_1351, n1900);
  not g3065 (n_1463, n1900);
  and g3066 (n1902, n1775, n_1463);
  not g3067 (n_1464, n1901);
  not g3068 (n_1465, n1902);
  and g3069 (n1903, n_1464, n_1465);
  and g3070 (n1904, \b[3] , n1627);
  and g3071 (n1905, \b[1] , n1763);
  and g3072 (n1906, \b[2] , n1622);
  and g3078 (n1909, n318, n1630);
  not g3081 (n_1470, n1910);
  and g3082 (n1911, \a[20] , n_1470);
  not g3083 (n_1471, n1911);
  and g3084 (n1912, \a[20] , n_1471);
  and g3085 (n1913, n_1470, n_1471);
  not g3086 (n_1472, n1912);
  not g3087 (n_1473, n1913);
  and g3088 (n1914, n_1472, n_1473);
  not g3089 (n_1474, n1903);
  not g3090 (n_1475, n1914);
  and g3091 (n1915, n_1474, n_1475);
  and g3092 (n1916, n1903, n1914);
  not g3093 (n_1476, n1915);
  not g3094 (n_1477, n1916);
  and g3095 (n1917, n_1476, n_1477);
  not g3096 (n_1478, n1896);
  and g3097 (n1918, n_1478, n1917);
  not g3098 (n_1479, n1918);
  and g3099 (n1919, n1917, n_1479);
  and g3100 (n1920, n_1478, n_1479);
  not g3101 (n_1480, n1919);
  not g3102 (n_1481, n1920);
  and g3103 (n1921, n_1480, n_1481);
  not g3104 (n_1482, n1793);
  and g3105 (n1922, n_1482, n1921);
  not g3106 (n_1483, n1921);
  and g3107 (n1923, n1793, n_1483);
  not g3108 (n_1484, n1922);
  not g3109 (n_1485, n1923);
  and g3110 (n1924, n_1484, n_1485);
  and g3111 (n1925, \b[9] , n951);
  and g3112 (n1926, \b[7] , n1056);
  and g3113 (n1927, \b[8] , n946);
  and g3119 (n1930, n651, n954);
  not g3122 (n_1490, n1931);
  and g3123 (n1932, \a[14] , n_1490);
  not g3124 (n_1491, n1932);
  and g3125 (n1933, \a[14] , n_1491);
  and g3126 (n1934, n_1490, n_1491);
  not g3127 (n_1492, n1933);
  not g3128 (n_1493, n1934);
  and g3129 (n1935, n_1492, n_1493);
  not g3130 (n_1494, n1924);
  not g3131 (n_1495, n1935);
  and g3132 (n1936, n_1494, n_1495);
  and g3133 (n1937, n1924, n1935);
  not g3134 (n_1496, n1936);
  not g3135 (n_1497, n1937);
  and g3136 (n1938, n_1496, n_1497);
  not g3137 (n_1498, n1885);
  and g3138 (n1939, n_1498, n1938);
  not g3139 (n_1499, n1938);
  and g3140 (n1940, n1885, n_1499);
  not g3141 (n_1500, n1939);
  not g3142 (n_1501, n1940);
  and g3143 (n1941, n_1500, n_1501);
  not g3144 (n_1502, n1941);
  and g3145 (n1942, n1884, n_1502);
  not g3146 (n_1503, n1884);
  and g3147 (n1943, n_1503, n1941);
  not g3148 (n_1504, n1942);
  not g3149 (n_1505, n1943);
  and g3150 (n1944, n_1504, n_1505);
  not g3151 (n_1506, n1873);
  and g3152 (n1945, n_1506, n1944);
  not g3153 (n_1507, n1944);
  and g3154 (n1946, n1873, n_1507);
  not g3155 (n_1508, n1945);
  not g3156 (n_1509, n1946);
  and g3157 (n1947, n_1508, n_1509);
  not g3158 (n_1510, n1872);
  and g3159 (n1948, n_1510, n1947);
  not g3160 (n_1511, n1947);
  and g3161 (n1949, n1872, n_1511);
  not g3162 (n_1512, n1948);
  not g3163 (n_1513, n1949);
  and g3164 (n1950, n_1512, n_1513);
  not g3165 (n_1514, n1861);
  and g3166 (n1951, n_1514, n1950);
  not g3167 (n_1515, n1950);
  and g3168 (n1952, n1861, n_1515);
  not g3169 (n_1516, n1951);
  not g3170 (n_1517, n1952);
  and g3171 (n1953, n_1516, n_1517);
  and g3172 (n1954, \b[18] , n362);
  and g3173 (n1955, \b[16] , n403);
  and g3174 (n1956, \b[17] , n357);
  and g3180 (n1959, n365, n1566);
  not g3183 (n_1522, n1960);
  and g3184 (n1961, \a[5] , n_1522);
  not g3185 (n_1523, n1961);
  and g3186 (n1962, \a[5] , n_1523);
  and g3187 (n1963, n_1522, n_1523);
  not g3188 (n_1524, n1962);
  not g3189 (n_1525, n1963);
  and g3190 (n1964, n_1524, n_1525);
  not g3191 (n_1526, n1964);
  and g3192 (n1965, n1953, n_1526);
  not g3193 (n_1527, n1965);
  and g3194 (n1966, n1953, n_1527);
  and g3195 (n1967, n_1526, n_1527);
  not g3196 (n_1528, n1966);
  not g3197 (n_1529, n1967);
  and g3198 (n1968, n_1528, n_1529);
  and g3199 (n1969, n_1401, n_1406);
  and g3200 (n1970, n1968, n1969);
  not g3201 (n_1530, n1968);
  not g3202 (n_1531, n1969);
  and g3203 (n1971, n_1530, n_1531);
  not g3204 (n_1532, n1970);
  not g3205 (n_1533, n1971);
  and g3206 (n1972, n_1532, n_1533);
  and g3207 (n1973, \b[21] , n266);
  and g3208 (n1974, \b[19] , n284);
  and g3209 (n1975, \b[20] , n261);
  and g3215 (n1978, n_1415, n_1418);
  not g3216 (n_1538, \b[21] );
  and g3217 (n1979, n_1413, n_1538);
  and g3218 (n1980, \b[20] , \b[21] );
  not g3219 (n_1539, n1979);
  not g3220 (n_1540, n1980);
  and g3221 (n1981, n_1539, n_1540);
  not g3222 (n_1541, n1978);
  and g3223 (n1982, n_1541, n1981);
  not g3224 (n_1542, n1981);
  and g3225 (n1983, n1978, n_1542);
  not g3226 (n_1543, n1982);
  not g3227 (n_1544, n1983);
  and g3228 (n1984, n_1543, n_1544);
  and g3229 (n1985, n269, n1984);
  not g3232 (n_1546, n1986);
  and g3233 (n1987, \a[2] , n_1546);
  not g3234 (n_1547, n1987);
  and g3235 (n1988, \a[2] , n_1547);
  and g3236 (n1989, n_1546, n_1547);
  not g3237 (n_1548, n1988);
  not g3238 (n_1549, n1989);
  and g3239 (n1990, n_1548, n_1549);
  not g3240 (n_1550, n1990);
  and g3241 (n1991, n1972, n_1550);
  not g3242 (n_1551, n1991);
  and g3243 (n1992, n1972, n_1551);
  and g3244 (n1993, n_1550, n_1551);
  not g3245 (n_1552, n1992);
  not g3246 (n_1553, n1993);
  and g3247 (n1994, n_1552, n_1553);
  and g3248 (n1995, n_1427, n_1432);
  not g3249 (n_1554, n1994);
  not g3250 (n_1555, n1995);
  and g3251 (n1996, n_1554, n_1555);
  and g3252 (n1997, n1994, n1995);
  not g3253 (n_1556, n1996);
  not g3254 (n_1557, n1997);
  and g3255 (\f[21] , n_1556, n_1557);
  and g3256 (n1999, n_1551, n_1556);
  and g3257 (n2000, n_1512, n_1516);
  and g3258 (n2001, \b[16] , n511);
  and g3259 (n2002, \b[14] , n541);
  and g3260 (n2003, \b[15] , n506);
  and g3266 (n2006, n514, n1237);
  not g3269 (n_1562, n2007);
  and g3270 (n2008, \a[8] , n_1562);
  not g3271 (n_1563, n2008);
  and g3272 (n2009, \a[8] , n_1563);
  and g3273 (n2010, n_1562, n_1563);
  not g3274 (n_1564, n2009);
  not g3275 (n_1565, n2010);
  and g3276 (n2011, n_1564, n_1565);
  and g3277 (n2012, n_1505, n_1508);
  and g3278 (n2013, n_1482, n_1483);
  not g3279 (n_1566, n2013);
  and g3280 (n2014, n_1479, n_1566);
  and g3281 (n2015, \b[7] , n1302);
  and g3282 (n2016, \b[5] , n1391);
  and g3283 (n2017, \b[6] , n1297);
  and g3289 (n2020, n484, n1305);
  not g3292 (n_1571, n2021);
  and g3293 (n2022, \a[17] , n_1571);
  not g3294 (n_1572, n2022);
  and g3295 (n2023, \a[17] , n_1572);
  and g3296 (n2024, n_1571, n_1572);
  not g3297 (n_1573, n2023);
  not g3298 (n_1574, n2024);
  and g3299 (n2025, n_1573, n_1574);
  and g3300 (n2026, n1775, n1900);
  not g3301 (n_1575, n2026);
  and g3302 (n2027, n_1476, n_1575);
  and g3303 (n2028, \b[4] , n1627);
  and g3304 (n2029, \b[2] , n1763);
  and g3305 (n2030, \b[3] , n1622);
  and g3311 (n2033, n346, n1630);
  not g3314 (n_1580, n2034);
  and g3315 (n2035, \a[20] , n_1580);
  not g3316 (n_1581, n2035);
  and g3317 (n2036, \a[20] , n_1581);
  and g3318 (n2037, n_1580, n_1581);
  not g3319 (n_1582, n2036);
  not g3320 (n_1583, n2037);
  and g3321 (n2038, n_1582, n_1583);
  and g3322 (n2039, \a[23] , n_1463);
  and g3323 (n2040, n_1459, \a[22] );
  not g3324 (n_1586, \a[22] );
  and g3325 (n2041, \a[21] , n_1586);
  not g3326 (n_1587, n2040);
  not g3327 (n_1588, n2041);
  and g3328 (n2042, n_1587, n_1588);
  not g3329 (n_1589, n2042);
  and g3330 (n2043, n1899, n_1589);
  and g3331 (n2044, \b[0] , n2043);
  and g3332 (n2045, n_1586, \a[23] );
  not g3333 (n_1590, \a[23] );
  and g3334 (n2046, \a[22] , n_1590);
  not g3335 (n_1591, n2045);
  not g3336 (n_1592, n2046);
  and g3337 (n2047, n_1591, n_1592);
  and g3338 (n2048, n_1462, n2047);
  and g3339 (n2049, \b[1] , n2048);
  not g3340 (n_1593, n2044);
  not g3341 (n_1594, n2049);
  and g3342 (n2050, n_1593, n_1594);
  not g3343 (n_1595, n2047);
  and g3344 (n2051, n_1462, n_1595);
  and g3345 (n2052, n_21, n2051);
  not g3346 (n_1596, n2052);
  and g3347 (n2053, n2050, n_1596);
  not g3348 (n_1597, n2053);
  and g3349 (n2054, \a[23] , n_1597);
  not g3350 (n_1598, n2054);
  and g3351 (n2055, \a[23] , n_1598);
  and g3352 (n2056, n_1597, n_1598);
  not g3353 (n_1599, n2055);
  not g3354 (n_1600, n2056);
  and g3355 (n2057, n_1599, n_1600);
  not g3356 (n_1601, n2057);
  and g3357 (n2058, n2039, n_1601);
  not g3358 (n_1602, n2039);
  and g3359 (n2059, n_1602, n2057);
  not g3360 (n_1603, n2058);
  not g3361 (n_1604, n2059);
  and g3362 (n2060, n_1603, n_1604);
  and g3363 (n2061, n2038, n2060);
  not g3364 (n_1605, n2038);
  not g3365 (n_1606, n2060);
  and g3366 (n2062, n_1605, n_1606);
  not g3367 (n_1607, n2061);
  not g3368 (n_1608, n2062);
  and g3369 (n2063, n_1607, n_1608);
  not g3370 (n_1609, n2027);
  not g3371 (n_1610, n2063);
  and g3372 (n2064, n_1609, n_1610);
  and g3373 (n2065, n2027, n2063);
  not g3374 (n_1611, n2064);
  not g3375 (n_1612, n2065);
  and g3376 (n2066, n_1611, n_1612);
  not g3377 (n_1613, n2025);
  and g3378 (n2067, n_1613, n2066);
  not g3379 (n_1614, n2066);
  and g3380 (n2068, n2025, n_1614);
  not g3381 (n_1615, n2067);
  not g3382 (n_1616, n2068);
  and g3383 (n2069, n_1615, n_1616);
  not g3384 (n_1617, n2014);
  and g3385 (n2070, n_1617, n2069);
  not g3386 (n_1618, n2069);
  and g3387 (n2071, n2014, n_1618);
  not g3388 (n_1619, n2070);
  not g3389 (n_1620, n2071);
  and g3390 (n2072, n_1619, n_1620);
  and g3391 (n2073, \b[10] , n951);
  and g3392 (n2074, \b[8] , n1056);
  and g3393 (n2075, \b[9] , n946);
  and g3399 (n2078, n738, n954);
  not g3402 (n_1625, n2079);
  and g3403 (n2080, \a[14] , n_1625);
  not g3404 (n_1626, n2080);
  and g3405 (n2081, \a[14] , n_1626);
  and g3406 (n2082, n_1625, n_1626);
  not g3407 (n_1627, n2081);
  not g3408 (n_1628, n2082);
  and g3409 (n2083, n_1627, n_1628);
  not g3410 (n_1629, n2083);
  and g3411 (n2084, n2072, n_1629);
  not g3412 (n_1630, n2084);
  and g3413 (n2085, n2072, n_1630);
  and g3414 (n2086, n_1629, n_1630);
  not g3415 (n_1631, n2085);
  not g3416 (n_1632, n2086);
  and g3417 (n2087, n_1631, n_1632);
  and g3418 (n2088, n_1496, n_1500);
  and g3419 (n2089, n2087, n2088);
  not g3420 (n_1633, n2087);
  not g3421 (n_1634, n2088);
  and g3422 (n2090, n_1633, n_1634);
  not g3423 (n_1635, n2089);
  not g3424 (n_1636, n2090);
  and g3425 (n2091, n_1635, n_1636);
  and g3426 (n2092, \b[13] , n700);
  and g3427 (n2093, \b[11] , n767);
  and g3428 (n2094, \b[12] , n695);
  and g3434 (n2097, n703, n1008);
  not g3437 (n_1641, n2098);
  and g3438 (n2099, \a[11] , n_1641);
  not g3439 (n_1642, n2099);
  and g3440 (n2100, \a[11] , n_1642);
  and g3441 (n2101, n_1641, n_1642);
  not g3442 (n_1643, n2100);
  not g3443 (n_1644, n2101);
  and g3444 (n2102, n_1643, n_1644);
  not g3445 (n_1645, n2091);
  and g3446 (n2103, n_1645, n2102);
  not g3447 (n_1646, n2102);
  and g3448 (n2104, n2091, n_1646);
  not g3449 (n_1647, n2103);
  not g3450 (n_1648, n2104);
  and g3451 (n2105, n_1647, n_1648);
  not g3452 (n_1649, n2012);
  and g3453 (n2106, n_1649, n2105);
  not g3454 (n_1650, n2105);
  and g3455 (n2107, n2012, n_1650);
  not g3456 (n_1651, n2106);
  not g3457 (n_1652, n2107);
  and g3458 (n2108, n_1651, n_1652);
  not g3459 (n_1653, n2011);
  and g3460 (n2109, n_1653, n2108);
  not g3461 (n_1654, n2108);
  and g3462 (n2110, n2011, n_1654);
  not g3463 (n_1655, n2109);
  not g3464 (n_1656, n2110);
  and g3465 (n2111, n_1655, n_1656);
  not g3466 (n_1657, n2000);
  and g3467 (n2112, n_1657, n2111);
  not g3468 (n_1658, n2111);
  and g3469 (n2113, n2000, n_1658);
  not g3470 (n_1659, n2112);
  not g3471 (n_1660, n2113);
  and g3472 (n2114, n_1659, n_1660);
  and g3473 (n2115, \b[19] , n362);
  and g3474 (n2116, \b[17] , n403);
  and g3475 (n2117, \b[18] , n357);
  and g3481 (n2120, n365, n1708);
  not g3484 (n_1665, n2121);
  and g3485 (n2122, \a[5] , n_1665);
  not g3486 (n_1666, n2122);
  and g3487 (n2123, \a[5] , n_1666);
  and g3488 (n2124, n_1665, n_1666);
  not g3489 (n_1667, n2123);
  not g3490 (n_1668, n2124);
  and g3491 (n2125, n_1667, n_1668);
  not g3492 (n_1669, n2125);
  and g3493 (n2126, n2114, n_1669);
  not g3494 (n_1670, n2126);
  and g3495 (n2127, n2114, n_1670);
  and g3496 (n2128, n_1669, n_1670);
  not g3497 (n_1671, n2127);
  not g3498 (n_1672, n2128);
  and g3499 (n2129, n_1671, n_1672);
  and g3500 (n2130, n_1527, n_1533);
  and g3501 (n2131, n2129, n2130);
  not g3502 (n_1673, n2129);
  not g3503 (n_1674, n2130);
  and g3504 (n2132, n_1673, n_1674);
  not g3505 (n_1675, n2131);
  not g3506 (n_1676, n2132);
  and g3507 (n2133, n_1675, n_1676);
  and g3508 (n2134, \b[22] , n266);
  and g3509 (n2135, \b[20] , n284);
  and g3510 (n2136, \b[21] , n261);
  and g3516 (n2139, n_1540, n_1543);
  not g3517 (n_1681, \b[22] );
  and g3518 (n2140, n_1538, n_1681);
  and g3519 (n2141, \b[21] , \b[22] );
  not g3520 (n_1682, n2140);
  not g3521 (n_1683, n2141);
  and g3522 (n2142, n_1682, n_1683);
  not g3523 (n_1684, n2139);
  and g3524 (n2143, n_1684, n2142);
  not g3525 (n_1685, n2142);
  and g3526 (n2144, n2139, n_1685);
  not g3527 (n_1686, n2143);
  not g3528 (n_1687, n2144);
  and g3529 (n2145, n_1686, n_1687);
  and g3530 (n2146, n269, n2145);
  not g3533 (n_1689, n2147);
  and g3534 (n2148, \a[2] , n_1689);
  not g3535 (n_1690, n2148);
  and g3536 (n2149, \a[2] , n_1690);
  and g3537 (n2150, n_1689, n_1690);
  not g3538 (n_1691, n2149);
  not g3539 (n_1692, n2150);
  and g3540 (n2151, n_1691, n_1692);
  not g3541 (n_1693, n2133);
  and g3542 (n2152, n_1693, n2151);
  not g3543 (n_1694, n2151);
  and g3544 (n2153, n2133, n_1694);
  not g3545 (n_1695, n2152);
  not g3546 (n_1696, n2153);
  and g3547 (n2154, n_1695, n_1696);
  not g3548 (n_1697, n1999);
  and g3549 (n2155, n_1697, n2154);
  not g3550 (n_1698, n2154);
  and g3551 (n2156, n1999, n_1698);
  not g3552 (n_1699, n2155);
  not g3553 (n_1700, n2156);
  and g3554 (\f[22] , n_1699, n_1700);
  and g3555 (n2158, n_1655, n_1659);
  and g3556 (n2159, \b[17] , n511);
  and g3557 (n2160, \b[15] , n541);
  and g3558 (n2161, \b[16] , n506);
  and g3564 (n2164, n514, n1356);
  not g3567 (n_1705, n2165);
  and g3568 (n2166, \a[8] , n_1705);
  not g3569 (n_1706, n2166);
  and g3570 (n2167, \a[8] , n_1706);
  and g3571 (n2168, n_1705, n_1706);
  not g3572 (n_1707, n2167);
  not g3573 (n_1708, n2168);
  and g3574 (n2169, n_1707, n_1708);
  and g3575 (n2170, \b[14] , n700);
  and g3576 (n2171, \b[12] , n767);
  and g3577 (n2172, \b[13] , n695);
  and g3583 (n2175, n703, n1034);
  not g3586 (n_1713, n2176);
  and g3587 (n2177, \a[11] , n_1713);
  not g3588 (n_1714, n2177);
  and g3589 (n2178, \a[11] , n_1714);
  and g3590 (n2179, n_1713, n_1714);
  not g3591 (n_1715, n2178);
  not g3592 (n_1716, n2179);
  and g3593 (n2180, n_1715, n_1716);
  and g3594 (n2181, n_1630, n_1636);
  and g3595 (n2182, \b[11] , n951);
  and g3596 (n2183, \b[9] , n1056);
  and g3597 (n2184, \b[10] , n946);
  and g3603 (n2187, n818, n954);
  not g3606 (n_1721, n2188);
  and g3607 (n2189, \a[14] , n_1721);
  not g3608 (n_1722, n2189);
  and g3609 (n2190, \a[14] , n_1722);
  and g3610 (n2191, n_1721, n_1722);
  not g3611 (n_1723, n2190);
  not g3612 (n_1724, n2191);
  and g3613 (n2192, n_1723, n_1724);
  and g3614 (n2193, n_1615, n_1619);
  and g3615 (n2194, n_1605, n2060);
  not g3616 (n_1725, n2194);
  and g3617 (n2195, n_1611, n_1725);
  and g3618 (n2196, \b[2] , n2048);
  and g3619 (n2197, n1899, n_1595);
  and g3620 (n2198, n2042, n2197);
  and g3621 (n2199, \b[0] , n2198);
  and g3622 (n2200, \b[1] , n2043);
  and g3628 (n2203, n296, n2051);
  not g3631 (n_1730, n2204);
  and g3632 (n2205, \a[23] , n_1730);
  not g3633 (n_1731, n2205);
  and g3634 (n2206, \a[23] , n_1731);
  and g3635 (n2207, n_1730, n_1731);
  not g3636 (n_1732, n2206);
  not g3637 (n_1733, n2207);
  and g3638 (n2208, n_1732, n_1733);
  and g3639 (n2209, n_1603, n2208);
  not g3640 (n_1734, n2208);
  and g3641 (n2210, n2058, n_1734);
  not g3642 (n_1735, n2209);
  not g3643 (n_1736, n2210);
  and g3644 (n2211, n_1735, n_1736);
  and g3645 (n2212, \b[5] , n1627);
  and g3646 (n2213, \b[3] , n1763);
  and g3647 (n2214, \b[4] , n1622);
  and g3653 (n2217, n394, n1630);
  not g3656 (n_1741, n2218);
  and g3657 (n2219, \a[20] , n_1741);
  not g3658 (n_1742, n2219);
  and g3659 (n2220, \a[20] , n_1742);
  and g3660 (n2221, n_1741, n_1742);
  not g3661 (n_1743, n2220);
  not g3662 (n_1744, n2221);
  and g3663 (n2222, n_1743, n_1744);
  not g3664 (n_1745, n2222);
  and g3665 (n2223, n2211, n_1745);
  not g3666 (n_1746, n2211);
  and g3667 (n2224, n_1746, n2222);
  not g3668 (n_1747, n2195);
  not g3669 (n_1748, n2224);
  and g3670 (n2225, n_1747, n_1748);
  not g3671 (n_1749, n2223);
  and g3672 (n2226, n_1749, n2225);
  not g3673 (n_1750, n2226);
  and g3674 (n2227, n_1747, n_1750);
  and g3675 (n2228, n_1749, n_1750);
  and g3676 (n2229, n_1748, n2228);
  not g3677 (n_1751, n2227);
  not g3678 (n_1752, n2229);
  and g3679 (n2230, n_1751, n_1752);
  and g3680 (n2231, \b[8] , n1302);
  and g3681 (n2232, \b[6] , n1391);
  and g3682 (n2233, \b[7] , n1297);
  and g3688 (n2236, n585, n1305);
  not g3691 (n_1757, n2237);
  and g3692 (n2238, \a[17] , n_1757);
  not g3693 (n_1758, n2238);
  and g3694 (n2239, \a[17] , n_1758);
  and g3695 (n2240, n_1757, n_1758);
  not g3696 (n_1759, n2239);
  not g3697 (n_1760, n2240);
  and g3698 (n2241, n_1759, n_1760);
  and g3699 (n2242, n2230, n2241);
  not g3700 (n_1761, n2230);
  not g3701 (n_1762, n2241);
  and g3702 (n2243, n_1761, n_1762);
  not g3703 (n_1763, n2242);
  not g3704 (n_1764, n2243);
  and g3705 (n2244, n_1763, n_1764);
  not g3706 (n_1765, n2193);
  and g3707 (n2245, n_1765, n2244);
  not g3708 (n_1766, n2244);
  and g3709 (n2246, n2193, n_1766);
  not g3710 (n_1767, n2245);
  not g3711 (n_1768, n2246);
  and g3712 (n2247, n_1767, n_1768);
  not g3713 (n_1769, n2247);
  and g3714 (n2248, n2192, n_1769);
  not g3715 (n_1770, n2192);
  and g3716 (n2249, n_1770, n2247);
  not g3717 (n_1771, n2248);
  not g3718 (n_1772, n2249);
  and g3719 (n2250, n_1771, n_1772);
  not g3720 (n_1773, n2181);
  and g3721 (n2251, n_1773, n2250);
  not g3722 (n_1774, n2250);
  and g3723 (n2252, n2181, n_1774);
  not g3724 (n_1775, n2251);
  not g3725 (n_1776, n2252);
  and g3726 (n2253, n_1775, n_1776);
  not g3727 (n_1777, n2180);
  and g3728 (n2254, n_1777, n2253);
  not g3729 (n_1778, n2254);
  and g3730 (n2255, n2253, n_1778);
  and g3731 (n2256, n_1777, n_1778);
  not g3732 (n_1779, n2255);
  not g3733 (n_1780, n2256);
  and g3734 (n2257, n_1779, n_1780);
  and g3735 (n2258, n_1648, n_1651);
  not g3736 (n_1781, n2257);
  not g3737 (n_1782, n2258);
  and g3738 (n2259, n_1781, n_1782);
  and g3739 (n2260, n2257, n2258);
  not g3740 (n_1783, n2259);
  not g3741 (n_1784, n2260);
  and g3742 (n2261, n_1783, n_1784);
  not g3743 (n_1785, n2169);
  and g3744 (n2262, n_1785, n2261);
  not g3745 (n_1786, n2262);
  and g3746 (n2263, n_1785, n_1786);
  and g3747 (n2264, n2261, n_1786);
  not g3748 (n_1787, n2263);
  not g3749 (n_1788, n2264);
  and g3750 (n2265, n_1787, n_1788);
  not g3751 (n_1789, n2158);
  not g3752 (n_1790, n2265);
  and g3753 (n2266, n_1789, n_1790);
  not g3754 (n_1791, n2266);
  and g3755 (n2267, n_1789, n_1791);
  and g3756 (n2268, n_1790, n_1791);
  not g3757 (n_1792, n2267);
  not g3758 (n_1793, n2268);
  and g3759 (n2269, n_1792, n_1793);
  and g3760 (n2270, \b[20] , n362);
  and g3761 (n2271, \b[18] , n403);
  and g3762 (n2272, \b[19] , n357);
  and g3768 (n2275, n365, n1846);
  not g3771 (n_1798, n2276);
  and g3772 (n2277, \a[5] , n_1798);
  not g3773 (n_1799, n2277);
  and g3774 (n2278, \a[5] , n_1799);
  and g3775 (n2279, n_1798, n_1799);
  not g3776 (n_1800, n2278);
  not g3777 (n_1801, n2279);
  and g3778 (n2280, n_1800, n_1801);
  not g3779 (n_1802, n2269);
  not g3780 (n_1803, n2280);
  and g3781 (n2281, n_1802, n_1803);
  not g3782 (n_1804, n2281);
  and g3783 (n2282, n_1802, n_1804);
  and g3784 (n2283, n_1803, n_1804);
  not g3785 (n_1805, n2282);
  not g3786 (n_1806, n2283);
  and g3787 (n2284, n_1805, n_1806);
  and g3788 (n2285, n_1670, n_1676);
  and g3789 (n2286, n2284, n2285);
  not g3790 (n_1807, n2284);
  not g3791 (n_1808, n2285);
  and g3792 (n2287, n_1807, n_1808);
  not g3793 (n_1809, n2286);
  not g3794 (n_1810, n2287);
  and g3795 (n2288, n_1809, n_1810);
  and g3796 (n2289, \b[23] , n266);
  and g3797 (n2290, \b[21] , n284);
  and g3798 (n2291, \b[22] , n261);
  and g3804 (n2294, n_1683, n_1686);
  not g3805 (n_1815, \b[23] );
  and g3806 (n2295, n_1681, n_1815);
  and g3807 (n2296, \b[22] , \b[23] );
  not g3808 (n_1816, n2295);
  not g3809 (n_1817, n2296);
  and g3810 (n2297, n_1816, n_1817);
  not g3811 (n_1818, n2294);
  and g3812 (n2298, n_1818, n2297);
  not g3813 (n_1819, n2297);
  and g3814 (n2299, n2294, n_1819);
  not g3815 (n_1820, n2298);
  not g3816 (n_1821, n2299);
  and g3817 (n2300, n_1820, n_1821);
  and g3818 (n2301, n269, n2300);
  not g3821 (n_1823, n2302);
  and g3822 (n2303, \a[2] , n_1823);
  not g3823 (n_1824, n2303);
  and g3824 (n2304, \a[2] , n_1824);
  and g3825 (n2305, n_1823, n_1824);
  not g3826 (n_1825, n2304);
  not g3827 (n_1826, n2305);
  and g3828 (n2306, n_1825, n_1826);
  not g3829 (n_1827, n2306);
  and g3830 (n2307, n2288, n_1827);
  not g3831 (n_1828, n2307);
  and g3832 (n2308, n2288, n_1828);
  and g3833 (n2309, n_1827, n_1828);
  not g3834 (n_1829, n2308);
  not g3835 (n_1830, n2309);
  and g3836 (n2310, n_1829, n_1830);
  and g3837 (n2311, n_1696, n_1699);
  not g3838 (n_1831, n2310);
  not g3839 (n_1832, n2311);
  and g3840 (n2312, n_1831, n_1832);
  and g3841 (n2313, n2310, n2311);
  not g3842 (n_1833, n2312);
  not g3843 (n_1834, n2313);
  and g3844 (\f[23] , n_1833, n_1834);
  and g3845 (n2315, n_1804, n_1810);
  and g3846 (n2316, \b[21] , n362);
  and g3847 (n2317, \b[19] , n403);
  and g3848 (n2318, \b[20] , n357);
  and g3854 (n2321, n365, n1984);
  not g3857 (n_1839, n2322);
  and g3858 (n2323, \a[5] , n_1839);
  not g3859 (n_1840, n2323);
  and g3860 (n2324, \a[5] , n_1840);
  and g3861 (n2325, n_1839, n_1840);
  not g3862 (n_1841, n2324);
  not g3863 (n_1842, n2325);
  and g3864 (n2326, n_1841, n_1842);
  and g3865 (n2327, n_1786, n_1791);
  and g3866 (n2328, \b[15] , n700);
  and g3867 (n2329, \b[13] , n767);
  and g3868 (n2330, \b[14] , n695);
  and g3874 (n2333, n703, n1131);
  not g3877 (n_1847, n2334);
  and g3878 (n2335, \a[11] , n_1847);
  not g3879 (n_1848, n2335);
  and g3880 (n2336, \a[11] , n_1848);
  and g3881 (n2337, n_1847, n_1848);
  not g3882 (n_1849, n2336);
  not g3883 (n_1850, n2337);
  and g3884 (n2338, n_1849, n_1850);
  and g3885 (n2339, n_1772, n_1775);
  and g3886 (n2340, \b[12] , n951);
  and g3887 (n2341, \b[10] , n1056);
  and g3888 (n2342, \b[11] , n946);
  and g3894 (n2345, n842, n954);
  not g3897 (n_1855, n2346);
  and g3898 (n2347, \a[14] , n_1855);
  not g3899 (n_1856, n2347);
  and g3900 (n2348, \a[14] , n_1856);
  and g3901 (n2349, n_1855, n_1856);
  not g3902 (n_1857, n2348);
  not g3903 (n_1858, n2349);
  and g3904 (n2350, n_1857, n_1858);
  and g3905 (n2351, n_1764, n_1767);
  and g3906 (n2352, \b[6] , n1627);
  and g3907 (n2353, \b[4] , n1763);
  and g3908 (n2354, \b[5] , n1622);
  and g3914 (n2357, n459, n1630);
  not g3917 (n_1863, n2358);
  and g3918 (n2359, \a[20] , n_1863);
  not g3919 (n_1864, n2359);
  and g3920 (n2360, \a[20] , n_1864);
  and g3921 (n2361, n_1863, n_1864);
  not g3922 (n_1865, n2360);
  not g3923 (n_1866, n2361);
  and g3924 (n2362, n_1865, n_1866);
  not g3925 (n_1868, \a[24] );
  and g3926 (n2363, \a[23] , n_1868);
  and g3927 (n2364, n_1590, \a[24] );
  not g3928 (n_1869, n2363);
  not g3929 (n_1870, n2364);
  and g3930 (n2365, n_1869, n_1870);
  not g3931 (n_1871, n2365);
  and g3932 (n2366, \b[0] , n_1871);
  and g3933 (n2367, n_1736, n2366);
  not g3934 (n_1872, n2366);
  and g3935 (n2368, n2210, n_1872);
  not g3936 (n_1873, n2367);
  not g3937 (n_1874, n2368);
  and g3938 (n2369, n_1873, n_1874);
  and g3939 (n2370, \b[3] , n2048);
  and g3940 (n2371, \b[1] , n2198);
  and g3941 (n2372, \b[2] , n2043);
  and g3947 (n2375, n318, n2051);
  not g3950 (n_1879, n2376);
  and g3951 (n2377, \a[23] , n_1879);
  not g3952 (n_1880, n2377);
  and g3953 (n2378, \a[23] , n_1880);
  and g3954 (n2379, n_1879, n_1880);
  not g3955 (n_1881, n2378);
  not g3956 (n_1882, n2379);
  and g3957 (n2380, n_1881, n_1882);
  not g3958 (n_1883, n2369);
  not g3959 (n_1884, n2380);
  and g3960 (n2381, n_1883, n_1884);
  and g3961 (n2382, n2369, n2380);
  not g3962 (n_1885, n2381);
  not g3963 (n_1886, n2382);
  and g3964 (n2383, n_1885, n_1886);
  not g3965 (n_1887, n2362);
  and g3966 (n2384, n_1887, n2383);
  not g3967 (n_1888, n2384);
  and g3968 (n2385, n2383, n_1888);
  and g3969 (n2386, n_1887, n_1888);
  not g3970 (n_1889, n2385);
  not g3971 (n_1890, n2386);
  and g3972 (n2387, n_1889, n_1890);
  not g3973 (n_1891, n2228);
  and g3974 (n2388, n_1891, n2387);
  not g3975 (n_1892, n2387);
  and g3976 (n2389, n2228, n_1892);
  not g3977 (n_1893, n2388);
  not g3978 (n_1894, n2389);
  and g3979 (n2390, n_1893, n_1894);
  and g3980 (n2391, \b[9] , n1302);
  and g3981 (n2392, \b[7] , n1391);
  and g3982 (n2393, \b[8] , n1297);
  and g3988 (n2396, n651, n1305);
  not g3991 (n_1899, n2397);
  and g3992 (n2398, \a[17] , n_1899);
  not g3993 (n_1900, n2398);
  and g3994 (n2399, \a[17] , n_1900);
  and g3995 (n2400, n_1899, n_1900);
  not g3996 (n_1901, n2399);
  not g3997 (n_1902, n2400);
  and g3998 (n2401, n_1901, n_1902);
  not g3999 (n_1903, n2390);
  not g4000 (n_1904, n2401);
  and g4001 (n2402, n_1903, n_1904);
  and g4002 (n2403, n2390, n2401);
  not g4003 (n_1905, n2402);
  not g4004 (n_1906, n2403);
  and g4005 (n2404, n_1905, n_1906);
  not g4006 (n_1907, n2351);
  and g4007 (n2405, n_1907, n2404);
  not g4008 (n_1908, n2404);
  and g4009 (n2406, n2351, n_1908);
  not g4010 (n_1909, n2405);
  not g4011 (n_1910, n2406);
  and g4012 (n2407, n_1909, n_1910);
  not g4013 (n_1911, n2407);
  and g4014 (n2408, n2350, n_1911);
  not g4015 (n_1912, n2350);
  and g4016 (n2409, n_1912, n2407);
  not g4017 (n_1913, n2408);
  not g4018 (n_1914, n2409);
  and g4019 (n2410, n_1913, n_1914);
  not g4020 (n_1915, n2339);
  and g4021 (n2411, n_1915, n2410);
  not g4022 (n_1916, n2410);
  and g4023 (n2412, n2339, n_1916);
  not g4024 (n_1917, n2411);
  not g4025 (n_1918, n2412);
  and g4026 (n2413, n_1917, n_1918);
  not g4027 (n_1919, n2338);
  and g4028 (n2414, n_1919, n2413);
  not g4029 (n_1920, n2414);
  and g4030 (n2415, n2413, n_1920);
  and g4031 (n2416, n_1919, n_1920);
  not g4032 (n_1921, n2415);
  not g4033 (n_1922, n2416);
  and g4034 (n2417, n_1921, n_1922);
  and g4035 (n2418, n_1778, n_1783);
  and g4036 (n2419, n2417, n2418);
  not g4037 (n_1923, n2417);
  not g4038 (n_1924, n2418);
  and g4039 (n2420, n_1923, n_1924);
  not g4040 (n_1925, n2419);
  not g4041 (n_1926, n2420);
  and g4042 (n2421, n_1925, n_1926);
  and g4043 (n2422, \b[18] , n511);
  and g4044 (n2423, \b[16] , n541);
  and g4045 (n2424, \b[17] , n506);
  and g4051 (n2427, n514, n1566);
  not g4054 (n_1931, n2428);
  and g4055 (n2429, \a[8] , n_1931);
  not g4056 (n_1932, n2429);
  and g4057 (n2430, \a[8] , n_1932);
  and g4058 (n2431, n_1931, n_1932);
  not g4059 (n_1933, n2430);
  not g4060 (n_1934, n2431);
  and g4061 (n2432, n_1933, n_1934);
  not g4062 (n_1935, n2421);
  and g4063 (n2433, n_1935, n2432);
  not g4064 (n_1936, n2432);
  and g4065 (n2434, n2421, n_1936);
  not g4066 (n_1937, n2433);
  not g4067 (n_1938, n2434);
  and g4068 (n2435, n_1937, n_1938);
  not g4069 (n_1939, n2327);
  and g4070 (n2436, n_1939, n2435);
  not g4071 (n_1940, n2435);
  and g4072 (n2437, n2327, n_1940);
  not g4073 (n_1941, n2436);
  not g4074 (n_1942, n2437);
  and g4075 (n2438, n_1941, n_1942);
  not g4076 (n_1943, n2326);
  and g4077 (n2439, n_1943, n2438);
  not g4078 (n_1944, n2439);
  and g4079 (n2440, n_1943, n_1944);
  and g4080 (n2441, n2438, n_1944);
  not g4081 (n_1945, n2440);
  not g4082 (n_1946, n2441);
  and g4083 (n2442, n_1945, n_1946);
  not g4084 (n_1947, n2315);
  not g4085 (n_1948, n2442);
  and g4086 (n2443, n_1947, n_1948);
  not g4087 (n_1949, n2443);
  and g4088 (n2444, n_1947, n_1949);
  and g4089 (n2445, n_1948, n_1949);
  not g4090 (n_1950, n2444);
  not g4091 (n_1951, n2445);
  and g4092 (n2446, n_1950, n_1951);
  and g4093 (n2447, \b[24] , n266);
  and g4094 (n2448, \b[22] , n284);
  and g4095 (n2449, \b[23] , n261);
  and g4101 (n2452, n_1817, n_1820);
  not g4102 (n_1956, \b[24] );
  and g4103 (n2453, n_1815, n_1956);
  and g4104 (n2454, \b[23] , \b[24] );
  not g4105 (n_1957, n2453);
  not g4106 (n_1958, n2454);
  and g4107 (n2455, n_1957, n_1958);
  not g4108 (n_1959, n2452);
  and g4109 (n2456, n_1959, n2455);
  not g4110 (n_1960, n2455);
  and g4111 (n2457, n2452, n_1960);
  not g4112 (n_1961, n2456);
  not g4113 (n_1962, n2457);
  and g4114 (n2458, n_1961, n_1962);
  and g4115 (n2459, n269, n2458);
  not g4118 (n_1964, n2460);
  and g4119 (n2461, \a[2] , n_1964);
  not g4120 (n_1965, n2461);
  and g4121 (n2462, \a[2] , n_1965);
  and g4122 (n2463, n_1964, n_1965);
  not g4123 (n_1966, n2462);
  not g4124 (n_1967, n2463);
  and g4125 (n2464, n_1966, n_1967);
  not g4126 (n_1968, n2446);
  not g4127 (n_1969, n2464);
  and g4128 (n2465, n_1968, n_1969);
  not g4129 (n_1970, n2465);
  and g4130 (n2466, n_1968, n_1970);
  and g4131 (n2467, n_1969, n_1970);
  not g4132 (n_1971, n2466);
  not g4133 (n_1972, n2467);
  and g4134 (n2468, n_1971, n_1972);
  and g4135 (n2469, n_1828, n_1833);
  not g4136 (n_1973, n2468);
  not g4137 (n_1974, n2469);
  and g4138 (n2470, n_1973, n_1974);
  and g4139 (n2471, n2468, n2469);
  not g4140 (n_1975, n2470);
  not g4141 (n_1976, n2471);
  and g4142 (\f[24] , n_1975, n_1976);
  and g4143 (n2473, n_1970, n_1975);
  and g4144 (n2474, \b[25] , n266);
  and g4145 (n2475, \b[23] , n284);
  and g4146 (n2476, \b[24] , n261);
  and g4152 (n2479, n_1958, n_1961);
  not g4153 (n_1981, \b[25] );
  and g4154 (n2480, n_1956, n_1981);
  and g4155 (n2481, \b[24] , \b[25] );
  not g4156 (n_1982, n2480);
  not g4157 (n_1983, n2481);
  and g4158 (n2482, n_1982, n_1983);
  not g4159 (n_1984, n2479);
  and g4160 (n2483, n_1984, n2482);
  not g4161 (n_1985, n2482);
  and g4162 (n2484, n2479, n_1985);
  not g4163 (n_1986, n2483);
  not g4164 (n_1987, n2484);
  and g4165 (n2485, n_1986, n_1987);
  and g4166 (n2486, n269, n2485);
  not g4169 (n_1989, n2487);
  and g4170 (n2488, \a[2] , n_1989);
  not g4171 (n_1990, n2488);
  and g4172 (n2489, \a[2] , n_1990);
  and g4173 (n2490, n_1989, n_1990);
  not g4174 (n_1991, n2489);
  not g4175 (n_1992, n2490);
  and g4176 (n2491, n_1991, n_1992);
  and g4177 (n2492, n_1944, n_1949);
  and g4178 (n2493, \b[16] , n700);
  and g4179 (n2494, \b[14] , n767);
  and g4180 (n2495, \b[15] , n695);
  and g4186 (n2498, n703, n1237);
  not g4189 (n_1997, n2499);
  and g4190 (n2500, \a[11] , n_1997);
  not g4191 (n_1998, n2500);
  and g4192 (n2501, \a[11] , n_1998);
  and g4193 (n2502, n_1997, n_1998);
  not g4194 (n_1999, n2501);
  not g4195 (n_2000, n2502);
  and g4196 (n2503, n_1999, n_2000);
  and g4197 (n2504, n_1891, n_1892);
  not g4198 (n_2001, n2504);
  and g4199 (n2505, n_1888, n_2001);
  and g4200 (n2506, \b[7] , n1627);
  and g4201 (n2507, \b[5] , n1763);
  and g4202 (n2508, \b[6] , n1622);
  and g4208 (n2511, n484, n1630);
  not g4211 (n_2006, n2512);
  and g4212 (n2513, \a[20] , n_2006);
  not g4213 (n_2007, n2513);
  and g4214 (n2514, \a[20] , n_2007);
  and g4215 (n2515, n_2006, n_2007);
  not g4216 (n_2008, n2514);
  not g4217 (n_2009, n2515);
  and g4218 (n2516, n_2008, n_2009);
  and g4219 (n2517, n2210, n2366);
  not g4220 (n_2010, n2517);
  and g4221 (n2518, n_1885, n_2010);
  and g4222 (n2519, \b[4] , n2048);
  and g4223 (n2520, \b[2] , n2198);
  and g4224 (n2521, \b[3] , n2043);
  and g4230 (n2524, n346, n2051);
  not g4233 (n_2015, n2525);
  and g4234 (n2526, \a[23] , n_2015);
  not g4235 (n_2016, n2526);
  and g4236 (n2527, \a[23] , n_2016);
  and g4237 (n2528, n_2015, n_2016);
  not g4238 (n_2017, n2527);
  not g4239 (n_2018, n2528);
  and g4240 (n2529, n_2017, n_2018);
  and g4241 (n2530, \a[26] , n_1872);
  and g4242 (n2531, n_1868, \a[25] );
  not g4243 (n_2021, \a[25] );
  and g4244 (n2532, \a[24] , n_2021);
  not g4245 (n_2022, n2531);
  not g4246 (n_2023, n2532);
  and g4247 (n2533, n_2022, n_2023);
  not g4248 (n_2024, n2533);
  and g4249 (n2534, n2365, n_2024);
  and g4250 (n2535, \b[0] , n2534);
  and g4251 (n2536, n_2021, \a[26] );
  not g4252 (n_2025, \a[26] );
  and g4253 (n2537, \a[25] , n_2025);
  not g4254 (n_2026, n2536);
  not g4255 (n_2027, n2537);
  and g4256 (n2538, n_2026, n_2027);
  and g4257 (n2539, n_1871, n2538);
  and g4258 (n2540, \b[1] , n2539);
  not g4259 (n_2028, n2535);
  not g4260 (n_2029, n2540);
  and g4261 (n2541, n_2028, n_2029);
  not g4262 (n_2030, n2538);
  and g4263 (n2542, n_1871, n_2030);
  and g4264 (n2543, n_21, n2542);
  not g4265 (n_2031, n2543);
  and g4266 (n2544, n2541, n_2031);
  not g4267 (n_2032, n2544);
  and g4268 (n2545, \a[26] , n_2032);
  not g4269 (n_2033, n2545);
  and g4270 (n2546, \a[26] , n_2033);
  and g4271 (n2547, n_2032, n_2033);
  not g4272 (n_2034, n2546);
  not g4273 (n_2035, n2547);
  and g4274 (n2548, n_2034, n_2035);
  not g4275 (n_2036, n2548);
  and g4276 (n2549, n2530, n_2036);
  not g4277 (n_2037, n2530);
  and g4278 (n2550, n_2037, n2548);
  not g4279 (n_2038, n2549);
  not g4280 (n_2039, n2550);
  and g4281 (n2551, n_2038, n_2039);
  and g4282 (n2552, n2529, n2551);
  not g4283 (n_2040, n2529);
  not g4284 (n_2041, n2551);
  and g4285 (n2553, n_2040, n_2041);
  not g4286 (n_2042, n2552);
  not g4287 (n_2043, n2553);
  and g4288 (n2554, n_2042, n_2043);
  not g4289 (n_2044, n2518);
  not g4290 (n_2045, n2554);
  and g4291 (n2555, n_2044, n_2045);
  and g4292 (n2556, n2518, n2554);
  not g4293 (n_2046, n2555);
  not g4294 (n_2047, n2556);
  and g4295 (n2557, n_2046, n_2047);
  not g4296 (n_2048, n2516);
  and g4297 (n2558, n_2048, n2557);
  not g4298 (n_2049, n2557);
  and g4299 (n2559, n2516, n_2049);
  not g4300 (n_2050, n2558);
  not g4301 (n_2051, n2559);
  and g4302 (n2560, n_2050, n_2051);
  not g4303 (n_2052, n2505);
  and g4304 (n2561, n_2052, n2560);
  not g4305 (n_2053, n2560);
  and g4306 (n2562, n2505, n_2053);
  not g4307 (n_2054, n2561);
  not g4308 (n_2055, n2562);
  and g4309 (n2563, n_2054, n_2055);
  and g4310 (n2564, \b[10] , n1302);
  and g4311 (n2565, \b[8] , n1391);
  and g4312 (n2566, \b[9] , n1297);
  and g4318 (n2569, n738, n1305);
  not g4321 (n_2060, n2570);
  and g4322 (n2571, \a[17] , n_2060);
  not g4323 (n_2061, n2571);
  and g4324 (n2572, \a[17] , n_2061);
  and g4325 (n2573, n_2060, n_2061);
  not g4326 (n_2062, n2572);
  not g4327 (n_2063, n2573);
  and g4328 (n2574, n_2062, n_2063);
  not g4329 (n_2064, n2574);
  and g4330 (n2575, n2563, n_2064);
  not g4331 (n_2065, n2575);
  and g4332 (n2576, n2563, n_2065);
  and g4333 (n2577, n_2064, n_2065);
  not g4334 (n_2066, n2576);
  not g4335 (n_2067, n2577);
  and g4336 (n2578, n_2066, n_2067);
  and g4337 (n2579, n_1905, n_1909);
  and g4338 (n2580, n2578, n2579);
  not g4339 (n_2068, n2578);
  not g4340 (n_2069, n2579);
  and g4341 (n2581, n_2068, n_2069);
  not g4342 (n_2070, n2580);
  not g4343 (n_2071, n2581);
  and g4344 (n2582, n_2070, n_2071);
  and g4345 (n2583, \b[13] , n951);
  and g4346 (n2584, \b[11] , n1056);
  and g4347 (n2585, \b[12] , n946);
  and g4353 (n2588, n954, n1008);
  not g4356 (n_2076, n2589);
  and g4357 (n2590, \a[14] , n_2076);
  not g4358 (n_2077, n2590);
  and g4359 (n2591, \a[14] , n_2077);
  and g4360 (n2592, n_2076, n_2077);
  not g4361 (n_2078, n2591);
  not g4362 (n_2079, n2592);
  and g4363 (n2593, n_2078, n_2079);
  not g4364 (n_2080, n2582);
  and g4365 (n2594, n_2080, n2593);
  not g4366 (n_2081, n2593);
  and g4367 (n2595, n2582, n_2081);
  not g4368 (n_2082, n2594);
  not g4369 (n_2083, n2595);
  and g4370 (n2596, n_2082, n_2083);
  and g4371 (n2597, n_1914, n_1917);
  not g4372 (n_2084, n2597);
  and g4373 (n2598, n2596, n_2084);
  not g4374 (n_2085, n2596);
  and g4375 (n2599, n_2085, n2597);
  not g4376 (n_2086, n2598);
  not g4377 (n_2087, n2599);
  and g4378 (n2600, n_2086, n_2087);
  not g4379 (n_2088, n2503);
  and g4380 (n2601, n_2088, n2600);
  not g4381 (n_2089, n2601);
  and g4382 (n2602, n2600, n_2089);
  and g4383 (n2603, n_2088, n_2089);
  not g4384 (n_2090, n2602);
  not g4385 (n_2091, n2603);
  and g4386 (n2604, n_2090, n_2091);
  and g4387 (n2605, n_1920, n_1926);
  and g4388 (n2606, n2604, n2605);
  not g4389 (n_2092, n2604);
  not g4390 (n_2093, n2605);
  and g4391 (n2607, n_2092, n_2093);
  not g4392 (n_2094, n2606);
  not g4393 (n_2095, n2607);
  and g4394 (n2608, n_2094, n_2095);
  and g4395 (n2609, \b[19] , n511);
  and g4396 (n2610, \b[17] , n541);
  and g4397 (n2611, \b[18] , n506);
  and g4403 (n2614, n514, n1708);
  not g4406 (n_2100, n2615);
  and g4407 (n2616, \a[8] , n_2100);
  not g4408 (n_2101, n2616);
  and g4409 (n2617, \a[8] , n_2101);
  and g4410 (n2618, n_2100, n_2101);
  not g4411 (n_2102, n2617);
  not g4412 (n_2103, n2618);
  and g4413 (n2619, n_2102, n_2103);
  not g4414 (n_2104, n2619);
  and g4415 (n2620, n2608, n_2104);
  not g4416 (n_2105, n2620);
  and g4417 (n2621, n2608, n_2105);
  and g4418 (n2622, n_2104, n_2105);
  not g4419 (n_2106, n2621);
  not g4420 (n_2107, n2622);
  and g4421 (n2623, n_2106, n_2107);
  and g4422 (n2624, n_1938, n_1941);
  not g4423 (n_2108, n2623);
  not g4424 (n_2109, n2624);
  and g4425 (n2625, n_2108, n_2109);
  not g4426 (n_2110, n2625);
  and g4427 (n2626, n_2108, n_2110);
  and g4428 (n2627, n_2109, n_2110);
  not g4429 (n_2111, n2626);
  not g4430 (n_2112, n2627);
  and g4431 (n2628, n_2111, n_2112);
  and g4432 (n2629, \b[22] , n362);
  and g4433 (n2630, \b[20] , n403);
  and g4434 (n2631, \b[21] , n357);
  and g4440 (n2634, n365, n2145);
  not g4443 (n_2117, n2635);
  and g4444 (n2636, \a[5] , n_2117);
  not g4445 (n_2118, n2636);
  and g4446 (n2637, \a[5] , n_2118);
  and g4447 (n2638, n_2117, n_2118);
  not g4448 (n_2119, n2637);
  not g4449 (n_2120, n2638);
  and g4450 (n2639, n_2119, n_2120);
  not g4451 (n_2121, n2628);
  and g4452 (n2640, n_2121, n2639);
  not g4453 (n_2122, n2639);
  and g4454 (n2641, n2628, n_2122);
  not g4455 (n_2123, n2640);
  not g4456 (n_2124, n2641);
  and g4457 (n2642, n_2123, n_2124);
  not g4458 (n_2125, n2492);
  not g4459 (n_2126, n2642);
  and g4460 (n2643, n_2125, n_2126);
  and g4461 (n2644, n2492, n2642);
  not g4462 (n_2127, n2643);
  not g4463 (n_2128, n2644);
  and g4464 (n2645, n_2127, n_2128);
  not g4465 (n_2129, n2491);
  and g4466 (n2646, n_2129, n2645);
  not g4467 (n_2130, n2645);
  and g4468 (n2647, n2491, n_2130);
  not g4469 (n_2131, n2646);
  not g4470 (n_2132, n2647);
  and g4471 (n2648, n_2131, n_2132);
  not g4472 (n_2133, n2473);
  and g4473 (n2649, n_2133, n2648);
  not g4474 (n_2134, n2648);
  and g4475 (n2650, n2473, n_2134);
  not g4476 (n_2135, n2649);
  not g4477 (n_2136, n2650);
  and g4478 (\f[25] , n_2135, n_2136);
  and g4479 (n2652, n_2131, n_2135);
  and g4480 (n2653, n_2121, n_2122);
  not g4481 (n_2137, n2653);
  and g4482 (n2654, n_2127, n_2137);
  and g4483 (n2655, n_2089, n_2095);
  and g4484 (n2656, n_2083, n_2086);
  and g4485 (n2657, \b[14] , n951);
  and g4486 (n2658, \b[12] , n1056);
  and g4487 (n2659, \b[13] , n946);
  and g4493 (n2662, n954, n1034);
  not g4496 (n_2142, n2663);
  and g4497 (n2664, \a[14] , n_2142);
  not g4498 (n_2143, n2664);
  and g4499 (n2665, \a[14] , n_2143);
  and g4500 (n2666, n_2142, n_2143);
  not g4501 (n_2144, n2665);
  not g4502 (n_2145, n2666);
  and g4503 (n2667, n_2144, n_2145);
  and g4504 (n2668, n_2065, n_2071);
  and g4505 (n2669, \b[11] , n1302);
  and g4506 (n2670, \b[9] , n1391);
  and g4507 (n2671, \b[10] , n1297);
  and g4513 (n2674, n818, n1305);
  not g4516 (n_2150, n2675);
  and g4517 (n2676, \a[17] , n_2150);
  not g4518 (n_2151, n2676);
  and g4519 (n2677, \a[17] , n_2151);
  and g4520 (n2678, n_2150, n_2151);
  not g4521 (n_2152, n2677);
  not g4522 (n_2153, n2678);
  and g4523 (n2679, n_2152, n_2153);
  and g4524 (n2680, n_2050, n_2054);
  and g4525 (n2681, n_2040, n2551);
  not g4526 (n_2154, n2681);
  and g4527 (n2682, n_2046, n_2154);
  and g4528 (n2683, \b[2] , n2539);
  and g4529 (n2684, n2365, n_2030);
  and g4530 (n2685, n2533, n2684);
  and g4531 (n2686, \b[0] , n2685);
  and g4532 (n2687, \b[1] , n2534);
  and g4538 (n2690, n296, n2542);
  not g4541 (n_2159, n2691);
  and g4542 (n2692, \a[26] , n_2159);
  not g4543 (n_2160, n2692);
  and g4544 (n2693, \a[26] , n_2160);
  and g4545 (n2694, n_2159, n_2160);
  not g4546 (n_2161, n2693);
  not g4547 (n_2162, n2694);
  and g4548 (n2695, n_2161, n_2162);
  and g4549 (n2696, n_2038, n2695);
  not g4550 (n_2163, n2695);
  and g4551 (n2697, n2549, n_2163);
  not g4552 (n_2164, n2696);
  not g4553 (n_2165, n2697);
  and g4554 (n2698, n_2164, n_2165);
  and g4555 (n2699, \b[5] , n2048);
  and g4556 (n2700, \b[3] , n2198);
  and g4557 (n2701, \b[4] , n2043);
  and g4563 (n2704, n394, n2051);
  not g4566 (n_2170, n2705);
  and g4567 (n2706, \a[23] , n_2170);
  not g4568 (n_2171, n2706);
  and g4569 (n2707, \a[23] , n_2171);
  and g4570 (n2708, n_2170, n_2171);
  not g4571 (n_2172, n2707);
  not g4572 (n_2173, n2708);
  and g4573 (n2709, n_2172, n_2173);
  not g4574 (n_2174, n2709);
  and g4575 (n2710, n2698, n_2174);
  not g4576 (n_2175, n2698);
  and g4577 (n2711, n_2175, n2709);
  not g4578 (n_2176, n2682);
  not g4579 (n_2177, n2711);
  and g4580 (n2712, n_2176, n_2177);
  not g4581 (n_2178, n2710);
  and g4582 (n2713, n_2178, n2712);
  not g4583 (n_2179, n2713);
  and g4584 (n2714, n_2176, n_2179);
  and g4585 (n2715, n_2178, n_2179);
  and g4586 (n2716, n_2177, n2715);
  not g4587 (n_2180, n2714);
  not g4588 (n_2181, n2716);
  and g4589 (n2717, n_2180, n_2181);
  and g4590 (n2718, \b[8] , n1627);
  and g4591 (n2719, \b[6] , n1763);
  and g4592 (n2720, \b[7] , n1622);
  and g4598 (n2723, n585, n1630);
  not g4601 (n_2186, n2724);
  and g4602 (n2725, \a[20] , n_2186);
  not g4603 (n_2187, n2725);
  and g4604 (n2726, \a[20] , n_2187);
  and g4605 (n2727, n_2186, n_2187);
  not g4606 (n_2188, n2726);
  not g4607 (n_2189, n2727);
  and g4608 (n2728, n_2188, n_2189);
  and g4609 (n2729, n2717, n2728);
  not g4610 (n_2190, n2717);
  not g4611 (n_2191, n2728);
  and g4612 (n2730, n_2190, n_2191);
  not g4613 (n_2192, n2729);
  not g4614 (n_2193, n2730);
  and g4615 (n2731, n_2192, n_2193);
  not g4616 (n_2194, n2680);
  and g4617 (n2732, n_2194, n2731);
  not g4618 (n_2195, n2731);
  and g4619 (n2733, n2680, n_2195);
  not g4620 (n_2196, n2732);
  not g4621 (n_2197, n2733);
  and g4622 (n2734, n_2196, n_2197);
  not g4623 (n_2198, n2734);
  and g4624 (n2735, n2679, n_2198);
  not g4625 (n_2199, n2679);
  and g4626 (n2736, n_2199, n2734);
  not g4627 (n_2200, n2735);
  not g4628 (n_2201, n2736);
  and g4629 (n2737, n_2200, n_2201);
  not g4630 (n_2202, n2668);
  and g4631 (n2738, n_2202, n2737);
  not g4632 (n_2203, n2737);
  and g4633 (n2739, n2668, n_2203);
  not g4634 (n_2204, n2738);
  not g4635 (n_2205, n2739);
  and g4636 (n2740, n_2204, n_2205);
  not g4637 (n_2206, n2667);
  and g4638 (n2741, n_2206, n2740);
  not g4639 (n_2207, n2741);
  and g4640 (n2742, n2740, n_2207);
  and g4641 (n2743, n_2206, n_2207);
  not g4642 (n_2208, n2742);
  not g4643 (n_2209, n2743);
  and g4644 (n2744, n_2208, n_2209);
  not g4645 (n_2210, n2656);
  and g4646 (n2745, n_2210, n2744);
  not g4647 (n_2211, n2744);
  and g4648 (n2746, n2656, n_2211);
  not g4649 (n_2212, n2745);
  not g4650 (n_2213, n2746);
  and g4651 (n2747, n_2212, n_2213);
  and g4652 (n2748, \b[17] , n700);
  and g4653 (n2749, \b[15] , n767);
  and g4654 (n2750, \b[16] , n695);
  and g4660 (n2753, n703, n1356);
  not g4663 (n_2218, n2754);
  and g4664 (n2755, \a[11] , n_2218);
  not g4665 (n_2219, n2755);
  and g4666 (n2756, \a[11] , n_2219);
  and g4667 (n2757, n_2218, n_2219);
  not g4668 (n_2220, n2756);
  not g4669 (n_2221, n2757);
  and g4670 (n2758, n_2220, n_2221);
  not g4671 (n_2222, n2747);
  not g4672 (n_2223, n2758);
  and g4673 (n2759, n_2222, n_2223);
  and g4674 (n2760, n2747, n2758);
  not g4675 (n_2224, n2759);
  not g4676 (n_2225, n2760);
  and g4677 (n2761, n_2224, n_2225);
  not g4678 (n_2226, n2761);
  and g4679 (n2762, n2655, n_2226);
  not g4680 (n_2227, n2655);
  and g4681 (n2763, n_2227, n2761);
  not g4682 (n_2228, n2762);
  not g4683 (n_2229, n2763);
  and g4684 (n2764, n_2228, n_2229);
  and g4685 (n2765, \b[20] , n511);
  and g4686 (n2766, \b[18] , n541);
  and g4687 (n2767, \b[19] , n506);
  and g4693 (n2770, n514, n1846);
  not g4696 (n_2234, n2771);
  and g4697 (n2772, \a[8] , n_2234);
  not g4698 (n_2235, n2772);
  and g4699 (n2773, \a[8] , n_2235);
  and g4700 (n2774, n_2234, n_2235);
  not g4701 (n_2236, n2773);
  not g4702 (n_2237, n2774);
  and g4703 (n2775, n_2236, n_2237);
  not g4704 (n_2238, n2775);
  and g4705 (n2776, n2764, n_2238);
  not g4706 (n_2239, n2776);
  and g4707 (n2777, n2764, n_2239);
  and g4708 (n2778, n_2238, n_2239);
  not g4709 (n_2240, n2777);
  not g4710 (n_2241, n2778);
  and g4711 (n2779, n_2240, n_2241);
  and g4712 (n2780, n_2105, n_2110);
  and g4713 (n2781, n2779, n2780);
  not g4714 (n_2242, n2779);
  not g4715 (n_2243, n2780);
  and g4716 (n2782, n_2242, n_2243);
  not g4717 (n_2244, n2781);
  not g4718 (n_2245, n2782);
  and g4719 (n2783, n_2244, n_2245);
  and g4720 (n2784, \b[23] , n362);
  and g4721 (n2785, \b[21] , n403);
  and g4722 (n2786, \b[22] , n357);
  and g4728 (n2789, n365, n2300);
  not g4731 (n_2250, n2790);
  and g4732 (n2791, \a[5] , n_2250);
  not g4733 (n_2251, n2791);
  and g4734 (n2792, \a[5] , n_2251);
  and g4735 (n2793, n_2250, n_2251);
  not g4736 (n_2252, n2792);
  not g4737 (n_2253, n2793);
  and g4738 (n2794, n_2252, n_2253);
  not g4739 (n_2254, n2794);
  and g4740 (n2795, n2783, n_2254);
  not g4741 (n_2255, n2795);
  and g4742 (n2796, n2783, n_2255);
  and g4743 (n2797, n_2254, n_2255);
  not g4744 (n_2256, n2796);
  not g4745 (n_2257, n2797);
  and g4746 (n2798, n_2256, n_2257);
  not g4747 (n_2258, n2654);
  and g4748 (n2799, n_2258, n2798);
  not g4749 (n_2259, n2798);
  and g4750 (n2800, n2654, n_2259);
  not g4751 (n_2260, n2799);
  not g4752 (n_2261, n2800);
  and g4753 (n2801, n_2260, n_2261);
  and g4754 (n2802, \b[26] , n266);
  and g4755 (n2803, \b[24] , n284);
  and g4756 (n2804, \b[25] , n261);
  and g4762 (n2807, n_1983, n_1986);
  not g4763 (n_2266, \b[26] );
  and g4764 (n2808, n_1981, n_2266);
  and g4765 (n2809, \b[25] , \b[26] );
  not g4766 (n_2267, n2808);
  not g4767 (n_2268, n2809);
  and g4768 (n2810, n_2267, n_2268);
  not g4769 (n_2269, n2807);
  and g4770 (n2811, n_2269, n2810);
  not g4771 (n_2270, n2810);
  and g4772 (n2812, n2807, n_2270);
  not g4773 (n_2271, n2811);
  not g4774 (n_2272, n2812);
  and g4775 (n2813, n_2271, n_2272);
  and g4776 (n2814, n269, n2813);
  not g4779 (n_2274, n2815);
  and g4780 (n2816, \a[2] , n_2274);
  not g4781 (n_2275, n2816);
  and g4782 (n2817, \a[2] , n_2275);
  and g4783 (n2818, n_2274, n_2275);
  not g4784 (n_2276, n2817);
  not g4785 (n_2277, n2818);
  and g4786 (n2819, n_2276, n_2277);
  not g4787 (n_2278, n2801);
  not g4788 (n_2279, n2819);
  and g4789 (n2820, n_2278, n_2279);
  and g4790 (n2821, n2801, n2819);
  not g4791 (n_2280, n2820);
  not g4792 (n_2281, n2821);
  and g4793 (n2822, n_2280, n_2281);
  not g4794 (n_2282, n2652);
  and g4795 (n2823, n_2282, n2822);
  not g4796 (n_2283, n2822);
  and g4797 (n2824, n2652, n_2283);
  not g4798 (n_2284, n2823);
  not g4799 (n_2285, n2824);
  and g4800 (\f[26] , n_2284, n_2285);
  and g4801 (n2826, n_2280, n_2284);
  and g4802 (n2827, \b[24] , n362);
  and g4803 (n2828, \b[22] , n403);
  and g4804 (n2829, \b[23] , n357);
  and g4810 (n2832, n365, n2458);
  not g4813 (n_2290, n2833);
  and g4814 (n2834, \a[5] , n_2290);
  not g4815 (n_2291, n2834);
  and g4816 (n2835, \a[5] , n_2291);
  and g4817 (n2836, n_2290, n_2291);
  not g4818 (n_2292, n2835);
  not g4819 (n_2293, n2836);
  and g4820 (n2837, n_2292, n_2293);
  and g4821 (n2838, \b[15] , n951);
  and g4822 (n2839, \b[13] , n1056);
  and g4823 (n2840, \b[14] , n946);
  and g4829 (n2843, n954, n1131);
  not g4832 (n_2298, n2844);
  and g4833 (n2845, \a[14] , n_2298);
  not g4834 (n_2299, n2845);
  and g4835 (n2846, \a[14] , n_2299);
  and g4836 (n2847, n_2298, n_2299);
  not g4837 (n_2300, n2846);
  not g4838 (n_2301, n2847);
  and g4839 (n2848, n_2300, n_2301);
  and g4840 (n2849, n_2201, n_2204);
  and g4841 (n2850, \b[12] , n1302);
  and g4842 (n2851, \b[10] , n1391);
  and g4843 (n2852, \b[11] , n1297);
  and g4849 (n2855, n842, n1305);
  not g4852 (n_2306, n2856);
  and g4853 (n2857, \a[17] , n_2306);
  not g4854 (n_2307, n2857);
  and g4855 (n2858, \a[17] , n_2307);
  and g4856 (n2859, n_2306, n_2307);
  not g4857 (n_2308, n2858);
  not g4858 (n_2309, n2859);
  and g4859 (n2860, n_2308, n_2309);
  and g4860 (n2861, n_2193, n_2196);
  and g4861 (n2862, \b[6] , n2048);
  and g4862 (n2863, \b[4] , n2198);
  and g4863 (n2864, \b[5] , n2043);
  and g4869 (n2867, n459, n2051);
  not g4872 (n_2314, n2868);
  and g4873 (n2869, \a[23] , n_2314);
  not g4874 (n_2315, n2869);
  and g4875 (n2870, \a[23] , n_2315);
  and g4876 (n2871, n_2314, n_2315);
  not g4877 (n_2316, n2870);
  not g4878 (n_2317, n2871);
  and g4879 (n2872, n_2316, n_2317);
  not g4880 (n_2319, \a[27] );
  and g4881 (n2873, \a[26] , n_2319);
  and g4882 (n2874, n_2025, \a[27] );
  not g4883 (n_2320, n2873);
  not g4884 (n_2321, n2874);
  and g4885 (n2875, n_2320, n_2321);
  not g4886 (n_2322, n2875);
  and g4887 (n2876, \b[0] , n_2322);
  and g4888 (n2877, n_2165, n2876);
  not g4889 (n_2323, n2876);
  and g4890 (n2878, n2697, n_2323);
  not g4891 (n_2324, n2877);
  not g4892 (n_2325, n2878);
  and g4893 (n2879, n_2324, n_2325);
  and g4894 (n2880, \b[3] , n2539);
  and g4895 (n2881, \b[1] , n2685);
  and g4896 (n2882, \b[2] , n2534);
  and g4902 (n2885, n318, n2542);
  not g4905 (n_2330, n2886);
  and g4906 (n2887, \a[26] , n_2330);
  not g4907 (n_2331, n2887);
  and g4908 (n2888, \a[26] , n_2331);
  and g4909 (n2889, n_2330, n_2331);
  not g4910 (n_2332, n2888);
  not g4911 (n_2333, n2889);
  and g4912 (n2890, n_2332, n_2333);
  not g4913 (n_2334, n2879);
  not g4914 (n_2335, n2890);
  and g4915 (n2891, n_2334, n_2335);
  and g4916 (n2892, n2879, n2890);
  not g4917 (n_2336, n2891);
  not g4918 (n_2337, n2892);
  and g4919 (n2893, n_2336, n_2337);
  not g4920 (n_2338, n2872);
  and g4921 (n2894, n_2338, n2893);
  not g4922 (n_2339, n2894);
  and g4923 (n2895, n2893, n_2339);
  and g4924 (n2896, n_2338, n_2339);
  not g4925 (n_2340, n2895);
  not g4926 (n_2341, n2896);
  and g4927 (n2897, n_2340, n_2341);
  not g4928 (n_2342, n2715);
  and g4929 (n2898, n_2342, n2897);
  not g4930 (n_2343, n2897);
  and g4931 (n2899, n2715, n_2343);
  not g4932 (n_2344, n2898);
  not g4933 (n_2345, n2899);
  and g4934 (n2900, n_2344, n_2345);
  and g4935 (n2901, \b[9] , n1627);
  and g4936 (n2902, \b[7] , n1763);
  and g4937 (n2903, \b[8] , n1622);
  and g4943 (n2906, n651, n1630);
  not g4946 (n_2350, n2907);
  and g4947 (n2908, \a[20] , n_2350);
  not g4948 (n_2351, n2908);
  and g4949 (n2909, \a[20] , n_2351);
  and g4950 (n2910, n_2350, n_2351);
  not g4951 (n_2352, n2909);
  not g4952 (n_2353, n2910);
  and g4953 (n2911, n_2352, n_2353);
  not g4954 (n_2354, n2900);
  not g4955 (n_2355, n2911);
  and g4956 (n2912, n_2354, n_2355);
  and g4957 (n2913, n2900, n2911);
  not g4958 (n_2356, n2912);
  not g4959 (n_2357, n2913);
  and g4960 (n2914, n_2356, n_2357);
  not g4961 (n_2358, n2861);
  and g4962 (n2915, n_2358, n2914);
  not g4963 (n_2359, n2914);
  and g4964 (n2916, n2861, n_2359);
  not g4965 (n_2360, n2915);
  not g4966 (n_2361, n2916);
  and g4967 (n2917, n_2360, n_2361);
  not g4968 (n_2362, n2917);
  and g4969 (n2918, n2860, n_2362);
  not g4970 (n_2363, n2860);
  and g4971 (n2919, n_2363, n2917);
  not g4972 (n_2364, n2918);
  not g4973 (n_2365, n2919);
  and g4974 (n2920, n_2364, n_2365);
  not g4975 (n_2366, n2849);
  and g4976 (n2921, n_2366, n2920);
  not g4977 (n_2367, n2920);
  and g4978 (n2922, n2849, n_2367);
  not g4979 (n_2368, n2921);
  not g4980 (n_2369, n2922);
  and g4981 (n2923, n_2368, n_2369);
  not g4982 (n_2370, n2848);
  and g4983 (n2924, n_2370, n2923);
  not g4984 (n_2371, n2924);
  and g4985 (n2925, n2923, n_2371);
  and g4986 (n2926, n_2370, n_2371);
  not g4987 (n_2372, n2925);
  not g4988 (n_2373, n2926);
  and g4989 (n2927, n_2372, n_2373);
  and g4990 (n2928, n_2210, n_2211);
  not g4991 (n_2374, n2928);
  and g4992 (n2929, n_2207, n_2374);
  and g4993 (n2930, n2927, n2929);
  not g4994 (n_2375, n2927);
  not g4995 (n_2376, n2929);
  and g4996 (n2931, n_2375, n_2376);
  not g4997 (n_2377, n2930);
  not g4998 (n_2378, n2931);
  and g4999 (n2932, n_2377, n_2378);
  and g5000 (n2933, \b[18] , n700);
  and g5001 (n2934, \b[16] , n767);
  and g5002 (n2935, \b[17] , n695);
  and g5008 (n2938, n703, n1566);
  not g5011 (n_2383, n2939);
  and g5012 (n2940, \a[11] , n_2383);
  not g5013 (n_2384, n2940);
  and g5014 (n2941, \a[11] , n_2384);
  and g5015 (n2942, n_2383, n_2384);
  not g5016 (n_2385, n2941);
  not g5017 (n_2386, n2942);
  and g5018 (n2943, n_2385, n_2386);
  not g5019 (n_2387, n2943);
  and g5020 (n2944, n2932, n_2387);
  not g5021 (n_2388, n2944);
  and g5022 (n2945, n2932, n_2388);
  and g5023 (n2946, n_2387, n_2388);
  not g5024 (n_2389, n2945);
  not g5025 (n_2390, n2946);
  and g5026 (n2947, n_2389, n_2390);
  and g5027 (n2948, n_2224, n_2229);
  and g5028 (n2949, n2947, n2948);
  not g5029 (n_2391, n2947);
  not g5030 (n_2392, n2948);
  and g5031 (n2950, n_2391, n_2392);
  not g5032 (n_2393, n2949);
  not g5033 (n_2394, n2950);
  and g5034 (n2951, n_2393, n_2394);
  and g5035 (n2952, \b[21] , n511);
  and g5036 (n2953, \b[19] , n541);
  and g5037 (n2954, \b[20] , n506);
  and g5043 (n2957, n514, n1984);
  not g5046 (n_2399, n2958);
  and g5047 (n2959, \a[8] , n_2399);
  not g5048 (n_2400, n2959);
  and g5049 (n2960, \a[8] , n_2400);
  and g5050 (n2961, n_2399, n_2400);
  not g5051 (n_2401, n2960);
  not g5052 (n_2402, n2961);
  and g5053 (n2962, n_2401, n_2402);
  not g5054 (n_2403, n2951);
  and g5055 (n2963, n_2403, n2962);
  not g5056 (n_2404, n2962);
  and g5057 (n2964, n2951, n_2404);
  not g5058 (n_2405, n2963);
  not g5059 (n_2406, n2964);
  and g5060 (n2965, n_2405, n_2406);
  and g5061 (n2966, n_2239, n_2245);
  not g5062 (n_2407, n2966);
  and g5063 (n2967, n2965, n_2407);
  not g5064 (n_2408, n2965);
  and g5065 (n2968, n_2408, n2966);
  not g5066 (n_2409, n2967);
  not g5067 (n_2410, n2968);
  and g5068 (n2969, n_2409, n_2410);
  not g5069 (n_2411, n2837);
  and g5070 (n2970, n_2411, n2969);
  not g5071 (n_2412, n2970);
  and g5072 (n2971, n2969, n_2412);
  and g5073 (n2972, n_2411, n_2412);
  not g5074 (n_2413, n2971);
  not g5075 (n_2414, n2972);
  and g5076 (n2973, n_2413, n_2414);
  and g5077 (n2974, n_2258, n_2259);
  not g5078 (n_2415, n2974);
  and g5079 (n2975, n_2255, n_2415);
  and g5080 (n2976, n2973, n2975);
  not g5081 (n_2416, n2973);
  not g5082 (n_2417, n2975);
  and g5083 (n2977, n_2416, n_2417);
  not g5084 (n_2418, n2976);
  not g5085 (n_2419, n2977);
  and g5086 (n2978, n_2418, n_2419);
  and g5087 (n2979, \b[27] , n266);
  and g5088 (n2980, \b[25] , n284);
  and g5089 (n2981, \b[26] , n261);
  and g5095 (n2984, n_2268, n_2271);
  not g5096 (n_2424, \b[27] );
  and g5097 (n2985, n_2266, n_2424);
  and g5098 (n2986, \b[26] , \b[27] );
  not g5099 (n_2425, n2985);
  not g5100 (n_2426, n2986);
  and g5101 (n2987, n_2425, n_2426);
  not g5102 (n_2427, n2984);
  and g5103 (n2988, n_2427, n2987);
  not g5104 (n_2428, n2987);
  and g5105 (n2989, n2984, n_2428);
  not g5106 (n_2429, n2988);
  not g5107 (n_2430, n2989);
  and g5108 (n2990, n_2429, n_2430);
  and g5109 (n2991, n269, n2990);
  not g5112 (n_2432, n2992);
  and g5113 (n2993, \a[2] , n_2432);
  not g5114 (n_2433, n2993);
  and g5115 (n2994, \a[2] , n_2433);
  and g5116 (n2995, n_2432, n_2433);
  not g5117 (n_2434, n2994);
  not g5118 (n_2435, n2995);
  and g5119 (n2996, n_2434, n_2435);
  not g5120 (n_2436, n2978);
  and g5121 (n2997, n_2436, n2996);
  not g5122 (n_2437, n2996);
  and g5123 (n2998, n2978, n_2437);
  not g5124 (n_2438, n2997);
  not g5125 (n_2439, n2998);
  and g5126 (n2999, n_2438, n_2439);
  not g5127 (n_2440, n2826);
  and g5128 (n3000, n_2440, n2999);
  not g5129 (n_2441, n2999);
  and g5130 (n3001, n2826, n_2441);
  not g5131 (n_2442, n3000);
  not g5132 (n_2443, n3001);
  and g5133 (\f[27] , n_2442, n_2443);
  and g5134 (n3003, n_2439, n_2442);
  and g5135 (n3004, \b[25] , n362);
  and g5136 (n3005, \b[23] , n403);
  and g5137 (n3006, \b[24] , n357);
  and g5143 (n3009, n365, n2485);
  not g5146 (n_2448, n3010);
  and g5147 (n3011, \a[5] , n_2448);
  not g5148 (n_2449, n3011);
  and g5149 (n3012, \a[5] , n_2449);
  and g5150 (n3013, n_2448, n_2449);
  not g5151 (n_2450, n3012);
  not g5152 (n_2451, n3013);
  and g5153 (n3014, n_2450, n_2451);
  and g5154 (n3015, n_2342, n_2343);
  not g5155 (n_2452, n3015);
  and g5156 (n3016, n_2339, n_2452);
  and g5157 (n3017, \b[7] , n2048);
  and g5158 (n3018, \b[5] , n2198);
  and g5159 (n3019, \b[6] , n2043);
  and g5165 (n3022, n484, n2051);
  not g5168 (n_2457, n3023);
  and g5169 (n3024, \a[23] , n_2457);
  not g5170 (n_2458, n3024);
  and g5171 (n3025, \a[23] , n_2458);
  and g5172 (n3026, n_2457, n_2458);
  not g5173 (n_2459, n3025);
  not g5174 (n_2460, n3026);
  and g5175 (n3027, n_2459, n_2460);
  and g5176 (n3028, n2697, n2876);
  not g5177 (n_2461, n3028);
  and g5178 (n3029, n_2336, n_2461);
  and g5179 (n3030, \b[4] , n2539);
  and g5180 (n3031, \b[2] , n2685);
  and g5181 (n3032, \b[3] , n2534);
  and g5187 (n3035, n346, n2542);
  not g5190 (n_2466, n3036);
  and g5191 (n3037, \a[26] , n_2466);
  not g5192 (n_2467, n3037);
  and g5193 (n3038, \a[26] , n_2467);
  and g5194 (n3039, n_2466, n_2467);
  not g5195 (n_2468, n3038);
  not g5196 (n_2469, n3039);
  and g5197 (n3040, n_2468, n_2469);
  and g5198 (n3041, \a[29] , n_2323);
  and g5199 (n3042, n_2319, \a[28] );
  not g5200 (n_2472, \a[28] );
  and g5201 (n3043, \a[27] , n_2472);
  not g5202 (n_2473, n3042);
  not g5203 (n_2474, n3043);
  and g5204 (n3044, n_2473, n_2474);
  not g5205 (n_2475, n3044);
  and g5206 (n3045, n2875, n_2475);
  and g5207 (n3046, \b[0] , n3045);
  and g5208 (n3047, n_2472, \a[29] );
  not g5209 (n_2476, \a[29] );
  and g5210 (n3048, \a[28] , n_2476);
  not g5211 (n_2477, n3047);
  not g5212 (n_2478, n3048);
  and g5213 (n3049, n_2477, n_2478);
  and g5214 (n3050, n_2322, n3049);
  and g5215 (n3051, \b[1] , n3050);
  not g5216 (n_2479, n3046);
  not g5217 (n_2480, n3051);
  and g5218 (n3052, n_2479, n_2480);
  not g5219 (n_2481, n3049);
  and g5220 (n3053, n_2322, n_2481);
  and g5221 (n3054, n_21, n3053);
  not g5222 (n_2482, n3054);
  and g5223 (n3055, n3052, n_2482);
  not g5224 (n_2483, n3055);
  and g5225 (n3056, \a[29] , n_2483);
  not g5226 (n_2484, n3056);
  and g5227 (n3057, \a[29] , n_2484);
  and g5228 (n3058, n_2483, n_2484);
  not g5229 (n_2485, n3057);
  not g5230 (n_2486, n3058);
  and g5231 (n3059, n_2485, n_2486);
  not g5232 (n_2487, n3059);
  and g5233 (n3060, n3041, n_2487);
  not g5234 (n_2488, n3041);
  and g5235 (n3061, n_2488, n3059);
  not g5236 (n_2489, n3060);
  not g5237 (n_2490, n3061);
  and g5238 (n3062, n_2489, n_2490);
  and g5239 (n3063, n3040, n3062);
  not g5240 (n_2491, n3040);
  not g5241 (n_2492, n3062);
  and g5242 (n3064, n_2491, n_2492);
  not g5243 (n_2493, n3063);
  not g5244 (n_2494, n3064);
  and g5245 (n3065, n_2493, n_2494);
  not g5246 (n_2495, n3029);
  not g5247 (n_2496, n3065);
  and g5248 (n3066, n_2495, n_2496);
  and g5249 (n3067, n3029, n3065);
  not g5250 (n_2497, n3066);
  not g5251 (n_2498, n3067);
  and g5252 (n3068, n_2497, n_2498);
  not g5253 (n_2499, n3027);
  and g5254 (n3069, n_2499, n3068);
  not g5255 (n_2500, n3068);
  and g5256 (n3070, n3027, n_2500);
  not g5257 (n_2501, n3069);
  not g5258 (n_2502, n3070);
  and g5259 (n3071, n_2501, n_2502);
  not g5260 (n_2503, n3016);
  and g5261 (n3072, n_2503, n3071);
  not g5262 (n_2504, n3071);
  and g5263 (n3073, n3016, n_2504);
  not g5264 (n_2505, n3072);
  not g5265 (n_2506, n3073);
  and g5266 (n3074, n_2505, n_2506);
  and g5267 (n3075, \b[10] , n1627);
  and g5268 (n3076, \b[8] , n1763);
  and g5269 (n3077, \b[9] , n1622);
  and g5275 (n3080, n738, n1630);
  not g5278 (n_2511, n3081);
  and g5279 (n3082, \a[20] , n_2511);
  not g5280 (n_2512, n3082);
  and g5281 (n3083, \a[20] , n_2512);
  and g5282 (n3084, n_2511, n_2512);
  not g5283 (n_2513, n3083);
  not g5284 (n_2514, n3084);
  and g5285 (n3085, n_2513, n_2514);
  not g5286 (n_2515, n3085);
  and g5287 (n3086, n3074, n_2515);
  not g5288 (n_2516, n3086);
  and g5289 (n3087, n3074, n_2516);
  and g5290 (n3088, n_2515, n_2516);
  not g5291 (n_2517, n3087);
  not g5292 (n_2518, n3088);
  and g5293 (n3089, n_2517, n_2518);
  and g5294 (n3090, n_2356, n_2360);
  and g5295 (n3091, n3089, n3090);
  not g5296 (n_2519, n3089);
  not g5297 (n_2520, n3090);
  and g5298 (n3092, n_2519, n_2520);
  not g5299 (n_2521, n3091);
  not g5300 (n_2522, n3092);
  and g5301 (n3093, n_2521, n_2522);
  and g5302 (n3094, \b[13] , n1302);
  and g5303 (n3095, \b[11] , n1391);
  and g5304 (n3096, \b[12] , n1297);
  and g5310 (n3099, n1008, n1305);
  not g5313 (n_2527, n3100);
  and g5314 (n3101, \a[17] , n_2527);
  not g5315 (n_2528, n3101);
  and g5316 (n3102, \a[17] , n_2528);
  and g5317 (n3103, n_2527, n_2528);
  not g5318 (n_2529, n3102);
  not g5319 (n_2530, n3103);
  and g5320 (n3104, n_2529, n_2530);
  not g5321 (n_2531, n3104);
  and g5322 (n3105, n3093, n_2531);
  not g5323 (n_2532, n3105);
  and g5324 (n3106, n3093, n_2532);
  and g5325 (n3107, n_2531, n_2532);
  not g5326 (n_2533, n3106);
  not g5327 (n_2534, n3107);
  and g5328 (n3108, n_2533, n_2534);
  and g5329 (n3109, n_2365, n_2368);
  not g5330 (n_2535, n3108);
  not g5331 (n_2536, n3109);
  and g5332 (n3110, n_2535, n_2536);
  not g5333 (n_2537, n3110);
  and g5334 (n3111, n_2535, n_2537);
  and g5335 (n3112, n_2536, n_2537);
  not g5336 (n_2538, n3111);
  not g5337 (n_2539, n3112);
  and g5338 (n3113, n_2538, n_2539);
  and g5339 (n3114, \b[16] , n951);
  and g5340 (n3115, \b[14] , n1056);
  and g5341 (n3116, \b[15] , n946);
  and g5347 (n3119, n954, n1237);
  not g5350 (n_2544, n3120);
  and g5351 (n3121, \a[14] , n_2544);
  not g5352 (n_2545, n3121);
  and g5353 (n3122, \a[14] , n_2545);
  and g5354 (n3123, n_2544, n_2545);
  not g5355 (n_2546, n3122);
  not g5356 (n_2547, n3123);
  and g5357 (n3124, n_2546, n_2547);
  not g5358 (n_2548, n3113);
  not g5359 (n_2549, n3124);
  and g5360 (n3125, n_2548, n_2549);
  not g5361 (n_2550, n3125);
  and g5362 (n3126, n_2548, n_2550);
  and g5363 (n3127, n_2549, n_2550);
  not g5364 (n_2551, n3126);
  not g5365 (n_2552, n3127);
  and g5366 (n3128, n_2551, n_2552);
  and g5367 (n3129, n_2371, n_2378);
  and g5368 (n3130, n3128, n3129);
  not g5369 (n_2553, n3128);
  not g5370 (n_2554, n3129);
  and g5371 (n3131, n_2553, n_2554);
  not g5372 (n_2555, n3130);
  not g5373 (n_2556, n3131);
  and g5374 (n3132, n_2555, n_2556);
  and g5375 (n3133, \b[19] , n700);
  and g5376 (n3134, \b[17] , n767);
  and g5377 (n3135, \b[18] , n695);
  and g5383 (n3138, n703, n1708);
  not g5386 (n_2561, n3139);
  and g5387 (n3140, \a[11] , n_2561);
  not g5388 (n_2562, n3140);
  and g5389 (n3141, \a[11] , n_2562);
  and g5390 (n3142, n_2561, n_2562);
  not g5391 (n_2563, n3141);
  not g5392 (n_2564, n3142);
  and g5393 (n3143, n_2563, n_2564);
  not g5394 (n_2565, n3143);
  and g5395 (n3144, n3132, n_2565);
  not g5396 (n_2566, n3144);
  and g5397 (n3145, n3132, n_2566);
  and g5398 (n3146, n_2565, n_2566);
  not g5399 (n_2567, n3145);
  not g5400 (n_2568, n3146);
  and g5401 (n3147, n_2567, n_2568);
  and g5402 (n3148, n_2388, n_2394);
  and g5403 (n3149, n3147, n3148);
  not g5404 (n_2569, n3147);
  not g5405 (n_2570, n3148);
  and g5406 (n3150, n_2569, n_2570);
  not g5407 (n_2571, n3149);
  not g5408 (n_2572, n3150);
  and g5409 (n3151, n_2571, n_2572);
  and g5410 (n3152, \b[22] , n511);
  and g5411 (n3153, \b[20] , n541);
  and g5412 (n3154, \b[21] , n506);
  and g5418 (n3157, n514, n2145);
  not g5421 (n_2577, n3158);
  and g5422 (n3159, \a[8] , n_2577);
  not g5423 (n_2578, n3159);
  and g5424 (n3160, \a[8] , n_2578);
  and g5425 (n3161, n_2577, n_2578);
  not g5426 (n_2579, n3160);
  not g5427 (n_2580, n3161);
  and g5428 (n3162, n_2579, n_2580);
  not g5429 (n_2581, n3151);
  and g5430 (n3163, n_2581, n3162);
  not g5431 (n_2582, n3162);
  and g5432 (n3164, n3151, n_2582);
  not g5433 (n_2583, n3163);
  not g5434 (n_2584, n3164);
  and g5435 (n3165, n_2583, n_2584);
  and g5436 (n3166, n_2406, n_2409);
  not g5437 (n_2585, n3166);
  and g5438 (n3167, n3165, n_2585);
  not g5439 (n_2586, n3165);
  and g5440 (n3168, n_2586, n3166);
  not g5441 (n_2587, n3167);
  not g5442 (n_2588, n3168);
  and g5443 (n3169, n_2587, n_2588);
  not g5444 (n_2589, n3014);
  and g5445 (n3170, n_2589, n3169);
  not g5446 (n_2590, n3170);
  and g5447 (n3171, n3169, n_2590);
  and g5448 (n3172, n_2589, n_2590);
  not g5449 (n_2591, n3171);
  not g5450 (n_2592, n3172);
  and g5451 (n3173, n_2591, n_2592);
  and g5452 (n3174, n_2412, n_2419);
  and g5453 (n3175, n3173, n3174);
  not g5454 (n_2593, n3173);
  not g5455 (n_2594, n3174);
  and g5456 (n3176, n_2593, n_2594);
  not g5457 (n_2595, n3175);
  not g5458 (n_2596, n3176);
  and g5459 (n3177, n_2595, n_2596);
  and g5460 (n3178, \b[28] , n266);
  and g5461 (n3179, \b[26] , n284);
  and g5462 (n3180, \b[27] , n261);
  and g5468 (n3183, n_2426, n_2429);
  not g5469 (n_2601, \b[28] );
  and g5470 (n3184, n_2424, n_2601);
  and g5471 (n3185, \b[27] , \b[28] );
  not g5472 (n_2602, n3184);
  not g5473 (n_2603, n3185);
  and g5474 (n3186, n_2602, n_2603);
  not g5475 (n_2604, n3183);
  and g5476 (n3187, n_2604, n3186);
  not g5477 (n_2605, n3186);
  and g5478 (n3188, n3183, n_2605);
  not g5479 (n_2606, n3187);
  not g5480 (n_2607, n3188);
  and g5481 (n3189, n_2606, n_2607);
  and g5482 (n3190, n269, n3189);
  not g5485 (n_2609, n3191);
  and g5486 (n3192, \a[2] , n_2609);
  not g5487 (n_2610, n3192);
  and g5488 (n3193, \a[2] , n_2610);
  and g5489 (n3194, n_2609, n_2610);
  not g5490 (n_2611, n3193);
  not g5491 (n_2612, n3194);
  and g5492 (n3195, n_2611, n_2612);
  not g5493 (n_2613, n3177);
  and g5494 (n3196, n_2613, n3195);
  not g5495 (n_2614, n3195);
  and g5496 (n3197, n3177, n_2614);
  not g5497 (n_2615, n3196);
  not g5498 (n_2616, n3197);
  and g5499 (n3198, n_2615, n_2616);
  not g5500 (n_2617, n3003);
  and g5501 (n3199, n_2617, n3198);
  not g5502 (n_2618, n3198);
  and g5503 (n3200, n3003, n_2618);
  not g5504 (n_2619, n3199);
  not g5505 (n_2620, n3200);
  and g5506 (\f[28] , n_2619, n_2620);
  and g5507 (n3202, n_2590, n_2596);
  and g5508 (n3203, \b[26] , n362);
  and g5509 (n3204, \b[24] , n403);
  and g5510 (n3205, \b[25] , n357);
  and g5516 (n3208, n365, n2813);
  not g5519 (n_2625, n3209);
  and g5520 (n3210, \a[5] , n_2625);
  not g5521 (n_2626, n3210);
  and g5522 (n3211, \a[5] , n_2626);
  and g5523 (n3212, n_2625, n_2626);
  not g5524 (n_2627, n3211);
  not g5525 (n_2628, n3212);
  and g5526 (n3213, n_2627, n_2628);
  and g5527 (n3214, n_2566, n_2572);
  and g5528 (n3215, \b[14] , n1302);
  and g5529 (n3216, \b[12] , n1391);
  and g5530 (n3217, \b[13] , n1297);
  and g5536 (n3220, n1034, n1305);
  not g5539 (n_2633, n3221);
  and g5540 (n3222, \a[17] , n_2633);
  not g5541 (n_2634, n3222);
  and g5542 (n3223, \a[17] , n_2634);
  and g5543 (n3224, n_2633, n_2634);
  not g5544 (n_2635, n3223);
  not g5545 (n_2636, n3224);
  and g5546 (n3225, n_2635, n_2636);
  and g5547 (n3226, n_2516, n_2522);
  and g5548 (n3227, \b[11] , n1627);
  and g5549 (n3228, \b[9] , n1763);
  and g5550 (n3229, \b[10] , n1622);
  and g5556 (n3232, n818, n1630);
  not g5559 (n_2641, n3233);
  and g5560 (n3234, \a[20] , n_2641);
  not g5561 (n_2642, n3234);
  and g5562 (n3235, \a[20] , n_2642);
  and g5563 (n3236, n_2641, n_2642);
  not g5564 (n_2643, n3235);
  not g5565 (n_2644, n3236);
  and g5566 (n3237, n_2643, n_2644);
  and g5567 (n3238, n_2501, n_2505);
  and g5568 (n3239, n_2491, n3062);
  not g5569 (n_2645, n3239);
  and g5570 (n3240, n_2497, n_2645);
  and g5571 (n3241, \b[2] , n3050);
  and g5572 (n3242, n2875, n_2481);
  and g5573 (n3243, n3044, n3242);
  and g5574 (n3244, \b[0] , n3243);
  and g5575 (n3245, \b[1] , n3045);
  and g5581 (n3248, n296, n3053);
  not g5584 (n_2650, n3249);
  and g5585 (n3250, \a[29] , n_2650);
  not g5586 (n_2651, n3250);
  and g5587 (n3251, \a[29] , n_2651);
  and g5588 (n3252, n_2650, n_2651);
  not g5589 (n_2652, n3251);
  not g5590 (n_2653, n3252);
  and g5591 (n3253, n_2652, n_2653);
  and g5592 (n3254, n_2489, n3253);
  not g5593 (n_2654, n3253);
  and g5594 (n3255, n3060, n_2654);
  not g5595 (n_2655, n3254);
  not g5596 (n_2656, n3255);
  and g5597 (n3256, n_2655, n_2656);
  and g5598 (n3257, \b[5] , n2539);
  and g5599 (n3258, \b[3] , n2685);
  and g5600 (n3259, \b[4] , n2534);
  and g5606 (n3262, n394, n2542);
  not g5609 (n_2661, n3263);
  and g5610 (n3264, \a[26] , n_2661);
  not g5611 (n_2662, n3264);
  and g5612 (n3265, \a[26] , n_2662);
  and g5613 (n3266, n_2661, n_2662);
  not g5614 (n_2663, n3265);
  not g5615 (n_2664, n3266);
  and g5616 (n3267, n_2663, n_2664);
  not g5617 (n_2665, n3267);
  and g5618 (n3268, n3256, n_2665);
  not g5619 (n_2666, n3256);
  and g5620 (n3269, n_2666, n3267);
  not g5621 (n_2667, n3240);
  not g5622 (n_2668, n3269);
  and g5623 (n3270, n_2667, n_2668);
  not g5624 (n_2669, n3268);
  and g5625 (n3271, n_2669, n3270);
  not g5626 (n_2670, n3271);
  and g5627 (n3272, n_2667, n_2670);
  and g5628 (n3273, n_2669, n_2670);
  and g5629 (n3274, n_2668, n3273);
  not g5630 (n_2671, n3272);
  not g5631 (n_2672, n3274);
  and g5632 (n3275, n_2671, n_2672);
  and g5633 (n3276, \b[8] , n2048);
  and g5634 (n3277, \b[6] , n2198);
  and g5635 (n3278, \b[7] , n2043);
  and g5641 (n3281, n585, n2051);
  not g5644 (n_2677, n3282);
  and g5645 (n3283, \a[23] , n_2677);
  not g5646 (n_2678, n3283);
  and g5647 (n3284, \a[23] , n_2678);
  and g5648 (n3285, n_2677, n_2678);
  not g5649 (n_2679, n3284);
  not g5650 (n_2680, n3285);
  and g5651 (n3286, n_2679, n_2680);
  and g5652 (n3287, n3275, n3286);
  not g5653 (n_2681, n3275);
  not g5654 (n_2682, n3286);
  and g5655 (n3288, n_2681, n_2682);
  not g5656 (n_2683, n3287);
  not g5657 (n_2684, n3288);
  and g5658 (n3289, n_2683, n_2684);
  not g5659 (n_2685, n3238);
  and g5660 (n3290, n_2685, n3289);
  not g5661 (n_2686, n3289);
  and g5662 (n3291, n3238, n_2686);
  not g5663 (n_2687, n3290);
  not g5664 (n_2688, n3291);
  and g5665 (n3292, n_2687, n_2688);
  not g5666 (n_2689, n3292);
  and g5667 (n3293, n3237, n_2689);
  not g5668 (n_2690, n3237);
  and g5669 (n3294, n_2690, n3292);
  not g5670 (n_2691, n3293);
  not g5671 (n_2692, n3294);
  and g5672 (n3295, n_2691, n_2692);
  not g5673 (n_2693, n3226);
  and g5674 (n3296, n_2693, n3295);
  not g5675 (n_2694, n3295);
  and g5676 (n3297, n3226, n_2694);
  not g5677 (n_2695, n3296);
  not g5678 (n_2696, n3297);
  and g5679 (n3298, n_2695, n_2696);
  not g5680 (n_2697, n3225);
  and g5681 (n3299, n_2697, n3298);
  not g5682 (n_2698, n3299);
  and g5683 (n3300, n3298, n_2698);
  and g5684 (n3301, n_2697, n_2698);
  not g5685 (n_2699, n3300);
  not g5686 (n_2700, n3301);
  and g5687 (n3302, n_2699, n_2700);
  and g5688 (n3303, n_2532, n_2537);
  and g5689 (n3304, n3302, n3303);
  not g5690 (n_2701, n3302);
  not g5691 (n_2702, n3303);
  and g5692 (n3305, n_2701, n_2702);
  not g5693 (n_2703, n3304);
  not g5694 (n_2704, n3305);
  and g5695 (n3306, n_2703, n_2704);
  and g5696 (n3307, \b[17] , n951);
  and g5697 (n3308, \b[15] , n1056);
  and g5698 (n3309, \b[16] , n946);
  and g5704 (n3312, n954, n1356);
  not g5707 (n_2709, n3313);
  and g5708 (n3314, \a[14] , n_2709);
  not g5709 (n_2710, n3314);
  and g5710 (n3315, \a[14] , n_2710);
  and g5711 (n3316, n_2709, n_2710);
  not g5712 (n_2711, n3315);
  not g5713 (n_2712, n3316);
  and g5714 (n3317, n_2711, n_2712);
  not g5715 (n_2713, n3317);
  and g5716 (n3318, n3306, n_2713);
  not g5717 (n_2714, n3318);
  and g5718 (n3319, n3306, n_2714);
  and g5719 (n3320, n_2713, n_2714);
  not g5720 (n_2715, n3319);
  not g5721 (n_2716, n3320);
  and g5722 (n3321, n_2715, n_2716);
  and g5723 (n3322, n_2550, n_2556);
  and g5724 (n3323, n3321, n3322);
  not g5725 (n_2717, n3321);
  not g5726 (n_2718, n3322);
  and g5727 (n3324, n_2717, n_2718);
  not g5728 (n_2719, n3323);
  not g5729 (n_2720, n3324);
  and g5730 (n3325, n_2719, n_2720);
  and g5731 (n3326, \b[20] , n700);
  and g5732 (n3327, \b[18] , n767);
  and g5733 (n3328, \b[19] , n695);
  and g5739 (n3331, n703, n1846);
  not g5742 (n_2725, n3332);
  and g5743 (n3333, \a[11] , n_2725);
  not g5744 (n_2726, n3333);
  and g5745 (n3334, \a[11] , n_2726);
  and g5746 (n3335, n_2725, n_2726);
  not g5747 (n_2727, n3334);
  not g5748 (n_2728, n3335);
  and g5749 (n3336, n_2727, n_2728);
  not g5750 (n_2729, n3336);
  and g5751 (n3337, n3325, n_2729);
  not g5752 (n_2730, n3325);
  and g5753 (n3338, n_2730, n3336);
  not g5754 (n_2731, n3214);
  not g5755 (n_2732, n3338);
  and g5756 (n3339, n_2731, n_2732);
  not g5757 (n_2733, n3337);
  and g5758 (n3340, n_2733, n3339);
  not g5759 (n_2734, n3340);
  and g5760 (n3341, n_2731, n_2734);
  and g5761 (n3342, n_2733, n_2734);
  and g5762 (n3343, n_2732, n3342);
  not g5763 (n_2735, n3341);
  not g5764 (n_2736, n3343);
  and g5765 (n3344, n_2735, n_2736);
  and g5766 (n3345, \b[23] , n511);
  and g5767 (n3346, \b[21] , n541);
  and g5768 (n3347, \b[22] , n506);
  and g5774 (n3350, n514, n2300);
  not g5777 (n_2741, n3351);
  and g5778 (n3352, \a[8] , n_2741);
  not g5779 (n_2742, n3352);
  and g5780 (n3353, \a[8] , n_2742);
  and g5781 (n3354, n_2741, n_2742);
  not g5782 (n_2743, n3353);
  not g5783 (n_2744, n3354);
  and g5784 (n3355, n_2743, n_2744);
  not g5785 (n_2745, n3344);
  not g5786 (n_2746, n3355);
  and g5787 (n3356, n_2745, n_2746);
  not g5788 (n_2747, n3356);
  and g5789 (n3357, n_2745, n_2747);
  and g5790 (n3358, n_2746, n_2747);
  not g5791 (n_2748, n3357);
  not g5792 (n_2749, n3358);
  and g5793 (n3359, n_2748, n_2749);
  and g5794 (n3360, n_2584, n_2587);
  not g5795 (n_2750, n3359);
  not g5796 (n_2751, n3360);
  and g5797 (n3361, n_2750, n_2751);
  and g5798 (n3362, n3359, n3360);
  not g5799 (n_2752, n3361);
  not g5800 (n_2753, n3362);
  and g5801 (n3363, n_2752, n_2753);
  not g5802 (n_2754, n3213);
  and g5803 (n3364, n_2754, n3363);
  not g5804 (n_2755, n3364);
  and g5805 (n3365, n_2754, n_2755);
  and g5806 (n3366, n3363, n_2755);
  not g5807 (n_2756, n3365);
  not g5808 (n_2757, n3366);
  and g5809 (n3367, n_2756, n_2757);
  not g5810 (n_2758, n3202);
  not g5811 (n_2759, n3367);
  and g5812 (n3368, n_2758, n_2759);
  not g5813 (n_2760, n3368);
  and g5814 (n3369, n_2758, n_2760);
  and g5815 (n3370, n_2759, n_2760);
  not g5816 (n_2761, n3369);
  not g5817 (n_2762, n3370);
  and g5818 (n3371, n_2761, n_2762);
  and g5819 (n3372, \b[29] , n266);
  and g5820 (n3373, \b[27] , n284);
  and g5821 (n3374, \b[28] , n261);
  and g5827 (n3377, n_2603, n_2606);
  not g5828 (n_2767, \b[29] );
  and g5829 (n3378, n_2601, n_2767);
  and g5830 (n3379, \b[28] , \b[29] );
  not g5831 (n_2768, n3378);
  not g5832 (n_2769, n3379);
  and g5833 (n3380, n_2768, n_2769);
  not g5834 (n_2770, n3377);
  and g5835 (n3381, n_2770, n3380);
  not g5836 (n_2771, n3380);
  and g5837 (n3382, n3377, n_2771);
  not g5838 (n_2772, n3381);
  not g5839 (n_2773, n3382);
  and g5840 (n3383, n_2772, n_2773);
  and g5841 (n3384, n269, n3383);
  not g5844 (n_2775, n3385);
  and g5845 (n3386, \a[2] , n_2775);
  not g5846 (n_2776, n3386);
  and g5847 (n3387, \a[2] , n_2776);
  and g5848 (n3388, n_2775, n_2776);
  not g5849 (n_2777, n3387);
  not g5850 (n_2778, n3388);
  and g5851 (n3389, n_2777, n_2778);
  not g5852 (n_2779, n3371);
  not g5853 (n_2780, n3389);
  and g5854 (n3390, n_2779, n_2780);
  not g5855 (n_2781, n3390);
  and g5856 (n3391, n_2779, n_2781);
  and g5857 (n3392, n_2780, n_2781);
  not g5858 (n_2782, n3391);
  not g5859 (n_2783, n3392);
  and g5860 (n3393, n_2782, n_2783);
  and g5861 (n3394, n_2616, n_2619);
  not g5862 (n_2784, n3393);
  not g5863 (n_2785, n3394);
  and g5864 (n3395, n_2784, n_2785);
  and g5865 (n3396, n3393, n3394);
  not g5866 (n_2786, n3395);
  not g5867 (n_2787, n3396);
  and g5868 (\f[29] , n_2786, n_2787);
  and g5869 (n3398, n_2747, n_2752);
  and g5870 (n3399, \b[15] , n1302);
  and g5871 (n3400, \b[13] , n1391);
  and g5872 (n3401, \b[14] , n1297);
  and g5878 (n3404, n1131, n1305);
  not g5881 (n_2792, n3405);
  and g5882 (n3406, \a[17] , n_2792);
  not g5883 (n_2793, n3406);
  and g5884 (n3407, \a[17] , n_2793);
  and g5885 (n3408, n_2792, n_2793);
  not g5886 (n_2794, n3407);
  not g5887 (n_2795, n3408);
  and g5888 (n3409, n_2794, n_2795);
  and g5889 (n3410, n_2692, n_2695);
  and g5890 (n3411, \b[12] , n1627);
  and g5891 (n3412, \b[10] , n1763);
  and g5892 (n3413, \b[11] , n1622);
  and g5898 (n3416, n842, n1630);
  not g5901 (n_2800, n3417);
  and g5902 (n3418, \a[20] , n_2800);
  not g5903 (n_2801, n3418);
  and g5904 (n3419, \a[20] , n_2801);
  and g5905 (n3420, n_2800, n_2801);
  not g5906 (n_2802, n3419);
  not g5907 (n_2803, n3420);
  and g5908 (n3421, n_2802, n_2803);
  and g5909 (n3422, n_2684, n_2687);
  and g5910 (n3423, \b[6] , n2539);
  and g5911 (n3424, \b[4] , n2685);
  and g5912 (n3425, \b[5] , n2534);
  and g5918 (n3428, n459, n2542);
  not g5921 (n_2808, n3429);
  and g5922 (n3430, \a[26] , n_2808);
  not g5923 (n_2809, n3430);
  and g5924 (n3431, \a[26] , n_2809);
  and g5925 (n3432, n_2808, n_2809);
  not g5926 (n_2810, n3431);
  not g5927 (n_2811, n3432);
  and g5928 (n3433, n_2810, n_2811);
  not g5929 (n_2813, \a[30] );
  and g5930 (n3434, \a[29] , n_2813);
  and g5931 (n3435, n_2476, \a[30] );
  not g5932 (n_2814, n3434);
  not g5933 (n_2815, n3435);
  and g5934 (n3436, n_2814, n_2815);
  not g5935 (n_2816, n3436);
  and g5936 (n3437, \b[0] , n_2816);
  and g5937 (n3438, n_2656, n3437);
  not g5938 (n_2817, n3437);
  and g5939 (n3439, n3255, n_2817);
  not g5940 (n_2818, n3438);
  not g5941 (n_2819, n3439);
  and g5942 (n3440, n_2818, n_2819);
  and g5943 (n3441, \b[3] , n3050);
  and g5944 (n3442, \b[1] , n3243);
  and g5945 (n3443, \b[2] , n3045);
  and g5951 (n3446, n318, n3053);
  not g5954 (n_2824, n3447);
  and g5955 (n3448, \a[29] , n_2824);
  not g5956 (n_2825, n3448);
  and g5957 (n3449, \a[29] , n_2825);
  and g5958 (n3450, n_2824, n_2825);
  not g5959 (n_2826, n3449);
  not g5960 (n_2827, n3450);
  and g5961 (n3451, n_2826, n_2827);
  not g5962 (n_2828, n3440);
  not g5963 (n_2829, n3451);
  and g5964 (n3452, n_2828, n_2829);
  and g5965 (n3453, n3440, n3451);
  not g5966 (n_2830, n3452);
  not g5967 (n_2831, n3453);
  and g5968 (n3454, n_2830, n_2831);
  not g5969 (n_2832, n3433);
  and g5970 (n3455, n_2832, n3454);
  not g5971 (n_2833, n3455);
  and g5972 (n3456, n3454, n_2833);
  and g5973 (n3457, n_2832, n_2833);
  not g5974 (n_2834, n3456);
  not g5975 (n_2835, n3457);
  and g5976 (n3458, n_2834, n_2835);
  not g5977 (n_2836, n3273);
  and g5978 (n3459, n_2836, n3458);
  not g5979 (n_2837, n3458);
  and g5980 (n3460, n3273, n_2837);
  not g5981 (n_2838, n3459);
  not g5982 (n_2839, n3460);
  and g5983 (n3461, n_2838, n_2839);
  and g5984 (n3462, \b[9] , n2048);
  and g5985 (n3463, \b[7] , n2198);
  and g5986 (n3464, \b[8] , n2043);
  and g5992 (n3467, n651, n2051);
  not g5995 (n_2844, n3468);
  and g5996 (n3469, \a[23] , n_2844);
  not g5997 (n_2845, n3469);
  and g5998 (n3470, \a[23] , n_2845);
  and g5999 (n3471, n_2844, n_2845);
  not g6000 (n_2846, n3470);
  not g6001 (n_2847, n3471);
  and g6002 (n3472, n_2846, n_2847);
  not g6003 (n_2848, n3461);
  not g6004 (n_2849, n3472);
  and g6005 (n3473, n_2848, n_2849);
  and g6006 (n3474, n3461, n3472);
  not g6007 (n_2850, n3473);
  not g6008 (n_2851, n3474);
  and g6009 (n3475, n_2850, n_2851);
  not g6010 (n_2852, n3422);
  and g6011 (n3476, n_2852, n3475);
  not g6012 (n_2853, n3475);
  and g6013 (n3477, n3422, n_2853);
  not g6014 (n_2854, n3476);
  not g6015 (n_2855, n3477);
  and g6016 (n3478, n_2854, n_2855);
  not g6017 (n_2856, n3478);
  and g6018 (n3479, n3421, n_2856);
  not g6019 (n_2857, n3421);
  and g6020 (n3480, n_2857, n3478);
  not g6021 (n_2858, n3479);
  not g6022 (n_2859, n3480);
  and g6023 (n3481, n_2858, n_2859);
  not g6024 (n_2860, n3410);
  and g6025 (n3482, n_2860, n3481);
  not g6026 (n_2861, n3481);
  and g6027 (n3483, n3410, n_2861);
  not g6028 (n_2862, n3482);
  not g6029 (n_2863, n3483);
  and g6030 (n3484, n_2862, n_2863);
  not g6031 (n_2864, n3409);
  and g6032 (n3485, n_2864, n3484);
  not g6033 (n_2865, n3485);
  and g6034 (n3486, n3484, n_2865);
  and g6035 (n3487, n_2864, n_2865);
  not g6036 (n_2866, n3486);
  not g6037 (n_2867, n3487);
  and g6038 (n3488, n_2866, n_2867);
  and g6039 (n3489, n_2698, n_2704);
  and g6040 (n3490, n3488, n3489);
  not g6041 (n_2868, n3488);
  not g6042 (n_2869, n3489);
  and g6043 (n3491, n_2868, n_2869);
  not g6044 (n_2870, n3490);
  not g6045 (n_2871, n3491);
  and g6046 (n3492, n_2870, n_2871);
  and g6047 (n3493, \b[18] , n951);
  and g6048 (n3494, \b[16] , n1056);
  and g6049 (n3495, \b[17] , n946);
  and g6055 (n3498, n954, n1566);
  not g6058 (n_2876, n3499);
  and g6059 (n3500, \a[14] , n_2876);
  not g6060 (n_2877, n3500);
  and g6061 (n3501, \a[14] , n_2877);
  and g6062 (n3502, n_2876, n_2877);
  not g6063 (n_2878, n3501);
  not g6064 (n_2879, n3502);
  and g6065 (n3503, n_2878, n_2879);
  not g6066 (n_2880, n3503);
  and g6067 (n3504, n3492, n_2880);
  not g6068 (n_2881, n3504);
  and g6069 (n3505, n3492, n_2881);
  and g6070 (n3506, n_2880, n_2881);
  not g6071 (n_2882, n3505);
  not g6072 (n_2883, n3506);
  and g6073 (n3507, n_2882, n_2883);
  and g6074 (n3508, n_2714, n_2720);
  and g6075 (n3509, n3507, n3508);
  not g6076 (n_2884, n3507);
  not g6077 (n_2885, n3508);
  and g6078 (n3510, n_2884, n_2885);
  not g6079 (n_2886, n3509);
  not g6080 (n_2887, n3510);
  and g6081 (n3511, n_2886, n_2887);
  and g6082 (n3512, \b[21] , n700);
  and g6083 (n3513, \b[19] , n767);
  and g6084 (n3514, \b[20] , n695);
  and g6090 (n3517, n703, n1984);
  not g6093 (n_2892, n3518);
  and g6094 (n3519, \a[11] , n_2892);
  not g6095 (n_2893, n3519);
  and g6096 (n3520, \a[11] , n_2893);
  and g6097 (n3521, n_2892, n_2893);
  not g6098 (n_2894, n3520);
  not g6099 (n_2895, n3521);
  and g6100 (n3522, n_2894, n_2895);
  not g6101 (n_2896, n3522);
  and g6102 (n3523, n3511, n_2896);
  not g6103 (n_2897, n3523);
  and g6104 (n3524, n3511, n_2897);
  and g6105 (n3525, n_2896, n_2897);
  not g6106 (n_2898, n3524);
  not g6107 (n_2899, n3525);
  and g6108 (n3526, n_2898, n_2899);
  not g6109 (n_2900, n3342);
  and g6110 (n3527, n_2900, n3526);
  not g6111 (n_2901, n3526);
  and g6112 (n3528, n3342, n_2901);
  not g6113 (n_2902, n3527);
  not g6114 (n_2903, n3528);
  and g6115 (n3529, n_2902, n_2903);
  and g6116 (n3530, \b[24] , n511);
  and g6117 (n3531, \b[22] , n541);
  and g6118 (n3532, \b[23] , n506);
  and g6124 (n3535, n514, n2458);
  not g6127 (n_2908, n3536);
  and g6128 (n3537, \a[8] , n_2908);
  not g6129 (n_2909, n3537);
  and g6130 (n3538, \a[8] , n_2909);
  and g6131 (n3539, n_2908, n_2909);
  not g6132 (n_2910, n3538);
  not g6133 (n_2911, n3539);
  and g6134 (n3540, n_2910, n_2911);
  not g6135 (n_2912, n3529);
  not g6136 (n_2913, n3540);
  and g6137 (n3541, n_2912, n_2913);
  and g6138 (n3542, n3529, n3540);
  not g6139 (n_2914, n3541);
  not g6140 (n_2915, n3542);
  and g6141 (n3543, n_2914, n_2915);
  not g6142 (n_2916, n3543);
  and g6143 (n3544, n3398, n_2916);
  not g6144 (n_2917, n3398);
  and g6145 (n3545, n_2917, n3543);
  not g6146 (n_2918, n3544);
  not g6147 (n_2919, n3545);
  and g6148 (n3546, n_2918, n_2919);
  and g6149 (n3547, \b[27] , n362);
  and g6150 (n3548, \b[25] , n403);
  and g6151 (n3549, \b[26] , n357);
  and g6157 (n3552, n365, n2990);
  not g6160 (n_2924, n3553);
  and g6161 (n3554, \a[5] , n_2924);
  not g6162 (n_2925, n3554);
  and g6163 (n3555, \a[5] , n_2925);
  and g6164 (n3556, n_2924, n_2925);
  not g6165 (n_2926, n3555);
  not g6166 (n_2927, n3556);
  and g6167 (n3557, n_2926, n_2927);
  not g6168 (n_2928, n3557);
  and g6169 (n3558, n3546, n_2928);
  not g6170 (n_2929, n3558);
  and g6171 (n3559, n3546, n_2929);
  and g6172 (n3560, n_2928, n_2929);
  not g6173 (n_2930, n3559);
  not g6174 (n_2931, n3560);
  and g6175 (n3561, n_2930, n_2931);
  and g6176 (n3562, n_2755, n_2760);
  and g6177 (n3563, n3561, n3562);
  not g6178 (n_2932, n3561);
  not g6179 (n_2933, n3562);
  and g6180 (n3564, n_2932, n_2933);
  not g6181 (n_2934, n3563);
  not g6182 (n_2935, n3564);
  and g6183 (n3565, n_2934, n_2935);
  and g6184 (n3566, \b[30] , n266);
  and g6185 (n3567, \b[28] , n284);
  and g6186 (n3568, \b[29] , n261);
  and g6192 (n3571, n_2769, n_2772);
  not g6193 (n_2940, \b[30] );
  and g6194 (n3572, n_2767, n_2940);
  and g6195 (n3573, \b[29] , \b[30] );
  not g6196 (n_2941, n3572);
  not g6197 (n_2942, n3573);
  and g6198 (n3574, n_2941, n_2942);
  not g6199 (n_2943, n3571);
  and g6200 (n3575, n_2943, n3574);
  not g6201 (n_2944, n3574);
  and g6202 (n3576, n3571, n_2944);
  not g6203 (n_2945, n3575);
  not g6204 (n_2946, n3576);
  and g6205 (n3577, n_2945, n_2946);
  and g6206 (n3578, n269, n3577);
  not g6209 (n_2948, n3579);
  and g6210 (n3580, \a[2] , n_2948);
  not g6211 (n_2949, n3580);
  and g6212 (n3581, \a[2] , n_2949);
  and g6213 (n3582, n_2948, n_2949);
  not g6214 (n_2950, n3581);
  not g6215 (n_2951, n3582);
  and g6216 (n3583, n_2950, n_2951);
  not g6217 (n_2952, n3583);
  and g6218 (n3584, n3565, n_2952);
  not g6219 (n_2953, n3584);
  and g6220 (n3585, n3565, n_2953);
  and g6221 (n3586, n_2952, n_2953);
  not g6222 (n_2954, n3585);
  not g6223 (n_2955, n3586);
  and g6224 (n3587, n_2954, n_2955);
  and g6225 (n3588, n_2781, n_2786);
  not g6226 (n_2956, n3587);
  not g6227 (n_2957, n3588);
  and g6228 (n3589, n_2956, n_2957);
  and g6229 (n3590, n3587, n3588);
  not g6230 (n_2958, n3589);
  not g6231 (n_2959, n3590);
  and g6232 (\f[30] , n_2958, n_2959);
  and g6233 (n3592, \b[16] , n1302);
  and g6234 (n3593, \b[14] , n1391);
  and g6235 (n3594, \b[15] , n1297);
  and g6241 (n3597, n1237, n1305);
  not g6244 (n_2964, n3598);
  and g6245 (n3599, \a[17] , n_2964);
  not g6246 (n_2965, n3599);
  and g6247 (n3600, \a[17] , n_2965);
  and g6248 (n3601, n_2964, n_2965);
  not g6249 (n_2966, n3600);
  not g6250 (n_2967, n3601);
  and g6251 (n3602, n_2966, n_2967);
  and g6252 (n3603, n_2836, n_2837);
  not g6253 (n_2968, n3603);
  and g6254 (n3604, n_2833, n_2968);
  and g6255 (n3605, \b[7] , n2539);
  and g6256 (n3606, \b[5] , n2685);
  and g6257 (n3607, \b[6] , n2534);
  and g6263 (n3610, n484, n2542);
  not g6266 (n_2973, n3611);
  and g6267 (n3612, \a[26] , n_2973);
  not g6268 (n_2974, n3612);
  and g6269 (n3613, \a[26] , n_2974);
  and g6270 (n3614, n_2973, n_2974);
  not g6271 (n_2975, n3613);
  not g6272 (n_2976, n3614);
  and g6273 (n3615, n_2975, n_2976);
  and g6274 (n3616, n3255, n3437);
  not g6275 (n_2977, n3616);
  and g6276 (n3617, n_2830, n_2977);
  and g6277 (n3618, \b[4] , n3050);
  and g6278 (n3619, \b[2] , n3243);
  and g6279 (n3620, \b[3] , n3045);
  and g6285 (n3623, n346, n3053);
  not g6288 (n_2982, n3624);
  and g6289 (n3625, \a[29] , n_2982);
  not g6290 (n_2983, n3625);
  and g6291 (n3626, \a[29] , n_2983);
  and g6292 (n3627, n_2982, n_2983);
  not g6293 (n_2984, n3626);
  not g6294 (n_2985, n3627);
  and g6295 (n3628, n_2984, n_2985);
  and g6296 (n3629, \a[32] , n_2817);
  and g6297 (n3630, n_2813, \a[31] );
  not g6298 (n_2988, \a[31] );
  and g6299 (n3631, \a[30] , n_2988);
  not g6300 (n_2989, n3630);
  not g6301 (n_2990, n3631);
  and g6302 (n3632, n_2989, n_2990);
  not g6303 (n_2991, n3632);
  and g6304 (n3633, n3436, n_2991);
  and g6305 (n3634, \b[0] , n3633);
  and g6306 (n3635, n_2988, \a[32] );
  not g6307 (n_2992, \a[32] );
  and g6308 (n3636, \a[31] , n_2992);
  not g6309 (n_2993, n3635);
  not g6310 (n_2994, n3636);
  and g6311 (n3637, n_2993, n_2994);
  and g6312 (n3638, n_2816, n3637);
  and g6313 (n3639, \b[1] , n3638);
  not g6314 (n_2995, n3634);
  not g6315 (n_2996, n3639);
  and g6316 (n3640, n_2995, n_2996);
  not g6317 (n_2997, n3637);
  and g6318 (n3641, n_2816, n_2997);
  and g6319 (n3642, n_21, n3641);
  not g6320 (n_2998, n3642);
  and g6321 (n3643, n3640, n_2998);
  not g6322 (n_2999, n3643);
  and g6323 (n3644, \a[32] , n_2999);
  not g6324 (n_3000, n3644);
  and g6325 (n3645, \a[32] , n_3000);
  and g6326 (n3646, n_2999, n_3000);
  not g6327 (n_3001, n3645);
  not g6328 (n_3002, n3646);
  and g6329 (n3647, n_3001, n_3002);
  not g6330 (n_3003, n3647);
  and g6331 (n3648, n3629, n_3003);
  not g6332 (n_3004, n3629);
  and g6333 (n3649, n_3004, n3647);
  not g6334 (n_3005, n3648);
  not g6335 (n_3006, n3649);
  and g6336 (n3650, n_3005, n_3006);
  and g6337 (n3651, n3628, n3650);
  not g6338 (n_3007, n3628);
  not g6339 (n_3008, n3650);
  and g6340 (n3652, n_3007, n_3008);
  not g6341 (n_3009, n3651);
  not g6342 (n_3010, n3652);
  and g6343 (n3653, n_3009, n_3010);
  not g6344 (n_3011, n3617);
  not g6345 (n_3012, n3653);
  and g6346 (n3654, n_3011, n_3012);
  and g6347 (n3655, n3617, n3653);
  not g6348 (n_3013, n3654);
  not g6349 (n_3014, n3655);
  and g6350 (n3656, n_3013, n_3014);
  not g6351 (n_3015, n3615);
  and g6352 (n3657, n_3015, n3656);
  not g6353 (n_3016, n3656);
  and g6354 (n3658, n3615, n_3016);
  not g6355 (n_3017, n3657);
  not g6356 (n_3018, n3658);
  and g6357 (n3659, n_3017, n_3018);
  not g6358 (n_3019, n3604);
  and g6359 (n3660, n_3019, n3659);
  not g6360 (n_3020, n3659);
  and g6361 (n3661, n3604, n_3020);
  not g6362 (n_3021, n3660);
  not g6363 (n_3022, n3661);
  and g6364 (n3662, n_3021, n_3022);
  and g6365 (n3663, \b[10] , n2048);
  and g6366 (n3664, \b[8] , n2198);
  and g6367 (n3665, \b[9] , n2043);
  and g6373 (n3668, n738, n2051);
  not g6376 (n_3027, n3669);
  and g6377 (n3670, \a[23] , n_3027);
  not g6378 (n_3028, n3670);
  and g6379 (n3671, \a[23] , n_3028);
  and g6380 (n3672, n_3027, n_3028);
  not g6381 (n_3029, n3671);
  not g6382 (n_3030, n3672);
  and g6383 (n3673, n_3029, n_3030);
  not g6384 (n_3031, n3673);
  and g6385 (n3674, n3662, n_3031);
  not g6386 (n_3032, n3674);
  and g6387 (n3675, n3662, n_3032);
  and g6388 (n3676, n_3031, n_3032);
  not g6389 (n_3033, n3675);
  not g6390 (n_3034, n3676);
  and g6391 (n3677, n_3033, n_3034);
  and g6392 (n3678, n_2850, n_2854);
  and g6393 (n3679, n3677, n3678);
  not g6394 (n_3035, n3677);
  not g6395 (n_3036, n3678);
  and g6396 (n3680, n_3035, n_3036);
  not g6397 (n_3037, n3679);
  not g6398 (n_3038, n3680);
  and g6399 (n3681, n_3037, n_3038);
  and g6400 (n3682, \b[13] , n1627);
  and g6401 (n3683, \b[11] , n1763);
  and g6402 (n3684, \b[12] , n1622);
  and g6408 (n3687, n1008, n1630);
  not g6411 (n_3043, n3688);
  and g6412 (n3689, \a[20] , n_3043);
  not g6413 (n_3044, n3689);
  and g6414 (n3690, \a[20] , n_3044);
  and g6415 (n3691, n_3043, n_3044);
  not g6416 (n_3045, n3690);
  not g6417 (n_3046, n3691);
  and g6418 (n3692, n_3045, n_3046);
  not g6419 (n_3047, n3681);
  and g6420 (n3693, n_3047, n3692);
  not g6421 (n_3048, n3692);
  and g6422 (n3694, n3681, n_3048);
  not g6423 (n_3049, n3693);
  not g6424 (n_3050, n3694);
  and g6425 (n3695, n_3049, n_3050);
  and g6426 (n3696, n_2859, n_2862);
  not g6427 (n_3051, n3696);
  and g6428 (n3697, n3695, n_3051);
  not g6429 (n_3052, n3695);
  and g6430 (n3698, n_3052, n3696);
  not g6431 (n_3053, n3697);
  not g6432 (n_3054, n3698);
  and g6433 (n3699, n_3053, n_3054);
  not g6434 (n_3055, n3602);
  and g6435 (n3700, n_3055, n3699);
  not g6436 (n_3056, n3700);
  and g6437 (n3701, n3699, n_3056);
  and g6438 (n3702, n_3055, n_3056);
  not g6439 (n_3057, n3701);
  not g6440 (n_3058, n3702);
  and g6441 (n3703, n_3057, n_3058);
  and g6442 (n3704, n_2865, n_2871);
  and g6443 (n3705, n3703, n3704);
  not g6444 (n_3059, n3703);
  not g6445 (n_3060, n3704);
  and g6446 (n3706, n_3059, n_3060);
  not g6447 (n_3061, n3705);
  not g6448 (n_3062, n3706);
  and g6449 (n3707, n_3061, n_3062);
  and g6450 (n3708, \b[19] , n951);
  and g6451 (n3709, \b[17] , n1056);
  and g6452 (n3710, \b[18] , n946);
  and g6458 (n3713, n954, n1708);
  not g6461 (n_3067, n3714);
  and g6462 (n3715, \a[14] , n_3067);
  not g6463 (n_3068, n3715);
  and g6464 (n3716, \a[14] , n_3068);
  and g6465 (n3717, n_3067, n_3068);
  not g6466 (n_3069, n3716);
  not g6467 (n_3070, n3717);
  and g6468 (n3718, n_3069, n_3070);
  not g6469 (n_3071, n3718);
  and g6470 (n3719, n3707, n_3071);
  not g6471 (n_3072, n3719);
  and g6472 (n3720, n3707, n_3072);
  and g6473 (n3721, n_3071, n_3072);
  not g6474 (n_3073, n3720);
  not g6475 (n_3074, n3721);
  and g6476 (n3722, n_3073, n_3074);
  and g6477 (n3723, n_2881, n_2887);
  and g6478 (n3724, n3722, n3723);
  not g6479 (n_3075, n3722);
  not g6480 (n_3076, n3723);
  and g6481 (n3725, n_3075, n_3076);
  not g6482 (n_3077, n3724);
  not g6483 (n_3078, n3725);
  and g6484 (n3726, n_3077, n_3078);
  and g6485 (n3727, \b[22] , n700);
  and g6486 (n3728, \b[20] , n767);
  and g6487 (n3729, \b[21] , n695);
  and g6493 (n3732, n703, n2145);
  not g6496 (n_3083, n3733);
  and g6497 (n3734, \a[11] , n_3083);
  not g6498 (n_3084, n3734);
  and g6499 (n3735, \a[11] , n_3084);
  and g6500 (n3736, n_3083, n_3084);
  not g6501 (n_3085, n3735);
  not g6502 (n_3086, n3736);
  and g6503 (n3737, n_3085, n_3086);
  not g6504 (n_3087, n3737);
  and g6505 (n3738, n3726, n_3087);
  not g6506 (n_3088, n3738);
  and g6507 (n3739, n3726, n_3088);
  and g6508 (n3740, n_3087, n_3088);
  not g6509 (n_3089, n3739);
  not g6510 (n_3090, n3740);
  and g6511 (n3741, n_3089, n_3090);
  and g6512 (n3742, n_2900, n_2901);
  not g6513 (n_3091, n3742);
  and g6514 (n3743, n_2897, n_3091);
  and g6515 (n3744, n3741, n3743);
  not g6516 (n_3092, n3741);
  not g6517 (n_3093, n3743);
  and g6518 (n3745, n_3092, n_3093);
  not g6519 (n_3094, n3744);
  not g6520 (n_3095, n3745);
  and g6521 (n3746, n_3094, n_3095);
  and g6522 (n3747, \b[25] , n511);
  and g6523 (n3748, \b[23] , n541);
  and g6524 (n3749, \b[24] , n506);
  and g6530 (n3752, n514, n2485);
  not g6533 (n_3100, n3753);
  and g6534 (n3754, \a[8] , n_3100);
  not g6535 (n_3101, n3754);
  and g6536 (n3755, \a[8] , n_3101);
  and g6537 (n3756, n_3100, n_3101);
  not g6538 (n_3102, n3755);
  not g6539 (n_3103, n3756);
  and g6540 (n3757, n_3102, n_3103);
  not g6541 (n_3104, n3757);
  and g6542 (n3758, n3746, n_3104);
  not g6543 (n_3105, n3758);
  and g6544 (n3759, n3746, n_3105);
  and g6545 (n3760, n_3104, n_3105);
  not g6546 (n_3106, n3759);
  not g6547 (n_3107, n3760);
  and g6548 (n3761, n_3106, n_3107);
  and g6549 (n3762, n_2914, n_2919);
  and g6550 (n3763, n3761, n3762);
  not g6551 (n_3108, n3761);
  not g6552 (n_3109, n3762);
  and g6553 (n3764, n_3108, n_3109);
  not g6554 (n_3110, n3763);
  not g6555 (n_3111, n3764);
  and g6556 (n3765, n_3110, n_3111);
  and g6557 (n3766, \b[28] , n362);
  and g6558 (n3767, \b[26] , n403);
  and g6559 (n3768, \b[27] , n357);
  and g6565 (n3771, n365, n3189);
  not g6568 (n_3116, n3772);
  and g6569 (n3773, \a[5] , n_3116);
  not g6570 (n_3117, n3773);
  and g6571 (n3774, \a[5] , n_3117);
  and g6572 (n3775, n_3116, n_3117);
  not g6573 (n_3118, n3774);
  not g6574 (n_3119, n3775);
  and g6575 (n3776, n_3118, n_3119);
  not g6576 (n_3120, n3776);
  and g6577 (n3777, n3765, n_3120);
  not g6578 (n_3121, n3777);
  and g6579 (n3778, n3765, n_3121);
  and g6580 (n3779, n_3120, n_3121);
  not g6581 (n_3122, n3778);
  not g6582 (n_3123, n3779);
  and g6583 (n3780, n_3122, n_3123);
  and g6584 (n3781, n_2929, n_2935);
  and g6585 (n3782, n3780, n3781);
  not g6586 (n_3124, n3780);
  not g6587 (n_3125, n3781);
  and g6588 (n3783, n_3124, n_3125);
  not g6589 (n_3126, n3782);
  not g6590 (n_3127, n3783);
  and g6591 (n3784, n_3126, n_3127);
  and g6592 (n3785, \b[31] , n266);
  and g6593 (n3786, \b[29] , n284);
  and g6594 (n3787, \b[30] , n261);
  and g6600 (n3790, n_2942, n_2945);
  not g6601 (n_3132, \b[31] );
  and g6602 (n3791, n_2940, n_3132);
  and g6603 (n3792, \b[30] , \b[31] );
  not g6604 (n_3133, n3791);
  not g6605 (n_3134, n3792);
  and g6606 (n3793, n_3133, n_3134);
  not g6607 (n_3135, n3790);
  and g6608 (n3794, n_3135, n3793);
  not g6609 (n_3136, n3793);
  and g6610 (n3795, n3790, n_3136);
  not g6611 (n_3137, n3794);
  not g6612 (n_3138, n3795);
  and g6613 (n3796, n_3137, n_3138);
  and g6614 (n3797, n269, n3796);
  not g6617 (n_3140, n3798);
  and g6618 (n3799, \a[2] , n_3140);
  not g6619 (n_3141, n3799);
  and g6620 (n3800, \a[2] , n_3141);
  and g6621 (n3801, n_3140, n_3141);
  not g6622 (n_3142, n3800);
  not g6623 (n_3143, n3801);
  and g6624 (n3802, n_3142, n_3143);
  not g6625 (n_3144, n3802);
  and g6626 (n3803, n3784, n_3144);
  not g6627 (n_3145, n3803);
  and g6628 (n3804, n3784, n_3145);
  and g6629 (n3805, n_3144, n_3145);
  not g6630 (n_3146, n3804);
  not g6631 (n_3147, n3805);
  and g6632 (n3806, n_3146, n_3147);
  and g6633 (n3807, n_2953, n_2958);
  not g6634 (n_3148, n3806);
  not g6635 (n_3149, n3807);
  and g6636 (n3808, n_3148, n_3149);
  and g6637 (n3809, n3806, n3807);
  not g6638 (n_3150, n3808);
  not g6639 (n_3151, n3809);
  and g6640 (\f[31] , n_3150, n_3151);
  and g6641 (n3811, n_3145, n_3150);
  and g6642 (n3812, n_3121, n_3127);
  and g6643 (n3813, \b[26] , n511);
  and g6644 (n3814, \b[24] , n541);
  and g6645 (n3815, \b[25] , n506);
  and g6651 (n3818, n514, n2813);
  not g6654 (n_3156, n3819);
  and g6655 (n3820, \a[8] , n_3156);
  not g6656 (n_3157, n3820);
  and g6657 (n3821, \a[8] , n_3157);
  and g6658 (n3822, n_3156, n_3157);
  not g6659 (n_3158, n3821);
  not g6660 (n_3159, n3822);
  and g6661 (n3823, n_3158, n_3159);
  and g6662 (n3824, n_3088, n_3095);
  and g6663 (n3825, n_3072, n_3078);
  and g6664 (n3826, \b[17] , n1302);
  and g6665 (n3827, \b[15] , n1391);
  and g6666 (n3828, \b[16] , n1297);
  and g6672 (n3831, n1305, n1356);
  not g6675 (n_3164, n3832);
  and g6676 (n3833, \a[17] , n_3164);
  not g6677 (n_3165, n3833);
  and g6678 (n3834, \a[17] , n_3165);
  and g6679 (n3835, n_3164, n_3165);
  not g6680 (n_3166, n3834);
  not g6681 (n_3167, n3835);
  and g6682 (n3836, n_3166, n_3167);
  and g6683 (n3837, n_3050, n_3053);
  and g6684 (n3838, n_3032, n_3038);
  and g6685 (n3839, n_3007, n3650);
  not g6686 (n_3168, n3839);
  and g6687 (n3840, n_3013, n_3168);
  and g6688 (n3841, \b[2] , n3638);
  and g6689 (n3842, n3436, n_2997);
  and g6690 (n3843, n3632, n3842);
  and g6691 (n3844, \b[0] , n3843);
  and g6692 (n3845, \b[1] , n3633);
  and g6698 (n3848, n296, n3641);
  not g6701 (n_3173, n3849);
  and g6702 (n3850, \a[32] , n_3173);
  not g6703 (n_3174, n3850);
  and g6704 (n3851, \a[32] , n_3174);
  and g6705 (n3852, n_3173, n_3174);
  not g6706 (n_3175, n3851);
  not g6707 (n_3176, n3852);
  and g6708 (n3853, n_3175, n_3176);
  and g6709 (n3854, n_3005, n3853);
  not g6710 (n_3177, n3853);
  and g6711 (n3855, n3648, n_3177);
  not g6712 (n_3178, n3854);
  not g6713 (n_3179, n3855);
  and g6714 (n3856, n_3178, n_3179);
  and g6715 (n3857, \b[5] , n3050);
  and g6716 (n3858, \b[3] , n3243);
  and g6717 (n3859, \b[4] , n3045);
  and g6723 (n3862, n394, n3053);
  not g6726 (n_3184, n3863);
  and g6727 (n3864, \a[29] , n_3184);
  not g6728 (n_3185, n3864);
  and g6729 (n3865, \a[29] , n_3185);
  and g6730 (n3866, n_3184, n_3185);
  not g6731 (n_3186, n3865);
  not g6732 (n_3187, n3866);
  and g6733 (n3867, n_3186, n_3187);
  not g6734 (n_3188, n3867);
  and g6735 (n3868, n3856, n_3188);
  not g6736 (n_3189, n3856);
  and g6737 (n3869, n_3189, n3867);
  not g6738 (n_3190, n3840);
  not g6739 (n_3191, n3869);
  and g6740 (n3870, n_3190, n_3191);
  not g6741 (n_3192, n3868);
  and g6742 (n3871, n_3192, n3870);
  not g6743 (n_3193, n3871);
  and g6744 (n3872, n_3190, n_3193);
  and g6745 (n3873, n_3192, n_3193);
  and g6746 (n3874, n_3191, n3873);
  not g6747 (n_3194, n3872);
  not g6748 (n_3195, n3874);
  and g6749 (n3875, n_3194, n_3195);
  and g6750 (n3876, \b[8] , n2539);
  and g6751 (n3877, \b[6] , n2685);
  and g6752 (n3878, \b[7] , n2534);
  and g6758 (n3881, n585, n2542);
  not g6761 (n_3200, n3882);
  and g6762 (n3883, \a[26] , n_3200);
  not g6763 (n_3201, n3883);
  and g6764 (n3884, \a[26] , n_3201);
  and g6765 (n3885, n_3200, n_3201);
  not g6766 (n_3202, n3884);
  not g6767 (n_3203, n3885);
  and g6768 (n3886, n_3202, n_3203);
  not g6769 (n_3204, n3875);
  not g6770 (n_3205, n3886);
  and g6771 (n3887, n_3204, n_3205);
  not g6772 (n_3206, n3887);
  and g6773 (n3888, n_3204, n_3206);
  and g6774 (n3889, n_3205, n_3206);
  not g6775 (n_3207, n3888);
  not g6776 (n_3208, n3889);
  and g6777 (n3890, n_3207, n_3208);
  and g6778 (n3891, n_3017, n_3021);
  and g6779 (n3892, n3890, n3891);
  not g6780 (n_3209, n3890);
  not g6781 (n_3210, n3891);
  and g6782 (n3893, n_3209, n_3210);
  not g6783 (n_3211, n3892);
  not g6784 (n_3212, n3893);
  and g6785 (n3894, n_3211, n_3212);
  and g6786 (n3895, \b[11] , n2048);
  and g6787 (n3896, \b[9] , n2198);
  and g6788 (n3897, \b[10] , n2043);
  and g6794 (n3900, n818, n2051);
  not g6797 (n_3217, n3901);
  and g6798 (n3902, \a[23] , n_3217);
  not g6799 (n_3218, n3902);
  and g6800 (n3903, \a[23] , n_3218);
  and g6801 (n3904, n_3217, n_3218);
  not g6802 (n_3219, n3903);
  not g6803 (n_3220, n3904);
  and g6804 (n3905, n_3219, n_3220);
  not g6805 (n_3221, n3905);
  and g6806 (n3906, n3894, n_3221);
  not g6807 (n_3222, n3894);
  and g6808 (n3907, n_3222, n3905);
  not g6809 (n_3223, n3838);
  not g6810 (n_3224, n3907);
  and g6811 (n3908, n_3223, n_3224);
  not g6812 (n_3225, n3906);
  and g6813 (n3909, n_3225, n3908);
  not g6814 (n_3226, n3909);
  and g6815 (n3910, n_3223, n_3226);
  and g6816 (n3911, n_3225, n_3226);
  and g6817 (n3912, n_3224, n3911);
  not g6818 (n_3227, n3910);
  not g6819 (n_3228, n3912);
  and g6820 (n3913, n_3227, n_3228);
  and g6821 (n3914, \b[14] , n1627);
  and g6822 (n3915, \b[12] , n1763);
  and g6823 (n3916, \b[13] , n1622);
  and g6829 (n3919, n1034, n1630);
  not g6832 (n_3233, n3920);
  and g6833 (n3921, \a[20] , n_3233);
  not g6834 (n_3234, n3921);
  and g6835 (n3922, \a[20] , n_3234);
  and g6836 (n3923, n_3233, n_3234);
  not g6837 (n_3235, n3922);
  not g6838 (n_3236, n3923);
  and g6839 (n3924, n_3235, n_3236);
  and g6840 (n3925, n3913, n3924);
  not g6841 (n_3237, n3913);
  not g6842 (n_3238, n3924);
  and g6843 (n3926, n_3237, n_3238);
  not g6844 (n_3239, n3925);
  not g6845 (n_3240, n3926);
  and g6846 (n3927, n_3239, n_3240);
  not g6847 (n_3241, n3837);
  and g6848 (n3928, n_3241, n3927);
  not g6849 (n_3242, n3927);
  and g6850 (n3929, n3837, n_3242);
  not g6851 (n_3243, n3928);
  not g6852 (n_3244, n3929);
  and g6853 (n3930, n_3243, n_3244);
  not g6854 (n_3245, n3836);
  and g6855 (n3931, n_3245, n3930);
  not g6856 (n_3246, n3931);
  and g6857 (n3932, n3930, n_3246);
  and g6858 (n3933, n_3245, n_3246);
  not g6859 (n_3247, n3932);
  not g6860 (n_3248, n3933);
  and g6861 (n3934, n_3247, n_3248);
  and g6862 (n3935, n_3056, n_3062);
  and g6863 (n3936, n3934, n3935);
  not g6864 (n_3249, n3934);
  not g6865 (n_3250, n3935);
  and g6866 (n3937, n_3249, n_3250);
  not g6867 (n_3251, n3936);
  not g6868 (n_3252, n3937);
  and g6869 (n3938, n_3251, n_3252);
  and g6870 (n3939, \b[20] , n951);
  and g6871 (n3940, \b[18] , n1056);
  and g6872 (n3941, \b[19] , n946);
  and g6878 (n3944, n954, n1846);
  not g6881 (n_3257, n3945);
  and g6882 (n3946, \a[14] , n_3257);
  not g6883 (n_3258, n3946);
  and g6884 (n3947, \a[14] , n_3258);
  and g6885 (n3948, n_3257, n_3258);
  not g6886 (n_3259, n3947);
  not g6887 (n_3260, n3948);
  and g6888 (n3949, n_3259, n_3260);
  not g6889 (n_3261, n3949);
  and g6890 (n3950, n3938, n_3261);
  not g6891 (n_3262, n3938);
  and g6892 (n3951, n_3262, n3949);
  not g6893 (n_3263, n3825);
  not g6894 (n_3264, n3951);
  and g6895 (n3952, n_3263, n_3264);
  not g6896 (n_3265, n3950);
  and g6897 (n3953, n_3265, n3952);
  not g6898 (n_3266, n3953);
  and g6899 (n3954, n_3263, n_3266);
  and g6900 (n3955, n_3265, n_3266);
  and g6901 (n3956, n_3264, n3955);
  not g6902 (n_3267, n3954);
  not g6903 (n_3268, n3956);
  and g6904 (n3957, n_3267, n_3268);
  and g6905 (n3958, \b[23] , n700);
  and g6906 (n3959, \b[21] , n767);
  and g6907 (n3960, \b[22] , n695);
  and g6913 (n3963, n703, n2300);
  not g6916 (n_3273, n3964);
  and g6917 (n3965, \a[11] , n_3273);
  not g6918 (n_3274, n3965);
  and g6919 (n3966, \a[11] , n_3274);
  and g6920 (n3967, n_3273, n_3274);
  not g6921 (n_3275, n3966);
  not g6922 (n_3276, n3967);
  and g6923 (n3968, n_3275, n_3276);
  and g6924 (n3969, n3957, n3968);
  not g6925 (n_3277, n3957);
  not g6926 (n_3278, n3968);
  and g6927 (n3970, n_3277, n_3278);
  not g6928 (n_3279, n3969);
  not g6929 (n_3280, n3970);
  and g6930 (n3971, n_3279, n_3280);
  not g6931 (n_3281, n3824);
  and g6932 (n3972, n_3281, n3971);
  not g6933 (n_3282, n3971);
  and g6934 (n3973, n3824, n_3282);
  not g6935 (n_3283, n3972);
  not g6936 (n_3284, n3973);
  and g6937 (n3974, n_3283, n_3284);
  not g6938 (n_3285, n3823);
  and g6939 (n3975, n_3285, n3974);
  not g6940 (n_3286, n3975);
  and g6941 (n3976, n3974, n_3286);
  and g6942 (n3977, n_3285, n_3286);
  not g6943 (n_3287, n3976);
  not g6944 (n_3288, n3977);
  and g6945 (n3978, n_3287, n_3288);
  and g6946 (n3979, n_3105, n_3111);
  and g6947 (n3980, n3978, n3979);
  not g6948 (n_3289, n3978);
  not g6949 (n_3290, n3979);
  and g6950 (n3981, n_3289, n_3290);
  not g6951 (n_3291, n3980);
  not g6952 (n_3292, n3981);
  and g6953 (n3982, n_3291, n_3292);
  and g6954 (n3983, \b[29] , n362);
  and g6955 (n3984, \b[27] , n403);
  and g6956 (n3985, \b[28] , n357);
  and g6962 (n3988, n365, n3383);
  not g6965 (n_3297, n3989);
  and g6966 (n3990, \a[5] , n_3297);
  not g6967 (n_3298, n3990);
  and g6968 (n3991, \a[5] , n_3298);
  and g6969 (n3992, n_3297, n_3298);
  not g6970 (n_3299, n3991);
  not g6971 (n_3300, n3992);
  and g6972 (n3993, n_3299, n_3300);
  not g6973 (n_3301, n3993);
  and g6974 (n3994, n3982, n_3301);
  not g6975 (n_3302, n3982);
  and g6976 (n3995, n_3302, n3993);
  not g6977 (n_3303, n3812);
  not g6978 (n_3304, n3995);
  and g6979 (n3996, n_3303, n_3304);
  not g6980 (n_3305, n3994);
  and g6981 (n3997, n_3305, n3996);
  not g6982 (n_3306, n3997);
  and g6983 (n3998, n_3303, n_3306);
  and g6984 (n3999, n_3305, n_3306);
  and g6985 (n4000, n_3304, n3999);
  not g6986 (n_3307, n3998);
  not g6987 (n_3308, n4000);
  and g6988 (n4001, n_3307, n_3308);
  and g6989 (n4002, \b[32] , n266);
  and g6990 (n4003, \b[30] , n284);
  and g6991 (n4004, \b[31] , n261);
  and g6997 (n4007, n_3134, n_3137);
  not g6998 (n_3313, \b[32] );
  and g6999 (n4008, n_3132, n_3313);
  and g7000 (n4009, \b[31] , \b[32] );
  not g7001 (n_3314, n4008);
  not g7002 (n_3315, n4009);
  and g7003 (n4010, n_3314, n_3315);
  not g7004 (n_3316, n4007);
  and g7005 (n4011, n_3316, n4010);
  not g7006 (n_3317, n4010);
  and g7007 (n4012, n4007, n_3317);
  not g7008 (n_3318, n4011);
  not g7009 (n_3319, n4012);
  and g7010 (n4013, n_3318, n_3319);
  and g7011 (n4014, n269, n4013);
  not g7014 (n_3321, n4015);
  and g7015 (n4016, \a[2] , n_3321);
  not g7016 (n_3322, n4016);
  and g7017 (n4017, \a[2] , n_3322);
  and g7018 (n4018, n_3321, n_3322);
  not g7019 (n_3323, n4017);
  not g7020 (n_3324, n4018);
  and g7021 (n4019, n_3323, n_3324);
  not g7022 (n_3325, n4001);
  and g7023 (n4020, n_3325, n4019);
  not g7024 (n_3326, n4019);
  and g7025 (n4021, n4001, n_3326);
  not g7026 (n_3327, n4020);
  not g7027 (n_3328, n4021);
  and g7028 (n4022, n_3327, n_3328);
  not g7029 (n_3329, n3811);
  not g7030 (n_3330, n4022);
  and g7031 (n4023, n_3329, n_3330);
  and g7032 (n4024, n3811, n4022);
  not g7033 (n_3331, n4023);
  not g7034 (n_3332, n4024);
  and g7035 (\f[32] , n_3331, n_3332);
  and g7036 (n4026, n_3325, n_3326);
  not g7037 (n_3333, n4026);
  and g7038 (n4027, n_3331, n_3333);
  and g7039 (n4028, \b[27] , n511);
  and g7040 (n4029, \b[25] , n541);
  and g7041 (n4030, \b[26] , n506);
  and g7047 (n4033, n514, n2990);
  not g7050 (n_3338, n4034);
  and g7051 (n4035, \a[8] , n_3338);
  not g7052 (n_3339, n4035);
  and g7053 (n4036, \a[8] , n_3339);
  and g7054 (n4037, n_3338, n_3339);
  not g7055 (n_3340, n4036);
  not g7056 (n_3341, n4037);
  and g7057 (n4038, n_3340, n_3341);
  and g7058 (n4039, n_3280, n_3283);
  and g7059 (n4040, n_3246, n_3252);
  and g7060 (n4041, n_3240, n_3243);
  and g7061 (n4042, \b[15] , n1627);
  and g7062 (n4043, \b[13] , n1763);
  and g7063 (n4044, \b[14] , n1622);
  and g7069 (n4047, n1131, n1630);
  not g7072 (n_3346, n4048);
  and g7073 (n4049, \a[20] , n_3346);
  not g7074 (n_3347, n4049);
  and g7075 (n4050, \a[20] , n_3347);
  and g7076 (n4051, n_3346, n_3347);
  not g7077 (n_3348, n4050);
  not g7078 (n_3349, n4051);
  and g7079 (n4052, n_3348, n_3349);
  and g7080 (n4053, n_3206, n_3212);
  and g7081 (n4054, \b[6] , n3050);
  and g7082 (n4055, \b[4] , n3243);
  and g7083 (n4056, \b[5] , n3045);
  and g7089 (n4059, n459, n3053);
  not g7092 (n_3354, n4060);
  and g7093 (n4061, \a[29] , n_3354);
  not g7094 (n_3355, n4061);
  and g7095 (n4062, \a[29] , n_3355);
  and g7096 (n4063, n_3354, n_3355);
  not g7097 (n_3356, n4062);
  not g7098 (n_3357, n4063);
  and g7099 (n4064, n_3356, n_3357);
  not g7100 (n_3359, \a[33] );
  and g7101 (n4065, \a[32] , n_3359);
  and g7102 (n4066, n_2992, \a[33] );
  not g7103 (n_3360, n4065);
  not g7104 (n_3361, n4066);
  and g7105 (n4067, n_3360, n_3361);
  not g7106 (n_3362, n4067);
  and g7107 (n4068, \b[0] , n_3362);
  and g7108 (n4069, n_3179, n4068);
  not g7109 (n_3363, n4068);
  and g7110 (n4070, n3855, n_3363);
  not g7111 (n_3364, n4069);
  not g7112 (n_3365, n4070);
  and g7113 (n4071, n_3364, n_3365);
  and g7114 (n4072, \b[3] , n3638);
  and g7115 (n4073, \b[1] , n3843);
  and g7116 (n4074, \b[2] , n3633);
  and g7122 (n4077, n318, n3641);
  not g7125 (n_3370, n4078);
  and g7126 (n4079, \a[32] , n_3370);
  not g7127 (n_3371, n4079);
  and g7128 (n4080, \a[32] , n_3371);
  and g7129 (n4081, n_3370, n_3371);
  not g7130 (n_3372, n4080);
  not g7131 (n_3373, n4081);
  and g7132 (n4082, n_3372, n_3373);
  not g7133 (n_3374, n4071);
  not g7134 (n_3375, n4082);
  and g7135 (n4083, n_3374, n_3375);
  and g7136 (n4084, n4071, n4082);
  not g7137 (n_3376, n4083);
  not g7138 (n_3377, n4084);
  and g7139 (n4085, n_3376, n_3377);
  not g7140 (n_3378, n4064);
  and g7141 (n4086, n_3378, n4085);
  not g7142 (n_3379, n4086);
  and g7143 (n4087, n4085, n_3379);
  and g7144 (n4088, n_3378, n_3379);
  not g7145 (n_3380, n4087);
  not g7146 (n_3381, n4088);
  and g7147 (n4089, n_3380, n_3381);
  not g7148 (n_3382, n3873);
  and g7149 (n4090, n_3382, n4089);
  not g7150 (n_3383, n4089);
  and g7151 (n4091, n3873, n_3383);
  not g7152 (n_3384, n4090);
  not g7153 (n_3385, n4091);
  and g7154 (n4092, n_3384, n_3385);
  and g7155 (n4093, \b[9] , n2539);
  and g7156 (n4094, \b[7] , n2685);
  and g7157 (n4095, \b[8] , n2534);
  and g7163 (n4098, n651, n2542);
  not g7166 (n_3390, n4099);
  and g7167 (n4100, \a[26] , n_3390);
  not g7168 (n_3391, n4100);
  and g7169 (n4101, \a[26] , n_3391);
  and g7170 (n4102, n_3390, n_3391);
  not g7171 (n_3392, n4101);
  not g7172 (n_3393, n4102);
  and g7173 (n4103, n_3392, n_3393);
  not g7174 (n_3394, n4092);
  not g7175 (n_3395, n4103);
  and g7176 (n4104, n_3394, n_3395);
  and g7177 (n4105, n4092, n4103);
  not g7178 (n_3396, n4104);
  not g7179 (n_3397, n4105);
  and g7180 (n4106, n_3396, n_3397);
  not g7181 (n_3398, n4106);
  and g7182 (n4107, n4053, n_3398);
  not g7183 (n_3399, n4053);
  and g7184 (n4108, n_3399, n4106);
  not g7185 (n_3400, n4107);
  not g7186 (n_3401, n4108);
  and g7187 (n4109, n_3400, n_3401);
  and g7188 (n4110, \b[12] , n2048);
  and g7189 (n4111, \b[10] , n2198);
  and g7190 (n4112, \b[11] , n2043);
  and g7196 (n4115, n842, n2051);
  not g7199 (n_3406, n4116);
  and g7200 (n4117, \a[23] , n_3406);
  not g7201 (n_3407, n4117);
  and g7202 (n4118, \a[23] , n_3407);
  and g7203 (n4119, n_3406, n_3407);
  not g7204 (n_3408, n4118);
  not g7205 (n_3409, n4119);
  and g7206 (n4120, n_3408, n_3409);
  not g7207 (n_3410, n4109);
  and g7208 (n4121, n_3410, n4120);
  not g7209 (n_3411, n4120);
  and g7210 (n4122, n4109, n_3411);
  not g7211 (n_3412, n4121);
  not g7212 (n_3413, n4122);
  and g7213 (n4123, n_3412, n_3413);
  not g7214 (n_3414, n3911);
  and g7215 (n4124, n_3414, n4123);
  not g7216 (n_3415, n4123);
  and g7217 (n4125, n3911, n_3415);
  not g7218 (n_3416, n4124);
  not g7219 (n_3417, n4125);
  and g7220 (n4126, n_3416, n_3417);
  not g7221 (n_3418, n4052);
  and g7222 (n4127, n_3418, n4126);
  not g7223 (n_3419, n4127);
  and g7224 (n4128, n4126, n_3419);
  and g7225 (n4129, n_3418, n_3419);
  not g7226 (n_3420, n4128);
  not g7227 (n_3421, n4129);
  and g7228 (n4130, n_3420, n_3421);
  not g7229 (n_3422, n4041);
  and g7230 (n4131, n_3422, n4130);
  not g7231 (n_3423, n4130);
  and g7232 (n4132, n4041, n_3423);
  not g7233 (n_3424, n4131);
  not g7234 (n_3425, n4132);
  and g7235 (n4133, n_3424, n_3425);
  and g7236 (n4134, \b[18] , n1302);
  and g7237 (n4135, \b[16] , n1391);
  and g7238 (n4136, \b[17] , n1297);
  and g7244 (n4139, n1305, n1566);
  not g7247 (n_3430, n4140);
  and g7248 (n4141, \a[17] , n_3430);
  not g7249 (n_3431, n4141);
  and g7250 (n4142, \a[17] , n_3431);
  and g7251 (n4143, n_3430, n_3431);
  not g7252 (n_3432, n4142);
  not g7253 (n_3433, n4143);
  and g7254 (n4144, n_3432, n_3433);
  not g7255 (n_3434, n4133);
  not g7256 (n_3435, n4144);
  and g7257 (n4145, n_3434, n_3435);
  and g7258 (n4146, n4133, n4144);
  not g7259 (n_3436, n4145);
  not g7260 (n_3437, n4146);
  and g7261 (n4147, n_3436, n_3437);
  not g7262 (n_3438, n4147);
  and g7263 (n4148, n4040, n_3438);
  not g7264 (n_3439, n4040);
  and g7265 (n4149, n_3439, n4147);
  not g7266 (n_3440, n4148);
  not g7267 (n_3441, n4149);
  and g7268 (n4150, n_3440, n_3441);
  and g7269 (n4151, \b[21] , n951);
  and g7270 (n4152, \b[19] , n1056);
  and g7271 (n4153, \b[20] , n946);
  and g7277 (n4156, n954, n1984);
  not g7280 (n_3446, n4157);
  and g7281 (n4158, \a[14] , n_3446);
  not g7282 (n_3447, n4158);
  and g7283 (n4159, \a[14] , n_3447);
  and g7284 (n4160, n_3446, n_3447);
  not g7285 (n_3448, n4159);
  not g7286 (n_3449, n4160);
  and g7287 (n4161, n_3448, n_3449);
  not g7288 (n_3450, n4161);
  and g7289 (n4162, n4150, n_3450);
  not g7290 (n_3451, n4162);
  and g7291 (n4163, n4150, n_3451);
  and g7292 (n4164, n_3450, n_3451);
  not g7293 (n_3452, n4163);
  not g7294 (n_3453, n4164);
  and g7295 (n4165, n_3452, n_3453);
  not g7296 (n_3454, n3955);
  and g7297 (n4166, n_3454, n4165);
  not g7298 (n_3455, n4165);
  and g7299 (n4167, n3955, n_3455);
  not g7300 (n_3456, n4166);
  not g7301 (n_3457, n4167);
  and g7302 (n4168, n_3456, n_3457);
  and g7303 (n4169, \b[24] , n700);
  and g7304 (n4170, \b[22] , n767);
  and g7305 (n4171, \b[23] , n695);
  and g7311 (n4174, n703, n2458);
  not g7314 (n_3462, n4175);
  and g7315 (n4176, \a[11] , n_3462);
  not g7316 (n_3463, n4176);
  and g7317 (n4177, \a[11] , n_3463);
  and g7318 (n4178, n_3462, n_3463);
  not g7319 (n_3464, n4177);
  not g7320 (n_3465, n4178);
  and g7321 (n4179, n_3464, n_3465);
  and g7322 (n4180, n4168, n4179);
  not g7323 (n_3466, n4168);
  not g7324 (n_3467, n4179);
  and g7325 (n4181, n_3466, n_3467);
  not g7326 (n_3468, n4180);
  not g7327 (n_3469, n4181);
  and g7328 (n4182, n_3468, n_3469);
  not g7329 (n_3470, n4039);
  and g7330 (n4183, n_3470, n4182);
  not g7331 (n_3471, n4182);
  and g7332 (n4184, n4039, n_3471);
  not g7333 (n_3472, n4183);
  not g7334 (n_3473, n4184);
  and g7335 (n4185, n_3472, n_3473);
  not g7336 (n_3474, n4038);
  and g7337 (n4186, n_3474, n4185);
  not g7338 (n_3475, n4186);
  and g7339 (n4187, n4185, n_3475);
  and g7340 (n4188, n_3474, n_3475);
  not g7341 (n_3476, n4187);
  not g7342 (n_3477, n4188);
  and g7343 (n4189, n_3476, n_3477);
  and g7344 (n4190, n_3286, n_3292);
  and g7345 (n4191, n4189, n4190);
  not g7346 (n_3478, n4189);
  not g7347 (n_3479, n4190);
  and g7348 (n4192, n_3478, n_3479);
  not g7349 (n_3480, n4191);
  not g7350 (n_3481, n4192);
  and g7351 (n4193, n_3480, n_3481);
  and g7352 (n4194, \b[30] , n362);
  and g7353 (n4195, \b[28] , n403);
  and g7354 (n4196, \b[29] , n357);
  and g7360 (n4199, n365, n3577);
  not g7363 (n_3486, n4200);
  and g7364 (n4201, \a[5] , n_3486);
  not g7365 (n_3487, n4201);
  and g7366 (n4202, \a[5] , n_3487);
  and g7367 (n4203, n_3486, n_3487);
  not g7368 (n_3488, n4202);
  not g7369 (n_3489, n4203);
  and g7370 (n4204, n_3488, n_3489);
  not g7371 (n_3490, n4204);
  and g7372 (n4205, n4193, n_3490);
  not g7373 (n_3491, n4205);
  and g7374 (n4206, n4193, n_3491);
  and g7375 (n4207, n_3490, n_3491);
  not g7376 (n_3492, n4206);
  not g7377 (n_3493, n4207);
  and g7378 (n4208, n_3492, n_3493);
  not g7379 (n_3494, n3999);
  and g7380 (n4209, n_3494, n4208);
  not g7381 (n_3495, n4208);
  and g7382 (n4210, n3999, n_3495);
  not g7383 (n_3496, n4209);
  not g7384 (n_3497, n4210);
  and g7385 (n4211, n_3496, n_3497);
  and g7386 (n4212, \b[33] , n266);
  and g7387 (n4213, \b[31] , n284);
  and g7388 (n4214, \b[32] , n261);
  and g7394 (n4217, n_3315, n_3318);
  not g7395 (n_3502, \b[33] );
  and g7396 (n4218, n_3313, n_3502);
  and g7397 (n4219, \b[32] , \b[33] );
  not g7398 (n_3503, n4218);
  not g7399 (n_3504, n4219);
  and g7400 (n4220, n_3503, n_3504);
  not g7401 (n_3505, n4217);
  and g7402 (n4221, n_3505, n4220);
  not g7403 (n_3506, n4220);
  and g7404 (n4222, n4217, n_3506);
  not g7405 (n_3507, n4221);
  not g7406 (n_3508, n4222);
  and g7407 (n4223, n_3507, n_3508);
  and g7408 (n4224, n269, n4223);
  not g7411 (n_3510, n4225);
  and g7412 (n4226, \a[2] , n_3510);
  not g7413 (n_3511, n4226);
  and g7414 (n4227, \a[2] , n_3511);
  and g7415 (n4228, n_3510, n_3511);
  not g7416 (n_3512, n4227);
  not g7417 (n_3513, n4228);
  and g7418 (n4229, n_3512, n_3513);
  not g7419 (n_3514, n4211);
  not g7420 (n_3515, n4229);
  and g7421 (n4230, n_3514, n_3515);
  and g7422 (n4231, n4211, n4229);
  not g7423 (n_3516, n4230);
  not g7424 (n_3517, n4231);
  and g7425 (n4232, n_3516, n_3517);
  not g7426 (n_3518, n4027);
  and g7427 (n4233, n_3518, n4232);
  not g7428 (n_3519, n4232);
  and g7429 (n4234, n4027, n_3519);
  not g7430 (n_3520, n4233);
  not g7431 (n_3521, n4234);
  and g7432 (\f[33] , n_3520, n_3521);
  and g7433 (n4236, n_3516, n_3520);
  and g7434 (n4237, n_3494, n_3495);
  not g7435 (n_3522, n4237);
  and g7436 (n4238, n_3491, n_3522);
  and g7437 (n4239, n_3469, n_3472);
  and g7438 (n4240, n_3413, n_3416);
  and g7439 (n4241, \b[10] , n2539);
  and g7440 (n4242, \b[8] , n2685);
  and g7441 (n4243, \b[9] , n2534);
  and g7447 (n4246, n738, n2542);
  not g7450 (n_3527, n4247);
  and g7451 (n4248, \a[26] , n_3527);
  not g7452 (n_3528, n4248);
  and g7453 (n4249, \a[26] , n_3528);
  and g7454 (n4250, n_3527, n_3528);
  not g7455 (n_3529, n4249);
  not g7456 (n_3530, n4250);
  and g7457 (n4251, n_3529, n_3530);
  and g7458 (n4252, n_3382, n_3383);
  not g7459 (n_3531, n4252);
  and g7460 (n4253, n_3379, n_3531);
  and g7461 (n4254, \b[7] , n3050);
  and g7462 (n4255, \b[5] , n3243);
  and g7463 (n4256, \b[6] , n3045);
  and g7469 (n4259, n484, n3053);
  not g7472 (n_3536, n4260);
  and g7473 (n4261, \a[29] , n_3536);
  not g7474 (n_3537, n4261);
  and g7475 (n4262, \a[29] , n_3537);
  and g7476 (n4263, n_3536, n_3537);
  not g7477 (n_3538, n4262);
  not g7478 (n_3539, n4263);
  and g7479 (n4264, n_3538, n_3539);
  and g7480 (n4265, n3855, n4068);
  not g7481 (n_3540, n4265);
  and g7482 (n4266, n_3376, n_3540);
  and g7483 (n4267, \b[4] , n3638);
  and g7484 (n4268, \b[2] , n3843);
  and g7485 (n4269, \b[3] , n3633);
  and g7491 (n4272, n346, n3641);
  not g7494 (n_3545, n4273);
  and g7495 (n4274, \a[32] , n_3545);
  not g7496 (n_3546, n4274);
  and g7497 (n4275, \a[32] , n_3546);
  and g7498 (n4276, n_3545, n_3546);
  not g7499 (n_3547, n4275);
  not g7500 (n_3548, n4276);
  and g7501 (n4277, n_3547, n_3548);
  and g7502 (n4278, \a[35] , n_3363);
  and g7503 (n4279, n_3359, \a[34] );
  not g7504 (n_3551, \a[34] );
  and g7505 (n4280, \a[33] , n_3551);
  not g7506 (n_3552, n4279);
  not g7507 (n_3553, n4280);
  and g7508 (n4281, n_3552, n_3553);
  not g7509 (n_3554, n4281);
  and g7510 (n4282, n4067, n_3554);
  and g7511 (n4283, \b[0] , n4282);
  and g7512 (n4284, n_3551, \a[35] );
  not g7513 (n_3555, \a[35] );
  and g7514 (n4285, \a[34] , n_3555);
  not g7515 (n_3556, n4284);
  not g7516 (n_3557, n4285);
  and g7517 (n4286, n_3556, n_3557);
  and g7518 (n4287, n_3362, n4286);
  and g7519 (n4288, \b[1] , n4287);
  not g7520 (n_3558, n4283);
  not g7521 (n_3559, n4288);
  and g7522 (n4289, n_3558, n_3559);
  not g7523 (n_3560, n4286);
  and g7524 (n4290, n_3362, n_3560);
  and g7525 (n4291, n_21, n4290);
  not g7526 (n_3561, n4291);
  and g7527 (n4292, n4289, n_3561);
  not g7528 (n_3562, n4292);
  and g7529 (n4293, \a[35] , n_3562);
  not g7530 (n_3563, n4293);
  and g7531 (n4294, \a[35] , n_3563);
  and g7532 (n4295, n_3562, n_3563);
  not g7533 (n_3564, n4294);
  not g7534 (n_3565, n4295);
  and g7535 (n4296, n_3564, n_3565);
  not g7536 (n_3566, n4296);
  and g7537 (n4297, n4278, n_3566);
  not g7538 (n_3567, n4278);
  and g7539 (n4298, n_3567, n4296);
  not g7540 (n_3568, n4297);
  not g7541 (n_3569, n4298);
  and g7542 (n4299, n_3568, n_3569);
  not g7543 (n_3570, n4299);
  and g7544 (n4300, n4277, n_3570);
  not g7545 (n_3571, n4277);
  and g7546 (n4301, n_3571, n4299);
  not g7547 (n_3572, n4300);
  not g7548 (n_3573, n4301);
  and g7549 (n4302, n_3572, n_3573);
  not g7550 (n_3574, n4266);
  and g7551 (n4303, n_3574, n4302);
  not g7552 (n_3575, n4302);
  and g7553 (n4304, n4266, n_3575);
  not g7554 (n_3576, n4303);
  not g7555 (n_3577, n4304);
  and g7556 (n4305, n_3576, n_3577);
  not g7557 (n_3578, n4305);
  and g7558 (n4306, n4264, n_3578);
  not g7559 (n_3579, n4264);
  and g7560 (n4307, n_3579, n4305);
  not g7561 (n_3580, n4306);
  not g7562 (n_3581, n4307);
  and g7563 (n4308, n_3580, n_3581);
  not g7564 (n_3582, n4253);
  and g7565 (n4309, n_3582, n4308);
  not g7566 (n_3583, n4308);
  and g7567 (n4310, n4253, n_3583);
  not g7568 (n_3584, n4309);
  not g7569 (n_3585, n4310);
  and g7570 (n4311, n_3584, n_3585);
  not g7571 (n_3586, n4251);
  and g7572 (n4312, n_3586, n4311);
  not g7573 (n_3587, n4312);
  and g7574 (n4313, n4311, n_3587);
  and g7575 (n4314, n_3586, n_3587);
  not g7576 (n_3588, n4313);
  not g7577 (n_3589, n4314);
  and g7578 (n4315, n_3588, n_3589);
  and g7579 (n4316, n_3396, n_3401);
  and g7580 (n4317, n4315, n4316);
  not g7581 (n_3590, n4315);
  not g7582 (n_3591, n4316);
  and g7583 (n4318, n_3590, n_3591);
  not g7584 (n_3592, n4317);
  not g7585 (n_3593, n4318);
  and g7586 (n4319, n_3592, n_3593);
  and g7587 (n4320, \b[13] , n2048);
  and g7588 (n4321, \b[11] , n2198);
  and g7589 (n4322, \b[12] , n2043);
  and g7595 (n4325, n1008, n2051);
  not g7598 (n_3598, n4326);
  and g7599 (n4327, \a[23] , n_3598);
  not g7600 (n_3599, n4327);
  and g7601 (n4328, \a[23] , n_3599);
  and g7602 (n4329, n_3598, n_3599);
  not g7603 (n_3600, n4328);
  not g7604 (n_3601, n4329);
  and g7605 (n4330, n_3600, n_3601);
  not g7606 (n_3602, n4330);
  and g7607 (n4331, n4319, n_3602);
  not g7608 (n_3603, n4319);
  and g7609 (n4332, n_3603, n4330);
  not g7610 (n_3604, n4240);
  not g7611 (n_3605, n4332);
  and g7612 (n4333, n_3604, n_3605);
  not g7613 (n_3606, n4331);
  and g7614 (n4334, n_3606, n4333);
  not g7615 (n_3607, n4334);
  and g7616 (n4335, n_3604, n_3607);
  and g7617 (n4336, n_3606, n_3607);
  and g7618 (n4337, n_3605, n4336);
  not g7619 (n_3608, n4335);
  not g7620 (n_3609, n4337);
  and g7621 (n4338, n_3608, n_3609);
  and g7622 (n4339, \b[16] , n1627);
  and g7623 (n4340, \b[14] , n1763);
  and g7624 (n4341, \b[15] , n1622);
  and g7630 (n4344, n1237, n1630);
  not g7633 (n_3614, n4345);
  and g7634 (n4346, \a[20] , n_3614);
  not g7635 (n_3615, n4346);
  and g7636 (n4347, \a[20] , n_3615);
  and g7637 (n4348, n_3614, n_3615);
  not g7638 (n_3616, n4347);
  not g7639 (n_3617, n4348);
  and g7640 (n4349, n_3616, n_3617);
  not g7641 (n_3618, n4338);
  not g7642 (n_3619, n4349);
  and g7643 (n4350, n_3618, n_3619);
  not g7644 (n_3620, n4350);
  and g7645 (n4351, n_3618, n_3620);
  and g7646 (n4352, n_3619, n_3620);
  not g7647 (n_3621, n4351);
  not g7648 (n_3622, n4352);
  and g7649 (n4353, n_3621, n_3622);
  and g7650 (n4354, n_3422, n_3423);
  not g7651 (n_3623, n4354);
  and g7652 (n4355, n_3419, n_3623);
  and g7653 (n4356, n4353, n4355);
  not g7654 (n_3624, n4353);
  not g7655 (n_3625, n4355);
  and g7656 (n4357, n_3624, n_3625);
  not g7657 (n_3626, n4356);
  not g7658 (n_3627, n4357);
  and g7659 (n4358, n_3626, n_3627);
  and g7660 (n4359, \b[19] , n1302);
  and g7661 (n4360, \b[17] , n1391);
  and g7662 (n4361, \b[18] , n1297);
  and g7668 (n4364, n1305, n1708);
  not g7671 (n_3632, n4365);
  and g7672 (n4366, \a[17] , n_3632);
  not g7673 (n_3633, n4366);
  and g7674 (n4367, \a[17] , n_3633);
  and g7675 (n4368, n_3632, n_3633);
  not g7676 (n_3634, n4367);
  not g7677 (n_3635, n4368);
  and g7678 (n4369, n_3634, n_3635);
  not g7679 (n_3636, n4369);
  and g7680 (n4370, n4358, n_3636);
  not g7681 (n_3637, n4370);
  and g7682 (n4371, n4358, n_3637);
  and g7683 (n4372, n_3636, n_3637);
  not g7684 (n_3638, n4371);
  not g7685 (n_3639, n4372);
  and g7686 (n4373, n_3638, n_3639);
  and g7687 (n4374, n_3436, n_3441);
  and g7688 (n4375, n4373, n4374);
  not g7689 (n_3640, n4373);
  not g7690 (n_3641, n4374);
  and g7691 (n4376, n_3640, n_3641);
  not g7692 (n_3642, n4375);
  not g7693 (n_3643, n4376);
  and g7694 (n4377, n_3642, n_3643);
  and g7695 (n4378, \b[22] , n951);
  and g7696 (n4379, \b[20] , n1056);
  and g7697 (n4380, \b[21] , n946);
  and g7703 (n4383, n954, n2145);
  not g7706 (n_3648, n4384);
  and g7707 (n4385, \a[14] , n_3648);
  not g7708 (n_3649, n4385);
  and g7709 (n4386, \a[14] , n_3649);
  and g7710 (n4387, n_3648, n_3649);
  not g7711 (n_3650, n4386);
  not g7712 (n_3651, n4387);
  and g7713 (n4388, n_3650, n_3651);
  not g7714 (n_3652, n4388);
  and g7715 (n4389, n4377, n_3652);
  not g7716 (n_3653, n4389);
  and g7717 (n4390, n4377, n_3653);
  and g7718 (n4391, n_3652, n_3653);
  not g7719 (n_3654, n4390);
  not g7720 (n_3655, n4391);
  and g7721 (n4392, n_3654, n_3655);
  and g7722 (n4393, n_3454, n_3455);
  not g7723 (n_3656, n4393);
  and g7724 (n4394, n_3451, n_3656);
  and g7725 (n4395, n4392, n4394);
  not g7726 (n_3657, n4392);
  not g7727 (n_3658, n4394);
  and g7728 (n4396, n_3657, n_3658);
  not g7729 (n_3659, n4395);
  not g7730 (n_3660, n4396);
  and g7731 (n4397, n_3659, n_3660);
  and g7732 (n4398, \b[25] , n700);
  and g7733 (n4399, \b[23] , n767);
  and g7734 (n4400, \b[24] , n695);
  and g7740 (n4403, n703, n2485);
  not g7743 (n_3665, n4404);
  and g7744 (n4405, \a[11] , n_3665);
  not g7745 (n_3666, n4405);
  and g7746 (n4406, \a[11] , n_3666);
  and g7747 (n4407, n_3665, n_3666);
  not g7748 (n_3667, n4406);
  not g7749 (n_3668, n4407);
  and g7750 (n4408, n_3667, n_3668);
  not g7751 (n_3669, n4408);
  and g7752 (n4409, n4397, n_3669);
  not g7753 (n_3670, n4397);
  and g7754 (n4410, n_3670, n4408);
  not g7755 (n_3671, n4239);
  not g7756 (n_3672, n4410);
  and g7757 (n4411, n_3671, n_3672);
  not g7758 (n_3673, n4409);
  and g7759 (n4412, n_3673, n4411);
  not g7760 (n_3674, n4412);
  and g7761 (n4413, n_3671, n_3674);
  and g7762 (n4414, n_3673, n_3674);
  and g7763 (n4415, n_3672, n4414);
  not g7764 (n_3675, n4413);
  not g7765 (n_3676, n4415);
  and g7766 (n4416, n_3675, n_3676);
  and g7767 (n4417, \b[28] , n511);
  and g7768 (n4418, \b[26] , n541);
  and g7769 (n4419, \b[27] , n506);
  and g7775 (n4422, n514, n3189);
  not g7778 (n_3681, n4423);
  and g7779 (n4424, \a[8] , n_3681);
  not g7780 (n_3682, n4424);
  and g7781 (n4425, \a[8] , n_3682);
  and g7782 (n4426, n_3681, n_3682);
  not g7783 (n_3683, n4425);
  not g7784 (n_3684, n4426);
  and g7785 (n4427, n_3683, n_3684);
  not g7786 (n_3685, n4416);
  not g7787 (n_3686, n4427);
  and g7788 (n4428, n_3685, n_3686);
  not g7789 (n_3687, n4428);
  and g7790 (n4429, n_3685, n_3687);
  and g7791 (n4430, n_3686, n_3687);
  not g7792 (n_3688, n4429);
  not g7793 (n_3689, n4430);
  and g7794 (n4431, n_3688, n_3689);
  and g7795 (n4432, n_3475, n_3481);
  and g7796 (n4433, n4431, n4432);
  not g7797 (n_3690, n4431);
  not g7798 (n_3691, n4432);
  and g7799 (n4434, n_3690, n_3691);
  not g7800 (n_3692, n4433);
  not g7801 (n_3693, n4434);
  and g7802 (n4435, n_3692, n_3693);
  and g7803 (n4436, \b[31] , n362);
  and g7804 (n4437, \b[29] , n403);
  and g7805 (n4438, \b[30] , n357);
  and g7811 (n4441, n365, n3796);
  not g7814 (n_3698, n4442);
  and g7815 (n4443, \a[5] , n_3698);
  not g7816 (n_3699, n4443);
  and g7817 (n4444, \a[5] , n_3699);
  and g7818 (n4445, n_3698, n_3699);
  not g7819 (n_3700, n4444);
  not g7820 (n_3701, n4445);
  and g7821 (n4446, n_3700, n_3701);
  not g7822 (n_3702, n4446);
  and g7823 (n4447, n4435, n_3702);
  not g7824 (n_3703, n4435);
  and g7825 (n4448, n_3703, n4446);
  not g7826 (n_3704, n4238);
  not g7827 (n_3705, n4448);
  and g7828 (n4449, n_3704, n_3705);
  not g7829 (n_3706, n4447);
  and g7830 (n4450, n_3706, n4449);
  not g7831 (n_3707, n4450);
  and g7832 (n4451, n_3704, n_3707);
  and g7833 (n4452, n_3706, n_3707);
  and g7834 (n4453, n_3705, n4452);
  not g7835 (n_3708, n4451);
  not g7836 (n_3709, n4453);
  and g7837 (n4454, n_3708, n_3709);
  and g7838 (n4455, \b[34] , n266);
  and g7839 (n4456, \b[32] , n284);
  and g7840 (n4457, \b[33] , n261);
  and g7846 (n4460, n_3504, n_3507);
  not g7847 (n_3714, \b[34] );
  and g7848 (n4461, n_3502, n_3714);
  and g7849 (n4462, \b[33] , \b[34] );
  not g7850 (n_3715, n4461);
  not g7851 (n_3716, n4462);
  and g7852 (n4463, n_3715, n_3716);
  not g7853 (n_3717, n4460);
  and g7854 (n4464, n_3717, n4463);
  not g7855 (n_3718, n4463);
  and g7856 (n4465, n4460, n_3718);
  not g7857 (n_3719, n4464);
  not g7858 (n_3720, n4465);
  and g7859 (n4466, n_3719, n_3720);
  and g7860 (n4467, n269, n4466);
  not g7863 (n_3722, n4468);
  and g7864 (n4469, \a[2] , n_3722);
  not g7865 (n_3723, n4469);
  and g7866 (n4470, \a[2] , n_3723);
  and g7867 (n4471, n_3722, n_3723);
  not g7868 (n_3724, n4470);
  not g7869 (n_3725, n4471);
  and g7870 (n4472, n_3724, n_3725);
  not g7871 (n_3726, n4454);
  and g7872 (n4473, n_3726, n4472);
  not g7873 (n_3727, n4472);
  and g7874 (n4474, n4454, n_3727);
  not g7875 (n_3728, n4473);
  not g7876 (n_3729, n4474);
  and g7877 (n4475, n_3728, n_3729);
  not g7878 (n_3730, n4236);
  not g7879 (n_3731, n4475);
  and g7880 (n4476, n_3730, n_3731);
  and g7881 (n4477, n4236, n4475);
  not g7882 (n_3732, n4476);
  not g7883 (n_3733, n4477);
  and g7884 (\f[34] , n_3732, n_3733);
  and g7885 (n4479, n_3726, n_3727);
  not g7886 (n_3734, n4479);
  and g7887 (n4480, n_3732, n_3734);
  and g7888 (n4481, \b[29] , n511);
  and g7889 (n4482, \b[27] , n541);
  and g7890 (n4483, \b[28] , n506);
  and g7896 (n4486, n514, n3383);
  not g7899 (n_3739, n4487);
  and g7900 (n4488, \a[8] , n_3739);
  not g7901 (n_3740, n4488);
  and g7902 (n4489, \a[8] , n_3740);
  and g7903 (n4490, n_3739, n_3740);
  not g7904 (n_3741, n4489);
  not g7905 (n_3742, n4490);
  and g7906 (n4491, n_3741, n_3742);
  and g7907 (n4492, \b[26] , n700);
  and g7908 (n4493, \b[24] , n767);
  and g7909 (n4494, \b[25] , n695);
  and g7915 (n4497, n703, n2813);
  not g7918 (n_3747, n4498);
  and g7919 (n4499, \a[11] , n_3747);
  not g7920 (n_3748, n4499);
  and g7921 (n4500, \a[11] , n_3748);
  and g7922 (n4501, n_3747, n_3748);
  not g7923 (n_3749, n4500);
  not g7924 (n_3750, n4501);
  and g7925 (n4502, n_3749, n_3750);
  and g7926 (n4503, n_3653, n_3660);
  and g7927 (n4504, n_3637, n_3643);
  and g7928 (n4505, \b[17] , n1627);
  and g7929 (n4506, \b[15] , n1763);
  and g7930 (n4507, \b[16] , n1622);
  and g7936 (n4510, n1356, n1630);
  not g7939 (n_3755, n4511);
  and g7940 (n4512, \a[20] , n_3755);
  not g7941 (n_3756, n4512);
  and g7942 (n4513, \a[20] , n_3756);
  and g7943 (n4514, n_3755, n_3756);
  not g7944 (n_3757, n4513);
  not g7945 (n_3758, n4514);
  and g7946 (n4515, n_3757, n_3758);
  and g7947 (n4516, n_3587, n_3593);
  and g7948 (n4517, \b[11] , n2539);
  and g7949 (n4518, \b[9] , n2685);
  and g7950 (n4519, \b[10] , n2534);
  and g7956 (n4522, n818, n2542);
  not g7959 (n_3763, n4523);
  and g7960 (n4524, \a[26] , n_3763);
  not g7961 (n_3764, n4524);
  and g7962 (n4525, \a[26] , n_3764);
  and g7963 (n4526, n_3763, n_3764);
  not g7964 (n_3765, n4525);
  not g7965 (n_3766, n4526);
  and g7966 (n4527, n_3765, n_3766);
  and g7967 (n4528, n_3581, n_3584);
  and g7968 (n4529, n_3573, n_3576);
  and g7969 (n4530, \b[2] , n4287);
  and g7970 (n4531, n4067, n_3560);
  and g7971 (n4532, n4281, n4531);
  and g7972 (n4533, \b[0] , n4532);
  and g7973 (n4534, \b[1] , n4282);
  and g7979 (n4537, n296, n4290);
  not g7982 (n_3771, n4538);
  and g7983 (n4539, \a[35] , n_3771);
  not g7984 (n_3772, n4539);
  and g7985 (n4540, \a[35] , n_3772);
  and g7986 (n4541, n_3771, n_3772);
  not g7987 (n_3773, n4540);
  not g7988 (n_3774, n4541);
  and g7989 (n4542, n_3773, n_3774);
  and g7990 (n4543, n_3568, n4542);
  not g7991 (n_3775, n4542);
  and g7992 (n4544, n4297, n_3775);
  not g7993 (n_3776, n4543);
  not g7994 (n_3777, n4544);
  and g7995 (n4545, n_3776, n_3777);
  and g7996 (n4546, \b[5] , n3638);
  and g7997 (n4547, \b[3] , n3843);
  and g7998 (n4548, \b[4] , n3633);
  and g8004 (n4551, n394, n3641);
  not g8007 (n_3782, n4552);
  and g8008 (n4553, \a[32] , n_3782);
  not g8009 (n_3783, n4553);
  and g8010 (n4554, \a[32] , n_3783);
  and g8011 (n4555, n_3782, n_3783);
  not g8012 (n_3784, n4554);
  not g8013 (n_3785, n4555);
  and g8014 (n4556, n_3784, n_3785);
  not g8015 (n_3786, n4556);
  and g8016 (n4557, n4545, n_3786);
  not g8017 (n_3787, n4545);
  and g8018 (n4558, n_3787, n4556);
  not g8019 (n_3788, n4529);
  not g8020 (n_3789, n4558);
  and g8021 (n4559, n_3788, n_3789);
  not g8022 (n_3790, n4557);
  and g8023 (n4560, n_3790, n4559);
  not g8024 (n_3791, n4560);
  and g8025 (n4561, n_3788, n_3791);
  and g8026 (n4562, n_3790, n_3791);
  and g8027 (n4563, n_3789, n4562);
  not g8028 (n_3792, n4561);
  not g8029 (n_3793, n4563);
  and g8030 (n4564, n_3792, n_3793);
  and g8031 (n4565, \b[8] , n3050);
  and g8032 (n4566, \b[6] , n3243);
  and g8033 (n4567, \b[7] , n3045);
  and g8039 (n4570, n585, n3053);
  not g8042 (n_3798, n4571);
  and g8043 (n4572, \a[29] , n_3798);
  not g8044 (n_3799, n4572);
  and g8045 (n4573, \a[29] , n_3799);
  and g8046 (n4574, n_3798, n_3799);
  not g8047 (n_3800, n4573);
  not g8048 (n_3801, n4574);
  and g8049 (n4575, n_3800, n_3801);
  not g8050 (n_3802, n4564);
  not g8051 (n_3803, n4575);
  and g8052 (n4576, n_3802, n_3803);
  not g8053 (n_3804, n4576);
  and g8054 (n4577, n_3802, n_3804);
  and g8055 (n4578, n_3803, n_3804);
  not g8056 (n_3805, n4577);
  not g8057 (n_3806, n4578);
  and g8058 (n4579, n_3805, n_3806);
  not g8059 (n_3807, n4528);
  not g8060 (n_3808, n4579);
  and g8061 (n4580, n_3807, n_3808);
  and g8062 (n4581, n4528, n4579);
  not g8063 (n_3809, n4580);
  not g8064 (n_3810, n4581);
  and g8065 (n4582, n_3809, n_3810);
  not g8066 (n_3811, n4527);
  and g8067 (n4583, n_3811, n4582);
  not g8068 (n_3812, n4583);
  and g8069 (n4584, n_3811, n_3812);
  and g8070 (n4585, n4582, n_3812);
  not g8071 (n_3813, n4584);
  not g8072 (n_3814, n4585);
  and g8073 (n4586, n_3813, n_3814);
  not g8074 (n_3815, n4516);
  not g8075 (n_3816, n4586);
  and g8076 (n4587, n_3815, n_3816);
  not g8077 (n_3817, n4587);
  and g8078 (n4588, n_3815, n_3817);
  and g8079 (n4589, n_3816, n_3817);
  not g8080 (n_3818, n4588);
  not g8081 (n_3819, n4589);
  and g8082 (n4590, n_3818, n_3819);
  and g8083 (n4591, \b[14] , n2048);
  and g8084 (n4592, \b[12] , n2198);
  and g8085 (n4593, \b[13] , n2043);
  and g8091 (n4596, n1034, n2051);
  not g8094 (n_3824, n4597);
  and g8095 (n4598, \a[23] , n_3824);
  not g8096 (n_3825, n4598);
  and g8097 (n4599, \a[23] , n_3825);
  and g8098 (n4600, n_3824, n_3825);
  not g8099 (n_3826, n4599);
  not g8100 (n_3827, n4600);
  and g8101 (n4601, n_3826, n_3827);
  and g8102 (n4602, n4590, n4601);
  not g8103 (n_3828, n4590);
  not g8104 (n_3829, n4601);
  and g8105 (n4603, n_3828, n_3829);
  not g8106 (n_3830, n4602);
  not g8107 (n_3831, n4603);
  and g8108 (n4604, n_3830, n_3831);
  not g8109 (n_3832, n4336);
  and g8110 (n4605, n_3832, n4604);
  not g8111 (n_3833, n4604);
  and g8112 (n4606, n4336, n_3833);
  not g8113 (n_3834, n4605);
  not g8114 (n_3835, n4606);
  and g8115 (n4607, n_3834, n_3835);
  not g8116 (n_3836, n4515);
  and g8117 (n4608, n_3836, n4607);
  not g8118 (n_3837, n4608);
  and g8119 (n4609, n4607, n_3837);
  and g8120 (n4610, n_3836, n_3837);
  not g8121 (n_3838, n4609);
  not g8122 (n_3839, n4610);
  and g8123 (n4611, n_3838, n_3839);
  and g8124 (n4612, n_3620, n_3627);
  and g8125 (n4613, n4611, n4612);
  not g8126 (n_3840, n4611);
  not g8127 (n_3841, n4612);
  and g8128 (n4614, n_3840, n_3841);
  not g8129 (n_3842, n4613);
  not g8130 (n_3843, n4614);
  and g8131 (n4615, n_3842, n_3843);
  and g8132 (n4616, \b[20] , n1302);
  and g8133 (n4617, \b[18] , n1391);
  and g8134 (n4618, \b[19] , n1297);
  and g8140 (n4621, n1305, n1846);
  not g8143 (n_3848, n4622);
  and g8144 (n4623, \a[17] , n_3848);
  not g8145 (n_3849, n4623);
  and g8146 (n4624, \a[17] , n_3849);
  and g8147 (n4625, n_3848, n_3849);
  not g8148 (n_3850, n4624);
  not g8149 (n_3851, n4625);
  and g8150 (n4626, n_3850, n_3851);
  not g8151 (n_3852, n4626);
  and g8152 (n4627, n4615, n_3852);
  not g8153 (n_3853, n4615);
  and g8154 (n4628, n_3853, n4626);
  not g8155 (n_3854, n4504);
  not g8156 (n_3855, n4628);
  and g8157 (n4629, n_3854, n_3855);
  not g8158 (n_3856, n4627);
  and g8159 (n4630, n_3856, n4629);
  not g8160 (n_3857, n4630);
  and g8161 (n4631, n_3854, n_3857);
  and g8162 (n4632, n_3856, n_3857);
  and g8163 (n4633, n_3855, n4632);
  not g8164 (n_3858, n4631);
  not g8165 (n_3859, n4633);
  and g8166 (n4634, n_3858, n_3859);
  and g8167 (n4635, \b[23] , n951);
  and g8168 (n4636, \b[21] , n1056);
  and g8169 (n4637, \b[22] , n946);
  and g8175 (n4640, n954, n2300);
  not g8178 (n_3864, n4641);
  and g8179 (n4642, \a[14] , n_3864);
  not g8180 (n_3865, n4642);
  and g8181 (n4643, \a[14] , n_3865);
  and g8182 (n4644, n_3864, n_3865);
  not g8183 (n_3866, n4643);
  not g8184 (n_3867, n4644);
  and g8185 (n4645, n_3866, n_3867);
  and g8186 (n4646, n4634, n4645);
  not g8187 (n_3868, n4634);
  not g8188 (n_3869, n4645);
  and g8189 (n4647, n_3868, n_3869);
  not g8190 (n_3870, n4646);
  not g8191 (n_3871, n4647);
  and g8192 (n4648, n_3870, n_3871);
  not g8193 (n_3872, n4503);
  and g8194 (n4649, n_3872, n4648);
  not g8195 (n_3873, n4648);
  and g8196 (n4650, n4503, n_3873);
  not g8197 (n_3874, n4649);
  not g8198 (n_3875, n4650);
  and g8199 (n4651, n_3874, n_3875);
  not g8200 (n_3876, n4651);
  and g8201 (n4652, n4502, n_3876);
  not g8202 (n_3877, n4502);
  and g8203 (n4653, n_3877, n4651);
  not g8204 (n_3878, n4652);
  not g8205 (n_3879, n4653);
  and g8206 (n4654, n_3878, n_3879);
  not g8207 (n_3880, n4414);
  and g8208 (n4655, n_3880, n4654);
  not g8209 (n_3881, n4654);
  and g8210 (n4656, n4414, n_3881);
  not g8211 (n_3882, n4655);
  not g8212 (n_3883, n4656);
  and g8213 (n4657, n_3882, n_3883);
  not g8214 (n_3884, n4491);
  and g8215 (n4658, n_3884, n4657);
  not g8216 (n_3885, n4658);
  and g8217 (n4659, n4657, n_3885);
  and g8218 (n4660, n_3884, n_3885);
  not g8219 (n_3886, n4659);
  not g8220 (n_3887, n4660);
  and g8221 (n4661, n_3886, n_3887);
  and g8222 (n4662, n_3687, n_3693);
  and g8223 (n4663, n4661, n4662);
  not g8224 (n_3888, n4661);
  not g8225 (n_3889, n4662);
  and g8226 (n4664, n_3888, n_3889);
  not g8227 (n_3890, n4663);
  not g8228 (n_3891, n4664);
  and g8229 (n4665, n_3890, n_3891);
  and g8230 (n4666, \b[32] , n362);
  and g8231 (n4667, \b[30] , n403);
  and g8232 (n4668, \b[31] , n357);
  and g8238 (n4671, n365, n4013);
  not g8241 (n_3896, n4672);
  and g8242 (n4673, \a[5] , n_3896);
  not g8243 (n_3897, n4673);
  and g8244 (n4674, \a[5] , n_3897);
  and g8245 (n4675, n_3896, n_3897);
  not g8246 (n_3898, n4674);
  not g8247 (n_3899, n4675);
  and g8248 (n4676, n_3898, n_3899);
  not g8249 (n_3900, n4676);
  and g8250 (n4677, n4665, n_3900);
  not g8251 (n_3901, n4665);
  and g8252 (n4678, n_3901, n4676);
  not g8253 (n_3902, n4452);
  not g8254 (n_3903, n4678);
  and g8255 (n4679, n_3902, n_3903);
  not g8256 (n_3904, n4677);
  and g8257 (n4680, n_3904, n4679);
  not g8258 (n_3905, n4680);
  and g8259 (n4681, n_3902, n_3905);
  and g8260 (n4682, n_3904, n_3905);
  and g8261 (n4683, n_3903, n4682);
  not g8262 (n_3906, n4681);
  not g8263 (n_3907, n4683);
  and g8264 (n4684, n_3906, n_3907);
  and g8265 (n4685, \b[35] , n266);
  and g8266 (n4686, \b[33] , n284);
  and g8267 (n4687, \b[34] , n261);
  and g8273 (n4690, n_3716, n_3719);
  not g8274 (n_3912, \b[35] );
  and g8275 (n4691, n_3714, n_3912);
  and g8276 (n4692, \b[34] , \b[35] );
  not g8277 (n_3913, n4691);
  not g8278 (n_3914, n4692);
  and g8279 (n4693, n_3913, n_3914);
  not g8280 (n_3915, n4690);
  and g8281 (n4694, n_3915, n4693);
  not g8282 (n_3916, n4693);
  and g8283 (n4695, n4690, n_3916);
  not g8284 (n_3917, n4694);
  not g8285 (n_3918, n4695);
  and g8286 (n4696, n_3917, n_3918);
  and g8287 (n4697, n269, n4696);
  not g8290 (n_3920, n4698);
  and g8291 (n4699, \a[2] , n_3920);
  not g8292 (n_3921, n4699);
  and g8293 (n4700, \a[2] , n_3921);
  and g8294 (n4701, n_3920, n_3921);
  not g8295 (n_3922, n4700);
  not g8296 (n_3923, n4701);
  and g8297 (n4702, n_3922, n_3923);
  not g8298 (n_3924, n4684);
  and g8299 (n4703, n_3924, n4702);
  not g8300 (n_3925, n4702);
  and g8301 (n4704, n4684, n_3925);
  not g8302 (n_3926, n4703);
  not g8303 (n_3927, n4704);
  and g8304 (n4705, n_3926, n_3927);
  not g8305 (n_3928, n4480);
  not g8306 (n_3929, n4705);
  and g8307 (n4706, n_3928, n_3929);
  and g8308 (n4707, n4480, n4705);
  not g8309 (n_3930, n4706);
  not g8310 (n_3931, n4707);
  and g8311 (\f[35] , n_3930, n_3931);
  and g8312 (n4709, \b[33] , n362);
  and g8313 (n4710, \b[31] , n403);
  and g8314 (n4711, \b[32] , n357);
  and g8320 (n4714, n365, n4223);
  not g8323 (n_3936, n4715);
  and g8324 (n4716, \a[5] , n_3936);
  not g8325 (n_3937, n4716);
  and g8326 (n4717, \a[5] , n_3937);
  and g8327 (n4718, n_3936, n_3937);
  not g8328 (n_3938, n4717);
  not g8329 (n_3939, n4718);
  and g8330 (n4719, n_3938, n_3939);
  and g8331 (n4720, n_3885, n_3891);
  and g8332 (n4721, n_3879, n_3882);
  and g8333 (n4722, \b[27] , n700);
  and g8334 (n4723, \b[25] , n767);
  and g8335 (n4724, \b[26] , n695);
  and g8341 (n4727, n703, n2990);
  not g8344 (n_3944, n4728);
  and g8345 (n4729, \a[11] , n_3944);
  not g8346 (n_3945, n4729);
  and g8347 (n4730, \a[11] , n_3945);
  and g8348 (n4731, n_3944, n_3945);
  not g8349 (n_3946, n4730);
  not g8350 (n_3947, n4731);
  and g8351 (n4732, n_3946, n_3947);
  and g8352 (n4733, n_3871, n_3874);
  and g8353 (n4734, n_3837, n_3843);
  and g8354 (n4735, n_3831, n_3834);
  and g8355 (n4736, \b[15] , n2048);
  and g8356 (n4737, \b[13] , n2198);
  and g8357 (n4738, \b[14] , n2043);
  and g8363 (n4741, n1131, n2051);
  not g8366 (n_3952, n4742);
  and g8367 (n4743, \a[23] , n_3952);
  not g8368 (n_3953, n4743);
  and g8369 (n4744, \a[23] , n_3953);
  and g8370 (n4745, n_3952, n_3953);
  not g8371 (n_3954, n4744);
  not g8372 (n_3955, n4745);
  and g8373 (n4746, n_3954, n_3955);
  and g8374 (n4747, n_3804, n_3809);
  and g8375 (n4748, \b[6] , n3638);
  and g8376 (n4749, \b[4] , n3843);
  and g8377 (n4750, \b[5] , n3633);
  and g8383 (n4753, n459, n3641);
  not g8386 (n_3960, n4754);
  and g8387 (n4755, \a[32] , n_3960);
  not g8388 (n_3961, n4755);
  and g8389 (n4756, \a[32] , n_3961);
  and g8390 (n4757, n_3960, n_3961);
  not g8391 (n_3962, n4756);
  not g8392 (n_3963, n4757);
  and g8393 (n4758, n_3962, n_3963);
  not g8394 (n_3965, \a[36] );
  and g8395 (n4759, \a[35] , n_3965);
  and g8396 (n4760, n_3555, \a[36] );
  not g8397 (n_3966, n4759);
  not g8398 (n_3967, n4760);
  and g8399 (n4761, n_3966, n_3967);
  not g8400 (n_3968, n4761);
  and g8401 (n4762, \b[0] , n_3968);
  and g8402 (n4763, n_3777, n4762);
  not g8403 (n_3969, n4762);
  and g8404 (n4764, n4544, n_3969);
  not g8405 (n_3970, n4763);
  not g8406 (n_3971, n4764);
  and g8407 (n4765, n_3970, n_3971);
  and g8408 (n4766, \b[3] , n4287);
  and g8409 (n4767, \b[1] , n4532);
  and g8410 (n4768, \b[2] , n4282);
  and g8416 (n4771, n318, n4290);
  not g8419 (n_3976, n4772);
  and g8420 (n4773, \a[35] , n_3976);
  not g8421 (n_3977, n4773);
  and g8422 (n4774, \a[35] , n_3977);
  and g8423 (n4775, n_3976, n_3977);
  not g8424 (n_3978, n4774);
  not g8425 (n_3979, n4775);
  and g8426 (n4776, n_3978, n_3979);
  not g8427 (n_3980, n4765);
  not g8428 (n_3981, n4776);
  and g8429 (n4777, n_3980, n_3981);
  and g8430 (n4778, n4765, n4776);
  not g8431 (n_3982, n4777);
  not g8432 (n_3983, n4778);
  and g8433 (n4779, n_3982, n_3983);
  not g8434 (n_3984, n4758);
  and g8435 (n4780, n_3984, n4779);
  not g8436 (n_3985, n4780);
  and g8437 (n4781, n4779, n_3985);
  and g8438 (n4782, n_3984, n_3985);
  not g8439 (n_3986, n4781);
  not g8440 (n_3987, n4782);
  and g8441 (n4783, n_3986, n_3987);
  not g8442 (n_3988, n4562);
  and g8443 (n4784, n_3988, n4783);
  not g8444 (n_3989, n4783);
  and g8445 (n4785, n4562, n_3989);
  not g8446 (n_3990, n4784);
  not g8447 (n_3991, n4785);
  and g8448 (n4786, n_3990, n_3991);
  and g8449 (n4787, \b[9] , n3050);
  and g8450 (n4788, \b[7] , n3243);
  and g8451 (n4789, \b[8] , n3045);
  and g8457 (n4792, n651, n3053);
  not g8460 (n_3996, n4793);
  and g8461 (n4794, \a[29] , n_3996);
  not g8462 (n_3997, n4794);
  and g8463 (n4795, \a[29] , n_3997);
  and g8464 (n4796, n_3996, n_3997);
  not g8465 (n_3998, n4795);
  not g8466 (n_3999, n4796);
  and g8467 (n4797, n_3998, n_3999);
  not g8468 (n_4000, n4786);
  not g8469 (n_4001, n4797);
  and g8470 (n4798, n_4000, n_4001);
  and g8471 (n4799, n4786, n4797);
  not g8472 (n_4002, n4798);
  not g8473 (n_4003, n4799);
  and g8474 (n4800, n_4002, n_4003);
  not g8475 (n_4004, n4800);
  and g8476 (n4801, n4747, n_4004);
  not g8477 (n_4005, n4747);
  and g8478 (n4802, n_4005, n4800);
  not g8479 (n_4006, n4801);
  not g8480 (n_4007, n4802);
  and g8481 (n4803, n_4006, n_4007);
  and g8482 (n4804, \b[12] , n2539);
  and g8483 (n4805, \b[10] , n2685);
  and g8484 (n4806, \b[11] , n2534);
  and g8490 (n4809, n842, n2542);
  not g8493 (n_4012, n4810);
  and g8494 (n4811, \a[26] , n_4012);
  not g8495 (n_4013, n4811);
  and g8496 (n4812, \a[26] , n_4013);
  and g8497 (n4813, n_4012, n_4013);
  not g8498 (n_4014, n4812);
  not g8499 (n_4015, n4813);
  and g8500 (n4814, n_4014, n_4015);
  not g8501 (n_4016, n4803);
  and g8502 (n4815, n_4016, n4814);
  not g8503 (n_4017, n4814);
  and g8504 (n4816, n4803, n_4017);
  not g8505 (n_4018, n4815);
  not g8506 (n_4019, n4816);
  and g8507 (n4817, n_4018, n_4019);
  and g8508 (n4818, n_3812, n_3817);
  not g8509 (n_4020, n4818);
  and g8510 (n4819, n4817, n_4020);
  not g8511 (n_4021, n4817);
  and g8512 (n4820, n_4021, n4818);
  not g8513 (n_4022, n4819);
  not g8514 (n_4023, n4820);
  and g8515 (n4821, n_4022, n_4023);
  not g8516 (n_4024, n4746);
  and g8517 (n4822, n_4024, n4821);
  not g8518 (n_4025, n4822);
  and g8519 (n4823, n4821, n_4025);
  and g8520 (n4824, n_4024, n_4025);
  not g8521 (n_4026, n4823);
  not g8522 (n_4027, n4824);
  and g8523 (n4825, n_4026, n_4027);
  not g8524 (n_4028, n4735);
  and g8525 (n4826, n_4028, n4825);
  not g8526 (n_4029, n4825);
  and g8527 (n4827, n4735, n_4029);
  not g8528 (n_4030, n4826);
  not g8529 (n_4031, n4827);
  and g8530 (n4828, n_4030, n_4031);
  and g8531 (n4829, \b[18] , n1627);
  and g8532 (n4830, \b[16] , n1763);
  and g8533 (n4831, \b[17] , n1622);
  and g8539 (n4834, n1566, n1630);
  not g8542 (n_4036, n4835);
  and g8543 (n4836, \a[20] , n_4036);
  not g8544 (n_4037, n4836);
  and g8545 (n4837, \a[20] , n_4037);
  and g8546 (n4838, n_4036, n_4037);
  not g8547 (n_4038, n4837);
  not g8548 (n_4039, n4838);
  and g8549 (n4839, n_4038, n_4039);
  not g8550 (n_4040, n4828);
  not g8551 (n_4041, n4839);
  and g8552 (n4840, n_4040, n_4041);
  and g8553 (n4841, n4828, n4839);
  not g8554 (n_4042, n4840);
  not g8555 (n_4043, n4841);
  and g8556 (n4842, n_4042, n_4043);
  not g8557 (n_4044, n4842);
  and g8558 (n4843, n4734, n_4044);
  not g8559 (n_4045, n4734);
  and g8560 (n4844, n_4045, n4842);
  not g8561 (n_4046, n4843);
  not g8562 (n_4047, n4844);
  and g8563 (n4845, n_4046, n_4047);
  and g8564 (n4846, \b[21] , n1302);
  and g8565 (n4847, \b[19] , n1391);
  and g8566 (n4848, \b[20] , n1297);
  and g8572 (n4851, n1305, n1984);
  not g8575 (n_4052, n4852);
  and g8576 (n4853, \a[17] , n_4052);
  not g8577 (n_4053, n4853);
  and g8578 (n4854, \a[17] , n_4053);
  and g8579 (n4855, n_4052, n_4053);
  not g8580 (n_4054, n4854);
  not g8581 (n_4055, n4855);
  and g8582 (n4856, n_4054, n_4055);
  not g8583 (n_4056, n4856);
  and g8584 (n4857, n4845, n_4056);
  not g8585 (n_4057, n4857);
  and g8586 (n4858, n4845, n_4057);
  and g8587 (n4859, n_4056, n_4057);
  not g8588 (n_4058, n4858);
  not g8589 (n_4059, n4859);
  and g8590 (n4860, n_4058, n_4059);
  not g8591 (n_4060, n4632);
  and g8592 (n4861, n_4060, n4860);
  not g8593 (n_4061, n4860);
  and g8594 (n4862, n4632, n_4061);
  not g8595 (n_4062, n4861);
  not g8596 (n_4063, n4862);
  and g8597 (n4863, n_4062, n_4063);
  and g8598 (n4864, \b[24] , n951);
  and g8599 (n4865, \b[22] , n1056);
  and g8600 (n4866, \b[23] , n946);
  and g8606 (n4869, n954, n2458);
  not g8609 (n_4068, n4870);
  and g8610 (n4871, \a[14] , n_4068);
  not g8611 (n_4069, n4871);
  and g8612 (n4872, \a[14] , n_4069);
  and g8613 (n4873, n_4068, n_4069);
  not g8614 (n_4070, n4872);
  not g8615 (n_4071, n4873);
  and g8616 (n4874, n_4070, n_4071);
  and g8617 (n4875, n4863, n4874);
  not g8618 (n_4072, n4863);
  not g8619 (n_4073, n4874);
  and g8620 (n4876, n_4072, n_4073);
  not g8621 (n_4074, n4875);
  not g8622 (n_4075, n4876);
  and g8623 (n4877, n_4074, n_4075);
  not g8624 (n_4076, n4733);
  and g8625 (n4878, n_4076, n4877);
  not g8626 (n_4077, n4877);
  and g8627 (n4879, n4733, n_4077);
  not g8628 (n_4078, n4878);
  not g8629 (n_4079, n4879);
  and g8630 (n4880, n_4078, n_4079);
  not g8631 (n_4080, n4732);
  and g8632 (n4881, n_4080, n4880);
  not g8633 (n_4081, n4881);
  and g8634 (n4882, n4880, n_4081);
  and g8635 (n4883, n_4080, n_4081);
  not g8636 (n_4082, n4882);
  not g8637 (n_4083, n4883);
  and g8638 (n4884, n_4082, n_4083);
  not g8639 (n_4084, n4721);
  and g8640 (n4885, n_4084, n4884);
  not g8641 (n_4085, n4884);
  and g8642 (n4886, n4721, n_4085);
  not g8643 (n_4086, n4885);
  not g8644 (n_4087, n4886);
  and g8645 (n4887, n_4086, n_4087);
  and g8646 (n4888, \b[30] , n511);
  and g8647 (n4889, \b[28] , n541);
  and g8648 (n4890, \b[29] , n506);
  and g8654 (n4893, n514, n3577);
  not g8657 (n_4092, n4894);
  and g8658 (n4895, \a[8] , n_4092);
  not g8659 (n_4093, n4895);
  and g8660 (n4896, \a[8] , n_4093);
  and g8661 (n4897, n_4092, n_4093);
  not g8662 (n_4094, n4896);
  not g8663 (n_4095, n4897);
  and g8664 (n4898, n_4094, n_4095);
  and g8665 (n4899, n4887, n4898);
  not g8666 (n_4096, n4887);
  not g8667 (n_4097, n4898);
  and g8668 (n4900, n_4096, n_4097);
  not g8669 (n_4098, n4899);
  not g8670 (n_4099, n4900);
  and g8671 (n4901, n_4098, n_4099);
  not g8672 (n_4100, n4720);
  and g8673 (n4902, n_4100, n4901);
  not g8674 (n_4101, n4901);
  and g8675 (n4903, n4720, n_4101);
  not g8676 (n_4102, n4902);
  not g8677 (n_4103, n4903);
  and g8678 (n4904, n_4102, n_4103);
  not g8679 (n_4104, n4719);
  and g8680 (n4905, n_4104, n4904);
  not g8681 (n_4105, n4904);
  and g8682 (n4906, n4719, n_4105);
  not g8683 (n_4106, n4905);
  not g8684 (n_4107, n4906);
  and g8685 (n4907, n_4106, n_4107);
  not g8686 (n_4108, n4682);
  and g8687 (n4908, n_4108, n4907);
  not g8688 (n_4109, n4907);
  and g8689 (n4909, n4682, n_4109);
  not g8690 (n_4110, n4908);
  not g8691 (n_4111, n4909);
  and g8692 (n4910, n_4110, n_4111);
  and g8693 (n4911, \b[36] , n266);
  and g8694 (n4912, \b[34] , n284);
  and g8695 (n4913, \b[35] , n261);
  and g8701 (n4916, n_3914, n_3917);
  not g8702 (n_4116, \b[36] );
  and g8703 (n4917, n_3912, n_4116);
  and g8704 (n4918, \b[35] , \b[36] );
  not g8705 (n_4117, n4917);
  not g8706 (n_4118, n4918);
  and g8707 (n4919, n_4117, n_4118);
  not g8708 (n_4119, n4916);
  and g8709 (n4920, n_4119, n4919);
  not g8710 (n_4120, n4919);
  and g8711 (n4921, n4916, n_4120);
  not g8712 (n_4121, n4920);
  not g8713 (n_4122, n4921);
  and g8714 (n4922, n_4121, n_4122);
  and g8715 (n4923, n269, n4922);
  not g8718 (n_4124, n4924);
  and g8719 (n4925, \a[2] , n_4124);
  not g8720 (n_4125, n4925);
  and g8721 (n4926, \a[2] , n_4125);
  and g8722 (n4927, n_4124, n_4125);
  not g8723 (n_4126, n4926);
  not g8724 (n_4127, n4927);
  and g8725 (n4928, n_4126, n_4127);
  not g8726 (n_4128, n4928);
  and g8727 (n4929, n4910, n_4128);
  not g8728 (n_4129, n4929);
  and g8729 (n4930, n4910, n_4129);
  and g8730 (n4931, n_4128, n_4129);
  not g8731 (n_4130, n4930);
  not g8732 (n_4131, n4931);
  and g8733 (n4932, n_4130, n_4131);
  and g8734 (n4933, n_3924, n_3925);
  not g8735 (n_4132, n4933);
  and g8736 (n4934, n_3930, n_4132);
  not g8737 (n_4133, n4932);
  not g8738 (n_4134, n4934);
  and g8739 (n4935, n_4133, n_4134);
  and g8740 (n4936, n4932, n4934);
  not g8741 (n_4135, n4935);
  not g8742 (n_4136, n4936);
  and g8743 (\f[36] , n_4135, n_4136);
  and g8744 (n4938, n_4129, n_4135);
  and g8745 (n4939, \b[34] , n362);
  and g8746 (n4940, \b[32] , n403);
  and g8747 (n4941, \b[33] , n357);
  and g8753 (n4944, n365, n4466);
  not g8756 (n_4141, n4945);
  and g8757 (n4946, \a[5] , n_4141);
  not g8758 (n_4142, n4946);
  and g8759 (n4947, \a[5] , n_4142);
  and g8760 (n4948, n_4141, n_4142);
  not g8761 (n_4143, n4947);
  not g8762 (n_4144, n4948);
  and g8763 (n4949, n_4143, n_4144);
  and g8764 (n4950, n_4099, n_4102);
  and g8765 (n4951, \b[31] , n511);
  and g8766 (n4952, \b[29] , n541);
  and g8767 (n4953, \b[30] , n506);
  and g8773 (n4956, n514, n3796);
  not g8776 (n_4149, n4957);
  and g8777 (n4958, \a[8] , n_4149);
  not g8778 (n_4150, n4958);
  and g8779 (n4959, \a[8] , n_4150);
  and g8780 (n4960, n_4149, n_4150);
  not g8781 (n_4151, n4959);
  not g8782 (n_4152, n4960);
  and g8783 (n4961, n_4151, n_4152);
  and g8784 (n4962, n_4084, n_4085);
  not g8785 (n_4153, n4962);
  and g8786 (n4963, n_4081, n_4153);
  and g8787 (n4964, n_4075, n_4078);
  and g8788 (n4965, \b[16] , n2048);
  and g8789 (n4966, \b[14] , n2198);
  and g8790 (n4967, \b[15] , n2043);
  and g8796 (n4970, n1237, n2051);
  not g8799 (n_4158, n4971);
  and g8800 (n4972, \a[23] , n_4158);
  not g8801 (n_4159, n4972);
  and g8802 (n4973, \a[23] , n_4159);
  and g8803 (n4974, n_4158, n_4159);
  not g8804 (n_4160, n4973);
  not g8805 (n_4161, n4974);
  and g8806 (n4975, n_4160, n_4161);
  and g8807 (n4976, n_4019, n_4022);
  and g8808 (n4977, \b[13] , n2539);
  and g8809 (n4978, \b[11] , n2685);
  and g8810 (n4979, \b[12] , n2534);
  and g8816 (n4982, n1008, n2542);
  not g8819 (n_4166, n4983);
  and g8820 (n4984, \a[26] , n_4166);
  not g8821 (n_4167, n4984);
  and g8822 (n4985, \a[26] , n_4167);
  and g8823 (n4986, n_4166, n_4167);
  not g8824 (n_4168, n4985);
  not g8825 (n_4169, n4986);
  and g8826 (n4987, n_4168, n_4169);
  and g8827 (n4988, n_4002, n_4007);
  and g8828 (n4989, \b[10] , n3050);
  and g8829 (n4990, \b[8] , n3243);
  and g8830 (n4991, \b[9] , n3045);
  and g8836 (n4994, n738, n3053);
  not g8839 (n_4174, n4995);
  and g8840 (n4996, \a[29] , n_4174);
  not g8841 (n_4175, n4996);
  and g8842 (n4997, \a[29] , n_4175);
  and g8843 (n4998, n_4174, n_4175);
  not g8844 (n_4176, n4997);
  not g8845 (n_4177, n4998);
  and g8846 (n4999, n_4176, n_4177);
  and g8847 (n5000, n_3988, n_3989);
  not g8848 (n_4178, n5000);
  and g8849 (n5001, n_3985, n_4178);
  and g8850 (n5002, \b[7] , n3638);
  and g8851 (n5003, \b[5] , n3843);
  and g8852 (n5004, \b[6] , n3633);
  and g8858 (n5007, n484, n3641);
  not g8861 (n_4183, n5008);
  and g8862 (n5009, \a[32] , n_4183);
  not g8863 (n_4184, n5009);
  and g8864 (n5010, \a[32] , n_4184);
  and g8865 (n5011, n_4183, n_4184);
  not g8866 (n_4185, n5010);
  not g8867 (n_4186, n5011);
  and g8868 (n5012, n_4185, n_4186);
  and g8869 (n5013, n4544, n4762);
  not g8870 (n_4187, n5013);
  and g8871 (n5014, n_3982, n_4187);
  and g8872 (n5015, \b[4] , n4287);
  and g8873 (n5016, \b[2] , n4532);
  and g8874 (n5017, \b[3] , n4282);
  and g8880 (n5020, n346, n4290);
  not g8883 (n_4192, n5021);
  and g8884 (n5022, \a[35] , n_4192);
  not g8885 (n_4193, n5022);
  and g8886 (n5023, \a[35] , n_4193);
  and g8887 (n5024, n_4192, n_4193);
  not g8888 (n_4194, n5023);
  not g8889 (n_4195, n5024);
  and g8890 (n5025, n_4194, n_4195);
  and g8891 (n5026, \a[38] , n_3969);
  and g8892 (n5027, n_3965, \a[37] );
  not g8893 (n_4198, \a[37] );
  and g8894 (n5028, \a[36] , n_4198);
  not g8895 (n_4199, n5027);
  not g8896 (n_4200, n5028);
  and g8897 (n5029, n_4199, n_4200);
  not g8898 (n_4201, n5029);
  and g8899 (n5030, n4761, n_4201);
  and g8900 (n5031, \b[0] , n5030);
  and g8901 (n5032, n_4198, \a[38] );
  not g8902 (n_4202, \a[38] );
  and g8903 (n5033, \a[37] , n_4202);
  not g8904 (n_4203, n5032);
  not g8905 (n_4204, n5033);
  and g8906 (n5034, n_4203, n_4204);
  and g8907 (n5035, n_3968, n5034);
  and g8908 (n5036, \b[1] , n5035);
  not g8909 (n_4205, n5031);
  not g8910 (n_4206, n5036);
  and g8911 (n5037, n_4205, n_4206);
  not g8912 (n_4207, n5034);
  and g8913 (n5038, n_3968, n_4207);
  and g8914 (n5039, n_21, n5038);
  not g8915 (n_4208, n5039);
  and g8916 (n5040, n5037, n_4208);
  not g8917 (n_4209, n5040);
  and g8918 (n5041, \a[38] , n_4209);
  not g8919 (n_4210, n5041);
  and g8920 (n5042, \a[38] , n_4210);
  and g8921 (n5043, n_4209, n_4210);
  not g8922 (n_4211, n5042);
  not g8923 (n_4212, n5043);
  and g8924 (n5044, n_4211, n_4212);
  not g8925 (n_4213, n5044);
  and g8926 (n5045, n5026, n_4213);
  not g8927 (n_4214, n5026);
  and g8928 (n5046, n_4214, n5044);
  not g8929 (n_4215, n5045);
  not g8930 (n_4216, n5046);
  and g8931 (n5047, n_4215, n_4216);
  not g8932 (n_4217, n5047);
  and g8933 (n5048, n5025, n_4217);
  not g8934 (n_4218, n5025);
  and g8935 (n5049, n_4218, n5047);
  not g8936 (n_4219, n5048);
  not g8937 (n_4220, n5049);
  and g8938 (n5050, n_4219, n_4220);
  not g8939 (n_4221, n5014);
  and g8940 (n5051, n_4221, n5050);
  not g8941 (n_4222, n5050);
  and g8942 (n5052, n5014, n_4222);
  not g8943 (n_4223, n5051);
  not g8944 (n_4224, n5052);
  and g8945 (n5053, n_4223, n_4224);
  not g8946 (n_4225, n5053);
  and g8947 (n5054, n5012, n_4225);
  not g8948 (n_4226, n5012);
  and g8949 (n5055, n_4226, n5053);
  not g8950 (n_4227, n5054);
  not g8951 (n_4228, n5055);
  and g8952 (n5056, n_4227, n_4228);
  not g8953 (n_4229, n5001);
  and g8954 (n5057, n_4229, n5056);
  not g8955 (n_4230, n5056);
  and g8956 (n5058, n5001, n_4230);
  not g8957 (n_4231, n5057);
  not g8958 (n_4232, n5058);
  and g8959 (n5059, n_4231, n_4232);
  not g8960 (n_4233, n5059);
  and g8961 (n5060, n4999, n_4233);
  not g8962 (n_4234, n4999);
  and g8963 (n5061, n_4234, n5059);
  not g8964 (n_4235, n5060);
  not g8965 (n_4236, n5061);
  and g8966 (n5062, n_4235, n_4236);
  not g8967 (n_4237, n4988);
  and g8968 (n5063, n_4237, n5062);
  not g8969 (n_4238, n5062);
  and g8970 (n5064, n4988, n_4238);
  not g8971 (n_4239, n5063);
  not g8972 (n_4240, n5064);
  and g8973 (n5065, n_4239, n_4240);
  not g8974 (n_4241, n5065);
  and g8975 (n5066, n4987, n_4241);
  not g8976 (n_4242, n4987);
  and g8977 (n5067, n_4242, n5065);
  not g8978 (n_4243, n5066);
  not g8979 (n_4244, n5067);
  and g8980 (n5068, n_4243, n_4244);
  not g8981 (n_4245, n4976);
  and g8982 (n5069, n_4245, n5068);
  not g8983 (n_4246, n5068);
  and g8984 (n5070, n4976, n_4246);
  not g8985 (n_4247, n5069);
  not g8986 (n_4248, n5070);
  and g8987 (n5071, n_4247, n_4248);
  not g8988 (n_4249, n4975);
  and g8989 (n5072, n_4249, n5071);
  not g8990 (n_4250, n5072);
  and g8991 (n5073, n5071, n_4250);
  and g8992 (n5074, n_4249, n_4250);
  not g8993 (n_4251, n5073);
  not g8994 (n_4252, n5074);
  and g8995 (n5075, n_4251, n_4252);
  and g8996 (n5076, n_4028, n_4029);
  not g8997 (n_4253, n5076);
  and g8998 (n5077, n_4025, n_4253);
  and g8999 (n5078, n5075, n5077);
  not g9000 (n_4254, n5075);
  not g9001 (n_4255, n5077);
  and g9002 (n5079, n_4254, n_4255);
  not g9003 (n_4256, n5078);
  not g9004 (n_4257, n5079);
  and g9005 (n5080, n_4256, n_4257);
  and g9006 (n5081, \b[19] , n1627);
  and g9007 (n5082, \b[17] , n1763);
  and g9008 (n5083, \b[18] , n1622);
  and g9014 (n5086, n1630, n1708);
  not g9017 (n_4262, n5087);
  and g9018 (n5088, \a[20] , n_4262);
  not g9019 (n_4263, n5088);
  and g9020 (n5089, \a[20] , n_4263);
  and g9021 (n5090, n_4262, n_4263);
  not g9022 (n_4264, n5089);
  not g9023 (n_4265, n5090);
  and g9024 (n5091, n_4264, n_4265);
  not g9025 (n_4266, n5091);
  and g9026 (n5092, n5080, n_4266);
  not g9027 (n_4267, n5092);
  and g9028 (n5093, n5080, n_4267);
  and g9029 (n5094, n_4266, n_4267);
  not g9030 (n_4268, n5093);
  not g9031 (n_4269, n5094);
  and g9032 (n5095, n_4268, n_4269);
  and g9033 (n5096, n_4042, n_4047);
  and g9034 (n5097, n5095, n5096);
  not g9035 (n_4270, n5095);
  not g9036 (n_4271, n5096);
  and g9037 (n5098, n_4270, n_4271);
  not g9038 (n_4272, n5097);
  not g9039 (n_4273, n5098);
  and g9040 (n5099, n_4272, n_4273);
  and g9041 (n5100, \b[22] , n1302);
  and g9042 (n5101, \b[20] , n1391);
  and g9043 (n5102, \b[21] , n1297);
  and g9049 (n5105, n1305, n2145);
  not g9052 (n_4278, n5106);
  and g9053 (n5107, \a[17] , n_4278);
  not g9054 (n_4279, n5107);
  and g9055 (n5108, \a[17] , n_4279);
  and g9056 (n5109, n_4278, n_4279);
  not g9057 (n_4280, n5108);
  not g9058 (n_4281, n5109);
  and g9059 (n5110, n_4280, n_4281);
  not g9060 (n_4282, n5110);
  and g9061 (n5111, n5099, n_4282);
  not g9062 (n_4283, n5111);
  and g9063 (n5112, n5099, n_4283);
  and g9064 (n5113, n_4282, n_4283);
  not g9065 (n_4284, n5112);
  not g9066 (n_4285, n5113);
  and g9067 (n5114, n_4284, n_4285);
  and g9068 (n5115, n_4060, n_4061);
  not g9069 (n_4286, n5115);
  and g9070 (n5116, n_4057, n_4286);
  and g9071 (n5117, n5114, n5116);
  not g9072 (n_4287, n5114);
  not g9073 (n_4288, n5116);
  and g9074 (n5118, n_4287, n_4288);
  not g9075 (n_4289, n5117);
  not g9076 (n_4290, n5118);
  and g9077 (n5119, n_4289, n_4290);
  and g9078 (n5120, \b[25] , n951);
  and g9079 (n5121, \b[23] , n1056);
  and g9080 (n5122, \b[24] , n946);
  and g9086 (n5125, n954, n2485);
  not g9089 (n_4295, n5126);
  and g9090 (n5127, \a[14] , n_4295);
  not g9091 (n_4296, n5127);
  and g9092 (n5128, \a[14] , n_4296);
  and g9093 (n5129, n_4295, n_4296);
  not g9094 (n_4297, n5128);
  not g9095 (n_4298, n5129);
  and g9096 (n5130, n_4297, n_4298);
  not g9097 (n_4299, n5130);
  and g9098 (n5131, n5119, n_4299);
  not g9099 (n_4300, n5119);
  and g9100 (n5132, n_4300, n5130);
  not g9101 (n_4301, n4964);
  not g9102 (n_4302, n5132);
  and g9103 (n5133, n_4301, n_4302);
  not g9104 (n_4303, n5131);
  and g9105 (n5134, n_4303, n5133);
  not g9106 (n_4304, n5134);
  and g9107 (n5135, n_4301, n_4304);
  and g9108 (n5136, n_4303, n_4304);
  and g9109 (n5137, n_4302, n5136);
  not g9110 (n_4305, n5135);
  not g9111 (n_4306, n5137);
  and g9112 (n5138, n_4305, n_4306);
  and g9113 (n5139, \b[28] , n700);
  and g9114 (n5140, \b[26] , n767);
  and g9115 (n5141, \b[27] , n695);
  and g9121 (n5144, n703, n3189);
  not g9124 (n_4311, n5145);
  and g9125 (n5146, \a[11] , n_4311);
  not g9126 (n_4312, n5146);
  and g9127 (n5147, \a[11] , n_4312);
  and g9128 (n5148, n_4311, n_4312);
  not g9129 (n_4313, n5147);
  not g9130 (n_4314, n5148);
  and g9131 (n5149, n_4313, n_4314);
  and g9132 (n5150, n5138, n5149);
  not g9133 (n_4315, n5138);
  not g9134 (n_4316, n5149);
  and g9135 (n5151, n_4315, n_4316);
  not g9136 (n_4317, n5150);
  not g9137 (n_4318, n5151);
  and g9138 (n5152, n_4317, n_4318);
  not g9139 (n_4319, n4963);
  and g9140 (n5153, n_4319, n5152);
  not g9141 (n_4320, n5152);
  and g9142 (n5154, n4963, n_4320);
  not g9143 (n_4321, n5153);
  not g9144 (n_4322, n5154);
  and g9145 (n5155, n_4321, n_4322);
  not g9146 (n_4323, n5155);
  and g9147 (n5156, n4961, n_4323);
  not g9148 (n_4324, n4961);
  and g9149 (n5157, n_4324, n5155);
  not g9150 (n_4325, n5156);
  not g9151 (n_4326, n5157);
  and g9152 (n5158, n_4325, n_4326);
  not g9153 (n_4327, n4950);
  and g9154 (n5159, n_4327, n5158);
  not g9155 (n_4328, n5158);
  and g9156 (n5160, n4950, n_4328);
  not g9157 (n_4329, n5159);
  not g9158 (n_4330, n5160);
  and g9159 (n5161, n_4329, n_4330);
  not g9160 (n_4331, n4949);
  and g9161 (n5162, n_4331, n5161);
  not g9162 (n_4332, n5162);
  and g9163 (n5163, n5161, n_4332);
  and g9164 (n5164, n_4331, n_4332);
  not g9165 (n_4333, n5163);
  not g9166 (n_4334, n5164);
  and g9167 (n5165, n_4333, n_4334);
  and g9168 (n5166, n_4106, n_4110);
  and g9169 (n5167, n5165, n5166);
  not g9170 (n_4335, n5165);
  not g9171 (n_4336, n5166);
  and g9172 (n5168, n_4335, n_4336);
  not g9173 (n_4337, n5167);
  not g9174 (n_4338, n5168);
  and g9175 (n5169, n_4337, n_4338);
  and g9176 (n5170, \b[37] , n266);
  and g9177 (n5171, \b[35] , n284);
  and g9178 (n5172, \b[36] , n261);
  and g9184 (n5175, n_4118, n_4121);
  not g9185 (n_4343, \b[37] );
  and g9186 (n5176, n_4116, n_4343);
  and g9187 (n5177, \b[36] , \b[37] );
  not g9188 (n_4344, n5176);
  not g9189 (n_4345, n5177);
  and g9190 (n5178, n_4344, n_4345);
  not g9191 (n_4346, n5175);
  and g9192 (n5179, n_4346, n5178);
  not g9193 (n_4347, n5178);
  and g9194 (n5180, n5175, n_4347);
  not g9195 (n_4348, n5179);
  not g9196 (n_4349, n5180);
  and g9197 (n5181, n_4348, n_4349);
  and g9198 (n5182, n269, n5181);
  not g9201 (n_4351, n5183);
  and g9202 (n5184, \a[2] , n_4351);
  not g9203 (n_4352, n5184);
  and g9204 (n5185, \a[2] , n_4352);
  and g9205 (n5186, n_4351, n_4352);
  not g9206 (n_4353, n5185);
  not g9207 (n_4354, n5186);
  and g9208 (n5187, n_4353, n_4354);
  not g9209 (n_4355, n5169);
  and g9210 (n5188, n_4355, n5187);
  not g9211 (n_4356, n5187);
  and g9212 (n5189, n5169, n_4356);
  not g9213 (n_4357, n5188);
  not g9214 (n_4358, n5189);
  and g9215 (n5190, n_4357, n_4358);
  not g9216 (n_4359, n4938);
  and g9217 (n5191, n_4359, n5190);
  not g9218 (n_4360, n5190);
  and g9219 (n5192, n4938, n_4360);
  not g9220 (n_4361, n5191);
  not g9221 (n_4362, n5192);
  and g9222 (\f[37] , n_4361, n_4362);
  and g9223 (n5194, \b[38] , n266);
  and g9224 (n5195, \b[36] , n284);
  and g9225 (n5196, \b[37] , n261);
  and g9231 (n5199, n_4345, n_4348);
  not g9232 (n_4367, \b[38] );
  and g9233 (n5200, n_4343, n_4367);
  and g9234 (n5201, \b[37] , \b[38] );
  not g9235 (n_4368, n5200);
  not g9236 (n_4369, n5201);
  and g9237 (n5202, n_4368, n_4369);
  not g9238 (n_4370, n5199);
  and g9239 (n5203, n_4370, n5202);
  not g9240 (n_4371, n5202);
  and g9241 (n5204, n5199, n_4371);
  not g9242 (n_4372, n5203);
  not g9243 (n_4373, n5204);
  and g9244 (n5205, n_4372, n_4373);
  and g9245 (n5206, n269, n5205);
  not g9248 (n_4375, n5207);
  and g9249 (n5208, \a[2] , n_4375);
  not g9250 (n_4376, n5208);
  and g9251 (n5209, \a[2] , n_4376);
  and g9252 (n5210, n_4375, n_4376);
  not g9253 (n_4377, n5209);
  not g9254 (n_4378, n5210);
  and g9255 (n5211, n_4377, n_4378);
  and g9256 (n5212, n_4332, n_4338);
  and g9257 (n5213, \b[35] , n362);
  and g9258 (n5214, \b[33] , n403);
  and g9259 (n5215, \b[34] , n357);
  and g9265 (n5218, n365, n4696);
  not g9268 (n_4383, n5219);
  and g9269 (n5220, \a[5] , n_4383);
  not g9270 (n_4384, n5220);
  and g9271 (n5221, \a[5] , n_4384);
  and g9272 (n5222, n_4383, n_4384);
  not g9273 (n_4385, n5221);
  not g9274 (n_4386, n5222);
  and g9275 (n5223, n_4385, n_4386);
  and g9276 (n5224, n_4326, n_4329);
  and g9277 (n5225, \b[32] , n511);
  and g9278 (n5226, \b[30] , n541);
  and g9279 (n5227, \b[31] , n506);
  and g9285 (n5230, n514, n4013);
  not g9288 (n_4391, n5231);
  and g9289 (n5232, \a[8] , n_4391);
  not g9290 (n_4392, n5232);
  and g9291 (n5233, \a[8] , n_4392);
  and g9292 (n5234, n_4391, n_4392);
  not g9293 (n_4393, n5233);
  not g9294 (n_4394, n5234);
  and g9295 (n5235, n_4393, n_4394);
  and g9296 (n5236, n_4318, n_4321);
  and g9297 (n5237, \b[29] , n700);
  and g9298 (n5238, \b[27] , n767);
  and g9299 (n5239, \b[28] , n695);
  and g9305 (n5242, n703, n3383);
  not g9308 (n_4399, n5243);
  and g9309 (n5244, \a[11] , n_4399);
  not g9310 (n_4400, n5244);
  and g9311 (n5245, \a[11] , n_4400);
  and g9312 (n5246, n_4399, n_4400);
  not g9313 (n_4401, n5245);
  not g9314 (n_4402, n5246);
  and g9315 (n5247, n_4401, n_4402);
  and g9316 (n5248, n_4283, n_4290);
  and g9317 (n5249, \b[17] , n2048);
  and g9318 (n5250, \b[15] , n2198);
  and g9319 (n5251, \b[16] , n2043);
  and g9325 (n5254, n1356, n2051);
  not g9328 (n_4407, n5255);
  and g9329 (n5256, \a[23] , n_4407);
  not g9330 (n_4408, n5256);
  and g9331 (n5257, \a[23] , n_4408);
  and g9332 (n5258, n_4407, n_4408);
  not g9333 (n_4409, n5257);
  not g9334 (n_4410, n5258);
  and g9335 (n5259, n_4409, n_4410);
  and g9336 (n5260, n_4244, n_4247);
  and g9337 (n5261, n_4236, n_4239);
  and g9338 (n5262, \b[11] , n3050);
  and g9339 (n5263, \b[9] , n3243);
  and g9340 (n5264, \b[10] , n3045);
  and g9346 (n5267, n818, n3053);
  not g9349 (n_4415, n5268);
  and g9350 (n5269, \a[29] , n_4415);
  not g9351 (n_4416, n5269);
  and g9352 (n5270, \a[29] , n_4416);
  and g9353 (n5271, n_4415, n_4416);
  not g9354 (n_4417, n5270);
  not g9355 (n_4418, n5271);
  and g9356 (n5272, n_4417, n_4418);
  and g9357 (n5273, n_4228, n_4231);
  and g9358 (n5274, n_4220, n_4223);
  and g9359 (n5275, \b[2] , n5035);
  and g9360 (n5276, n4761, n_4207);
  and g9361 (n5277, n5029, n5276);
  and g9362 (n5278, \b[0] , n5277);
  and g9363 (n5279, \b[1] , n5030);
  and g9369 (n5282, n296, n5038);
  not g9372 (n_4423, n5283);
  and g9373 (n5284, \a[38] , n_4423);
  not g9374 (n_4424, n5284);
  and g9375 (n5285, \a[38] , n_4424);
  and g9376 (n5286, n_4423, n_4424);
  not g9377 (n_4425, n5285);
  not g9378 (n_4426, n5286);
  and g9379 (n5287, n_4425, n_4426);
  and g9380 (n5288, n_4215, n5287);
  not g9381 (n_4427, n5287);
  and g9382 (n5289, n5045, n_4427);
  not g9383 (n_4428, n5288);
  not g9384 (n_4429, n5289);
  and g9385 (n5290, n_4428, n_4429);
  and g9386 (n5291, \b[5] , n4287);
  and g9387 (n5292, \b[3] , n4532);
  and g9388 (n5293, \b[4] , n4282);
  and g9394 (n5296, n394, n4290);
  not g9397 (n_4434, n5297);
  and g9398 (n5298, \a[35] , n_4434);
  not g9399 (n_4435, n5298);
  and g9400 (n5299, \a[35] , n_4435);
  and g9401 (n5300, n_4434, n_4435);
  not g9402 (n_4436, n5299);
  not g9403 (n_4437, n5300);
  and g9404 (n5301, n_4436, n_4437);
  not g9405 (n_4438, n5301);
  and g9406 (n5302, n5290, n_4438);
  not g9407 (n_4439, n5302);
  and g9408 (n5303, n5290, n_4439);
  and g9409 (n5304, n_4438, n_4439);
  not g9410 (n_4440, n5303);
  not g9411 (n_4441, n5304);
  and g9412 (n5305, n_4440, n_4441);
  not g9413 (n_4442, n5274);
  and g9414 (n5306, n_4442, n5305);
  not g9415 (n_4443, n5305);
  and g9416 (n5307, n5274, n_4443);
  not g9417 (n_4444, n5306);
  not g9418 (n_4445, n5307);
  and g9419 (n5308, n_4444, n_4445);
  and g9420 (n5309, \b[8] , n3638);
  and g9421 (n5310, \b[6] , n3843);
  and g9422 (n5311, \b[7] , n3633);
  and g9428 (n5314, n585, n3641);
  not g9431 (n_4450, n5315);
  and g9432 (n5316, \a[32] , n_4450);
  not g9433 (n_4451, n5316);
  and g9434 (n5317, \a[32] , n_4451);
  and g9435 (n5318, n_4450, n_4451);
  not g9436 (n_4452, n5317);
  not g9437 (n_4453, n5318);
  and g9438 (n5319, n_4452, n_4453);
  not g9439 (n_4454, n5308);
  not g9440 (n_4455, n5319);
  and g9441 (n5320, n_4454, n_4455);
  and g9442 (n5321, n5308, n5319);
  not g9443 (n_4456, n5320);
  not g9444 (n_4457, n5321);
  and g9445 (n5322, n_4456, n_4457);
  not g9446 (n_4458, n5273);
  and g9447 (n5323, n_4458, n5322);
  not g9448 (n_4459, n5322);
  and g9449 (n5324, n5273, n_4459);
  not g9450 (n_4460, n5323);
  not g9451 (n_4461, n5324);
  and g9452 (n5325, n_4460, n_4461);
  not g9453 (n_4462, n5272);
  and g9454 (n5326, n_4462, n5325);
  not g9455 (n_4463, n5326);
  and g9456 (n5327, n_4462, n_4463);
  and g9457 (n5328, n5325, n_4463);
  not g9458 (n_4464, n5327);
  not g9459 (n_4465, n5328);
  and g9460 (n5329, n_4464, n_4465);
  not g9461 (n_4466, n5261);
  not g9462 (n_4467, n5329);
  and g9463 (n5330, n_4466, n_4467);
  not g9464 (n_4468, n5330);
  and g9465 (n5331, n_4466, n_4468);
  and g9466 (n5332, n_4467, n_4468);
  not g9467 (n_4469, n5331);
  not g9468 (n_4470, n5332);
  and g9469 (n5333, n_4469, n_4470);
  and g9470 (n5334, \b[14] , n2539);
  and g9471 (n5335, \b[12] , n2685);
  and g9472 (n5336, \b[13] , n2534);
  and g9478 (n5339, n1034, n2542);
  not g9481 (n_4475, n5340);
  and g9482 (n5341, \a[26] , n_4475);
  not g9483 (n_4476, n5341);
  and g9484 (n5342, \a[26] , n_4476);
  and g9485 (n5343, n_4475, n_4476);
  not g9486 (n_4477, n5342);
  not g9487 (n_4478, n5343);
  and g9488 (n5344, n_4477, n_4478);
  and g9489 (n5345, n5333, n5344);
  not g9490 (n_4479, n5333);
  not g9491 (n_4480, n5344);
  and g9492 (n5346, n_4479, n_4480);
  not g9493 (n_4481, n5345);
  not g9494 (n_4482, n5346);
  and g9495 (n5347, n_4481, n_4482);
  not g9496 (n_4483, n5260);
  and g9497 (n5348, n_4483, n5347);
  not g9498 (n_4484, n5347);
  and g9499 (n5349, n5260, n_4484);
  not g9500 (n_4485, n5348);
  not g9501 (n_4486, n5349);
  and g9502 (n5350, n_4485, n_4486);
  not g9503 (n_4487, n5259);
  and g9504 (n5351, n_4487, n5350);
  not g9505 (n_4488, n5351);
  and g9506 (n5352, n5350, n_4488);
  and g9507 (n5353, n_4487, n_4488);
  not g9508 (n_4489, n5352);
  not g9509 (n_4490, n5353);
  and g9510 (n5354, n_4489, n_4490);
  and g9511 (n5355, n_4250, n_4257);
  and g9512 (n5356, n5354, n5355);
  not g9513 (n_4491, n5354);
  not g9514 (n_4492, n5355);
  and g9515 (n5357, n_4491, n_4492);
  not g9516 (n_4493, n5356);
  not g9517 (n_4494, n5357);
  and g9518 (n5358, n_4493, n_4494);
  and g9519 (n5359, \b[20] , n1627);
  and g9520 (n5360, \b[18] , n1763);
  and g9521 (n5361, \b[19] , n1622);
  and g9527 (n5364, n1630, n1846);
  not g9530 (n_4499, n5365);
  and g9531 (n5366, \a[20] , n_4499);
  not g9532 (n_4500, n5366);
  and g9533 (n5367, \a[20] , n_4500);
  and g9534 (n5368, n_4499, n_4500);
  not g9535 (n_4501, n5367);
  not g9536 (n_4502, n5368);
  and g9537 (n5369, n_4501, n_4502);
  not g9538 (n_4503, n5369);
  and g9539 (n5370, n5358, n_4503);
  not g9540 (n_4504, n5370);
  and g9541 (n5371, n5358, n_4504);
  and g9542 (n5372, n_4503, n_4504);
  not g9543 (n_4505, n5371);
  not g9544 (n_4506, n5372);
  and g9545 (n5373, n_4505, n_4506);
  and g9546 (n5374, n_4267, n_4273);
  and g9547 (n5375, n5373, n5374);
  not g9548 (n_4507, n5373);
  not g9549 (n_4508, n5374);
  and g9550 (n5376, n_4507, n_4508);
  not g9551 (n_4509, n5375);
  not g9552 (n_4510, n5376);
  and g9553 (n5377, n_4509, n_4510);
  and g9554 (n5378, \b[23] , n1302);
  and g9555 (n5379, \b[21] , n1391);
  and g9556 (n5380, \b[22] , n1297);
  and g9562 (n5383, n1305, n2300);
  not g9565 (n_4515, n5384);
  and g9566 (n5385, \a[17] , n_4515);
  not g9567 (n_4516, n5385);
  and g9568 (n5386, \a[17] , n_4516);
  and g9569 (n5387, n_4515, n_4516);
  not g9570 (n_4517, n5386);
  not g9571 (n_4518, n5387);
  and g9572 (n5388, n_4517, n_4518);
  not g9573 (n_4519, n5388);
  and g9574 (n5389, n5377, n_4519);
  not g9575 (n_4520, n5377);
  and g9576 (n5390, n_4520, n5388);
  not g9577 (n_4521, n5248);
  not g9578 (n_4522, n5390);
  and g9579 (n5391, n_4521, n_4522);
  not g9580 (n_4523, n5389);
  and g9581 (n5392, n_4523, n5391);
  not g9582 (n_4524, n5392);
  and g9583 (n5393, n_4521, n_4524);
  and g9584 (n5394, n_4523, n_4524);
  and g9585 (n5395, n_4522, n5394);
  not g9586 (n_4525, n5393);
  not g9587 (n_4526, n5395);
  and g9588 (n5396, n_4525, n_4526);
  and g9589 (n5397, \b[26] , n951);
  and g9590 (n5398, \b[24] , n1056);
  and g9591 (n5399, \b[25] , n946);
  and g9597 (n5402, n954, n2813);
  not g9600 (n_4531, n5403);
  and g9601 (n5404, \a[14] , n_4531);
  not g9602 (n_4532, n5404);
  and g9603 (n5405, \a[14] , n_4532);
  and g9604 (n5406, n_4531, n_4532);
  not g9605 (n_4533, n5405);
  not g9606 (n_4534, n5406);
  and g9607 (n5407, n_4533, n_4534);
  and g9608 (n5408, n5396, n5407);
  not g9609 (n_4535, n5396);
  not g9610 (n_4536, n5407);
  and g9611 (n5409, n_4535, n_4536);
  not g9612 (n_4537, n5408);
  not g9613 (n_4538, n5409);
  and g9614 (n5410, n_4537, n_4538);
  not g9615 (n_4539, n5136);
  and g9616 (n5411, n_4539, n5410);
  not g9617 (n_4540, n5410);
  and g9618 (n5412, n5136, n_4540);
  not g9619 (n_4541, n5411);
  not g9620 (n_4542, n5412);
  and g9621 (n5413, n_4541, n_4542);
  not g9622 (n_4543, n5413);
  and g9623 (n5414, n5247, n_4543);
  not g9624 (n_4544, n5247);
  and g9625 (n5415, n_4544, n5413);
  not g9626 (n_4545, n5414);
  not g9627 (n_4546, n5415);
  and g9628 (n5416, n_4545, n_4546);
  not g9629 (n_4547, n5236);
  and g9630 (n5417, n_4547, n5416);
  not g9631 (n_4548, n5416);
  and g9632 (n5418, n5236, n_4548);
  not g9633 (n_4549, n5417);
  not g9634 (n_4550, n5418);
  and g9635 (n5419, n_4549, n_4550);
  not g9636 (n_4551, n5419);
  and g9637 (n5420, n5235, n_4551);
  not g9638 (n_4552, n5235);
  and g9639 (n5421, n_4552, n5419);
  not g9640 (n_4553, n5420);
  not g9641 (n_4554, n5421);
  and g9642 (n5422, n_4553, n_4554);
  not g9643 (n_4555, n5224);
  and g9644 (n5423, n_4555, n5422);
  not g9645 (n_4556, n5422);
  and g9646 (n5424, n5224, n_4556);
  not g9647 (n_4557, n5423);
  not g9648 (n_4558, n5424);
  and g9649 (n5425, n_4557, n_4558);
  not g9650 (n_4559, n5425);
  and g9651 (n5426, n5223, n_4559);
  not g9652 (n_4560, n5223);
  and g9653 (n5427, n_4560, n5425);
  not g9654 (n_4561, n5426);
  not g9655 (n_4562, n5427);
  and g9656 (n5428, n_4561, n_4562);
  not g9657 (n_4563, n5212);
  and g9658 (n5429, n_4563, n5428);
  not g9659 (n_4564, n5428);
  and g9660 (n5430, n5212, n_4564);
  not g9661 (n_4565, n5429);
  not g9662 (n_4566, n5430);
  and g9663 (n5431, n_4565, n_4566);
  not g9664 (n_4567, n5211);
  and g9665 (n5432, n_4567, n5431);
  not g9666 (n_4568, n5432);
  and g9667 (n5433, n5431, n_4568);
  and g9668 (n5434, n_4567, n_4568);
  not g9669 (n_4569, n5433);
  not g9670 (n_4570, n5434);
  and g9671 (n5435, n_4569, n_4570);
  and g9672 (n5436, n_4358, n_4361);
  not g9673 (n_4571, n5435);
  not g9674 (n_4572, n5436);
  and g9675 (n5437, n_4571, n_4572);
  and g9676 (n5438, n5435, n5436);
  not g9677 (n_4573, n5437);
  not g9678 (n_4574, n5438);
  and g9679 (\f[38] , n_4573, n_4574);
  and g9680 (n5440, \b[39] , n266);
  and g9681 (n5441, \b[37] , n284);
  and g9682 (n5442, \b[38] , n261);
  and g9688 (n5445, n_4369, n_4372);
  not g9689 (n_4579, \b[39] );
  and g9690 (n5446, n_4367, n_4579);
  and g9691 (n5447, \b[38] , \b[39] );
  not g9692 (n_4580, n5446);
  not g9693 (n_4581, n5447);
  and g9694 (n5448, n_4580, n_4581);
  not g9695 (n_4582, n5445);
  and g9696 (n5449, n_4582, n5448);
  not g9697 (n_4583, n5448);
  and g9698 (n5450, n5445, n_4583);
  not g9699 (n_4584, n5449);
  not g9700 (n_4585, n5450);
  and g9701 (n5451, n_4584, n_4585);
  and g9702 (n5452, n269, n5451);
  not g9705 (n_4587, n5453);
  and g9706 (n5454, \a[2] , n_4587);
  not g9707 (n_4588, n5454);
  and g9708 (n5455, \a[2] , n_4588);
  and g9709 (n5456, n_4587, n_4588);
  not g9710 (n_4589, n5455);
  not g9711 (n_4590, n5456);
  and g9712 (n5457, n_4589, n_4590);
  and g9713 (n5458, n_4562, n_4565);
  and g9714 (n5459, n_4554, n_4557);
  and g9715 (n5460, \b[33] , n511);
  and g9716 (n5461, \b[31] , n541);
  and g9717 (n5462, \b[32] , n506);
  and g9723 (n5465, n514, n4223);
  not g9726 (n_4595, n5466);
  and g9727 (n5467, \a[8] , n_4595);
  not g9728 (n_4596, n5467);
  and g9729 (n5468, \a[8] , n_4596);
  and g9730 (n5469, n_4595, n_4596);
  not g9731 (n_4597, n5468);
  not g9732 (n_4598, n5469);
  and g9733 (n5470, n_4597, n_4598);
  and g9734 (n5471, n_4546, n_4549);
  and g9735 (n5472, n_4538, n_4541);
  and g9736 (n5473, \b[27] , n951);
  and g9737 (n5474, \b[25] , n1056);
  and g9738 (n5475, \b[26] , n946);
  and g9744 (n5478, n954, n2990);
  not g9747 (n_4603, n5479);
  and g9748 (n5480, \a[14] , n_4603);
  not g9749 (n_4604, n5480);
  and g9750 (n5481, \a[14] , n_4604);
  and g9751 (n5482, n_4603, n_4604);
  not g9752 (n_4605, n5481);
  not g9753 (n_4606, n5482);
  and g9754 (n5483, n_4605, n_4606);
  and g9755 (n5484, n_4488, n_4494);
  and g9756 (n5485, n_4482, n_4485);
  and g9757 (n5486, \b[15] , n2539);
  and g9758 (n5487, \b[13] , n2685);
  and g9759 (n5488, \b[14] , n2534);
  and g9765 (n5491, n1131, n2542);
  not g9768 (n_4611, n5492);
  and g9769 (n5493, \a[26] , n_4611);
  not g9770 (n_4612, n5493);
  and g9771 (n5494, \a[26] , n_4612);
  and g9772 (n5495, n_4611, n_4612);
  not g9773 (n_4613, n5494);
  not g9774 (n_4614, n5495);
  and g9775 (n5496, n_4613, n_4614);
  and g9776 (n5497, \b[6] , n4287);
  and g9777 (n5498, \b[4] , n4532);
  and g9778 (n5499, \b[5] , n4282);
  and g9784 (n5502, n459, n4290);
  not g9787 (n_4619, n5503);
  and g9788 (n5504, \a[35] , n_4619);
  not g9789 (n_4620, n5504);
  and g9790 (n5505, \a[35] , n_4620);
  and g9791 (n5506, n_4619, n_4620);
  not g9792 (n_4621, n5505);
  not g9793 (n_4622, n5506);
  and g9794 (n5507, n_4621, n_4622);
  not g9795 (n_4624, \a[39] );
  and g9796 (n5508, \a[38] , n_4624);
  and g9797 (n5509, n_4202, \a[39] );
  not g9798 (n_4625, n5508);
  not g9799 (n_4626, n5509);
  and g9800 (n5510, n_4625, n_4626);
  not g9801 (n_4627, n5510);
  and g9802 (n5511, \b[0] , n_4627);
  and g9803 (n5512, n_4429, n5511);
  not g9804 (n_4628, n5511);
  and g9805 (n5513, n5289, n_4628);
  not g9806 (n_4629, n5512);
  not g9807 (n_4630, n5513);
  and g9808 (n5514, n_4629, n_4630);
  and g9809 (n5515, \b[3] , n5035);
  and g9810 (n5516, \b[1] , n5277);
  and g9811 (n5517, \b[2] , n5030);
  and g9817 (n5520, n318, n5038);
  not g9820 (n_4635, n5521);
  and g9821 (n5522, \a[38] , n_4635);
  not g9822 (n_4636, n5522);
  and g9823 (n5523, \a[38] , n_4636);
  and g9824 (n5524, n_4635, n_4636);
  not g9825 (n_4637, n5523);
  not g9826 (n_4638, n5524);
  and g9827 (n5525, n_4637, n_4638);
  not g9828 (n_4639, n5514);
  not g9829 (n_4640, n5525);
  and g9830 (n5526, n_4639, n_4640);
  and g9831 (n5527, n5514, n5525);
  not g9832 (n_4641, n5526);
  not g9833 (n_4642, n5527);
  and g9834 (n5528, n_4641, n_4642);
  not g9835 (n_4643, n5507);
  and g9836 (n5529, n_4643, n5528);
  not g9837 (n_4644, n5529);
  and g9838 (n5530, n5528, n_4644);
  and g9839 (n5531, n_4643, n_4644);
  not g9840 (n_4645, n5530);
  not g9841 (n_4646, n5531);
  and g9842 (n5532, n_4645, n_4646);
  and g9843 (n5533, n_4442, n_4443);
  not g9844 (n_4647, n5533);
  and g9845 (n5534, n_4439, n_4647);
  and g9846 (n5535, n5532, n5534);
  not g9847 (n_4648, n5532);
  not g9848 (n_4649, n5534);
  and g9849 (n5536, n_4648, n_4649);
  not g9850 (n_4650, n5535);
  not g9851 (n_4651, n5536);
  and g9852 (n5537, n_4650, n_4651);
  and g9853 (n5538, \b[9] , n3638);
  and g9854 (n5539, \b[7] , n3843);
  and g9855 (n5540, \b[8] , n3633);
  and g9861 (n5543, n651, n3641);
  not g9864 (n_4656, n5544);
  and g9865 (n5545, \a[32] , n_4656);
  not g9866 (n_4657, n5545);
  and g9867 (n5546, \a[32] , n_4657);
  and g9868 (n5547, n_4656, n_4657);
  not g9869 (n_4658, n5546);
  not g9870 (n_4659, n5547);
  and g9871 (n5548, n_4658, n_4659);
  not g9872 (n_4660, n5548);
  and g9873 (n5549, n5537, n_4660);
  not g9874 (n_4661, n5549);
  and g9875 (n5550, n5537, n_4661);
  and g9876 (n5551, n_4660, n_4661);
  not g9877 (n_4662, n5550);
  not g9878 (n_4663, n5551);
  and g9879 (n5552, n_4662, n_4663);
  and g9880 (n5553, n_4456, n_4460);
  and g9881 (n5554, n5552, n5553);
  not g9882 (n_4664, n5552);
  not g9883 (n_4665, n5553);
  and g9884 (n5555, n_4664, n_4665);
  not g9885 (n_4666, n5554);
  not g9886 (n_4667, n5555);
  and g9887 (n5556, n_4666, n_4667);
  and g9888 (n5557, \b[12] , n3050);
  and g9889 (n5558, \b[10] , n3243);
  and g9890 (n5559, \b[11] , n3045);
  and g9896 (n5562, n842, n3053);
  not g9899 (n_4672, n5563);
  and g9900 (n5564, \a[29] , n_4672);
  not g9901 (n_4673, n5564);
  and g9902 (n5565, \a[29] , n_4673);
  and g9903 (n5566, n_4672, n_4673);
  not g9904 (n_4674, n5565);
  not g9905 (n_4675, n5566);
  and g9906 (n5567, n_4674, n_4675);
  not g9907 (n_4676, n5556);
  and g9908 (n5568, n_4676, n5567);
  not g9909 (n_4677, n5567);
  and g9910 (n5569, n5556, n_4677);
  not g9911 (n_4678, n5568);
  not g9912 (n_4679, n5569);
  and g9913 (n5570, n_4678, n_4679);
  and g9914 (n5571, n_4463, n_4468);
  not g9915 (n_4680, n5571);
  and g9916 (n5572, n5570, n_4680);
  not g9917 (n_4681, n5570);
  and g9918 (n5573, n_4681, n5571);
  not g9919 (n_4682, n5572);
  not g9920 (n_4683, n5573);
  and g9921 (n5574, n_4682, n_4683);
  not g9922 (n_4684, n5496);
  and g9923 (n5575, n_4684, n5574);
  not g9924 (n_4685, n5575);
  and g9925 (n5576, n5574, n_4685);
  and g9926 (n5577, n_4684, n_4685);
  not g9927 (n_4686, n5576);
  not g9928 (n_4687, n5577);
  and g9929 (n5578, n_4686, n_4687);
  not g9930 (n_4688, n5485);
  and g9931 (n5579, n_4688, n5578);
  not g9932 (n_4689, n5578);
  and g9933 (n5580, n5485, n_4689);
  not g9934 (n_4690, n5579);
  not g9935 (n_4691, n5580);
  and g9936 (n5581, n_4690, n_4691);
  and g9937 (n5582, \b[18] , n2048);
  and g9938 (n5583, \b[16] , n2198);
  and g9939 (n5584, \b[17] , n2043);
  and g9945 (n5587, n1566, n2051);
  not g9948 (n_4696, n5588);
  and g9949 (n5589, \a[23] , n_4696);
  not g9950 (n_4697, n5589);
  and g9951 (n5590, \a[23] , n_4697);
  and g9952 (n5591, n_4696, n_4697);
  not g9953 (n_4698, n5590);
  not g9954 (n_4699, n5591);
  and g9955 (n5592, n_4698, n_4699);
  not g9956 (n_4700, n5581);
  not g9957 (n_4701, n5592);
  and g9958 (n5593, n_4700, n_4701);
  and g9959 (n5594, n5581, n5592);
  not g9960 (n_4702, n5593);
  not g9961 (n_4703, n5594);
  and g9962 (n5595, n_4702, n_4703);
  not g9963 (n_4704, n5595);
  and g9964 (n5596, n5484, n_4704);
  not g9965 (n_4705, n5484);
  and g9966 (n5597, n_4705, n5595);
  not g9967 (n_4706, n5596);
  not g9968 (n_4707, n5597);
  and g9969 (n5598, n_4706, n_4707);
  and g9970 (n5599, \b[21] , n1627);
  and g9971 (n5600, \b[19] , n1763);
  and g9972 (n5601, \b[20] , n1622);
  and g9978 (n5604, n1630, n1984);
  not g9981 (n_4712, n5605);
  and g9982 (n5606, \a[20] , n_4712);
  not g9983 (n_4713, n5606);
  and g9984 (n5607, \a[20] , n_4713);
  and g9985 (n5608, n_4712, n_4713);
  not g9986 (n_4714, n5607);
  not g9987 (n_4715, n5608);
  and g9988 (n5609, n_4714, n_4715);
  not g9989 (n_4716, n5609);
  and g9990 (n5610, n5598, n_4716);
  not g9991 (n_4717, n5610);
  and g9992 (n5611, n5598, n_4717);
  and g9993 (n5612, n_4716, n_4717);
  not g9994 (n_4718, n5611);
  not g9995 (n_4719, n5612);
  and g9996 (n5613, n_4718, n_4719);
  and g9997 (n5614, n_4504, n_4510);
  and g9998 (n5615, n5613, n5614);
  not g9999 (n_4720, n5613);
  not g10000 (n_4721, n5614);
  and g10001 (n5616, n_4720, n_4721);
  not g10002 (n_4722, n5615);
  not g10003 (n_4723, n5616);
  and g10004 (n5617, n_4722, n_4723);
  and g10005 (n5618, \b[24] , n1302);
  and g10006 (n5619, \b[22] , n1391);
  and g10007 (n5620, \b[23] , n1297);
  and g10013 (n5623, n1305, n2458);
  not g10016 (n_4728, n5624);
  and g10017 (n5625, \a[17] , n_4728);
  not g10018 (n_4729, n5625);
  and g10019 (n5626, \a[17] , n_4729);
  and g10020 (n5627, n_4728, n_4729);
  not g10021 (n_4730, n5626);
  not g10022 (n_4731, n5627);
  and g10023 (n5628, n_4730, n_4731);
  not g10024 (n_4732, n5617);
  and g10025 (n5629, n_4732, n5628);
  not g10026 (n_4733, n5628);
  and g10027 (n5630, n5617, n_4733);
  not g10028 (n_4734, n5629);
  not g10029 (n_4735, n5630);
  and g10030 (n5631, n_4734, n_4735);
  not g10031 (n_4736, n5394);
  and g10032 (n5632, n_4736, n5631);
  not g10033 (n_4737, n5631);
  and g10034 (n5633, n5394, n_4737);
  not g10035 (n_4738, n5632);
  not g10036 (n_4739, n5633);
  and g10037 (n5634, n_4738, n_4739);
  not g10038 (n_4740, n5483);
  and g10039 (n5635, n_4740, n5634);
  not g10040 (n_4741, n5635);
  and g10041 (n5636, n5634, n_4741);
  and g10042 (n5637, n_4740, n_4741);
  not g10043 (n_4742, n5636);
  not g10044 (n_4743, n5637);
  and g10045 (n5638, n_4742, n_4743);
  not g10046 (n_4744, n5472);
  and g10047 (n5639, n_4744, n5638);
  not g10048 (n_4745, n5638);
  and g10049 (n5640, n5472, n_4745);
  not g10050 (n_4746, n5639);
  not g10051 (n_4747, n5640);
  and g10052 (n5641, n_4746, n_4747);
  and g10053 (n5642, \b[30] , n700);
  and g10054 (n5643, \b[28] , n767);
  and g10055 (n5644, \b[29] , n695);
  and g10061 (n5647, n703, n3577);
  not g10064 (n_4752, n5648);
  and g10065 (n5649, \a[11] , n_4752);
  not g10066 (n_4753, n5649);
  and g10067 (n5650, \a[11] , n_4753);
  and g10068 (n5651, n_4752, n_4753);
  not g10069 (n_4754, n5650);
  not g10070 (n_4755, n5651);
  and g10071 (n5652, n_4754, n_4755);
  not g10072 (n_4756, n5641);
  not g10073 (n_4757, n5652);
  and g10074 (n5653, n_4756, n_4757);
  and g10075 (n5654, n5641, n5652);
  not g10076 (n_4758, n5653);
  not g10077 (n_4759, n5654);
  and g10078 (n5655, n_4758, n_4759);
  not g10079 (n_4760, n5471);
  and g10080 (n5656, n_4760, n5655);
  not g10081 (n_4761, n5655);
  and g10082 (n5657, n5471, n_4761);
  not g10083 (n_4762, n5656);
  not g10084 (n_4763, n5657);
  and g10085 (n5658, n_4762, n_4763);
  not g10086 (n_4764, n5470);
  and g10087 (n5659, n_4764, n5658);
  not g10088 (n_4765, n5659);
  and g10089 (n5660, n5658, n_4765);
  and g10090 (n5661, n_4764, n_4765);
  not g10091 (n_4766, n5660);
  not g10092 (n_4767, n5661);
  and g10093 (n5662, n_4766, n_4767);
  not g10094 (n_4768, n5459);
  and g10095 (n5663, n_4768, n5662);
  not g10096 (n_4769, n5662);
  and g10097 (n5664, n5459, n_4769);
  not g10098 (n_4770, n5663);
  not g10099 (n_4771, n5664);
  and g10100 (n5665, n_4770, n_4771);
  and g10101 (n5666, \b[36] , n362);
  and g10102 (n5667, \b[34] , n403);
  and g10103 (n5668, \b[35] , n357);
  and g10109 (n5671, n365, n4922);
  not g10112 (n_4776, n5672);
  and g10113 (n5673, \a[5] , n_4776);
  not g10114 (n_4777, n5673);
  and g10115 (n5674, \a[5] , n_4777);
  and g10116 (n5675, n_4776, n_4777);
  not g10117 (n_4778, n5674);
  not g10118 (n_4779, n5675);
  and g10119 (n5676, n_4778, n_4779);
  and g10120 (n5677, n5665, n5676);
  not g10121 (n_4780, n5665);
  not g10122 (n_4781, n5676);
  and g10123 (n5678, n_4780, n_4781);
  not g10124 (n_4782, n5677);
  not g10125 (n_4783, n5678);
  and g10126 (n5679, n_4782, n_4783);
  not g10127 (n_4784, n5458);
  and g10128 (n5680, n_4784, n5679);
  not g10129 (n_4785, n5679);
  and g10130 (n5681, n5458, n_4785);
  not g10131 (n_4786, n5680);
  not g10132 (n_4787, n5681);
  and g10133 (n5682, n_4786, n_4787);
  not g10134 (n_4788, n5457);
  and g10135 (n5683, n_4788, n5682);
  not g10136 (n_4789, n5683);
  and g10137 (n5684, n5682, n_4789);
  and g10138 (n5685, n_4788, n_4789);
  not g10139 (n_4790, n5684);
  not g10140 (n_4791, n5685);
  and g10141 (n5686, n_4790, n_4791);
  and g10142 (n5687, n_4568, n_4573);
  not g10143 (n_4792, n5686);
  not g10144 (n_4793, n5687);
  and g10145 (n5688, n_4792, n_4793);
  and g10146 (n5689, n5686, n5687);
  not g10147 (n_4794, n5688);
  not g10148 (n_4795, n5689);
  and g10149 (\f[39] , n_4794, n_4795);
  and g10150 (n5691, n_4789, n_4794);
  and g10151 (n5692, n_4783, n_4786);
  and g10152 (n5693, \b[37] , n362);
  and g10153 (n5694, \b[35] , n403);
  and g10154 (n5695, \b[36] , n357);
  and g10160 (n5698, n365, n5181);
  not g10163 (n_4800, n5699);
  and g10164 (n5700, \a[5] , n_4800);
  not g10165 (n_4801, n5700);
  and g10166 (n5701, \a[5] , n_4801);
  and g10167 (n5702, n_4800, n_4801);
  not g10168 (n_4802, n5701);
  not g10169 (n_4803, n5702);
  and g10170 (n5703, n_4802, n_4803);
  and g10171 (n5704, n_4768, n_4769);
  not g10172 (n_4804, n5704);
  and g10173 (n5705, n_4765, n_4804);
  and g10174 (n5706, \b[34] , n511);
  and g10175 (n5707, \b[32] , n541);
  and g10176 (n5708, \b[33] , n506);
  and g10182 (n5711, n514, n4466);
  not g10185 (n_4809, n5712);
  and g10186 (n5713, \a[8] , n_4809);
  not g10187 (n_4810, n5713);
  and g10188 (n5714, \a[8] , n_4810);
  and g10189 (n5715, n_4809, n_4810);
  not g10190 (n_4811, n5714);
  not g10191 (n_4812, n5715);
  and g10192 (n5716, n_4811, n_4812);
  and g10193 (n5717, n_4758, n_4762);
  and g10194 (n5718, n_4744, n_4745);
  not g10195 (n_4813, n5718);
  and g10196 (n5719, n_4741, n_4813);
  and g10197 (n5720, \b[28] , n951);
  and g10198 (n5721, \b[26] , n1056);
  and g10199 (n5722, \b[27] , n946);
  and g10205 (n5725, n954, n3189);
  not g10208 (n_4818, n5726);
  and g10209 (n5727, \a[14] , n_4818);
  not g10210 (n_4819, n5727);
  and g10211 (n5728, \a[14] , n_4819);
  and g10212 (n5729, n_4818, n_4819);
  not g10213 (n_4820, n5728);
  not g10214 (n_4821, n5729);
  and g10215 (n5730, n_4820, n_4821);
  and g10216 (n5731, \b[16] , n2539);
  and g10217 (n5732, \b[14] , n2685);
  and g10218 (n5733, \b[15] , n2534);
  and g10224 (n5736, n1237, n2542);
  not g10227 (n_4826, n5737);
  and g10228 (n5738, \a[26] , n_4826);
  not g10229 (n_4827, n5738);
  and g10230 (n5739, \a[26] , n_4827);
  and g10231 (n5740, n_4826, n_4827);
  not g10232 (n_4828, n5739);
  not g10233 (n_4829, n5740);
  and g10234 (n5741, n_4828, n_4829);
  and g10235 (n5742, n_4679, n_4682);
  and g10236 (n5743, n_4661, n_4667);
  and g10237 (n5744, \b[7] , n4287);
  and g10238 (n5745, \b[5] , n4532);
  and g10239 (n5746, \b[6] , n4282);
  and g10245 (n5749, n484, n4290);
  not g10248 (n_4834, n5750);
  and g10249 (n5751, \a[35] , n_4834);
  not g10250 (n_4835, n5751);
  and g10251 (n5752, \a[35] , n_4835);
  and g10252 (n5753, n_4834, n_4835);
  not g10253 (n_4836, n5752);
  not g10254 (n_4837, n5753);
  and g10255 (n5754, n_4836, n_4837);
  and g10256 (n5755, n5289, n5511);
  not g10257 (n_4838, n5755);
  and g10258 (n5756, n_4641, n_4838);
  and g10259 (n5757, \b[4] , n5035);
  and g10260 (n5758, \b[2] , n5277);
  and g10261 (n5759, \b[3] , n5030);
  and g10267 (n5762, n346, n5038);
  not g10270 (n_4843, n5763);
  and g10271 (n5764, \a[38] , n_4843);
  not g10272 (n_4844, n5764);
  and g10273 (n5765, \a[38] , n_4844);
  and g10274 (n5766, n_4843, n_4844);
  not g10275 (n_4845, n5765);
  not g10276 (n_4846, n5766);
  and g10277 (n5767, n_4845, n_4846);
  and g10278 (n5768, \a[41] , n_4628);
  and g10279 (n5769, n_4624, \a[40] );
  not g10280 (n_4849, \a[40] );
  and g10281 (n5770, \a[39] , n_4849);
  not g10282 (n_4850, n5769);
  not g10283 (n_4851, n5770);
  and g10284 (n5771, n_4850, n_4851);
  not g10285 (n_4852, n5771);
  and g10286 (n5772, n5510, n_4852);
  and g10287 (n5773, \b[0] , n5772);
  and g10288 (n5774, n_4849, \a[41] );
  not g10289 (n_4853, \a[41] );
  and g10290 (n5775, \a[40] , n_4853);
  not g10291 (n_4854, n5774);
  not g10292 (n_4855, n5775);
  and g10293 (n5776, n_4854, n_4855);
  and g10294 (n5777, n_4627, n5776);
  and g10295 (n5778, \b[1] , n5777);
  not g10296 (n_4856, n5773);
  not g10297 (n_4857, n5778);
  and g10298 (n5779, n_4856, n_4857);
  not g10299 (n_4858, n5776);
  and g10300 (n5780, n_4627, n_4858);
  and g10301 (n5781, n_21, n5780);
  not g10302 (n_4859, n5781);
  and g10303 (n5782, n5779, n_4859);
  not g10304 (n_4860, n5782);
  and g10305 (n5783, \a[41] , n_4860);
  not g10306 (n_4861, n5783);
  and g10307 (n5784, \a[41] , n_4861);
  and g10308 (n5785, n_4860, n_4861);
  not g10309 (n_4862, n5784);
  not g10310 (n_4863, n5785);
  and g10311 (n5786, n_4862, n_4863);
  not g10312 (n_4864, n5786);
  and g10313 (n5787, n5768, n_4864);
  not g10314 (n_4865, n5768);
  and g10315 (n5788, n_4865, n5786);
  not g10316 (n_4866, n5787);
  not g10317 (n_4867, n5788);
  and g10318 (n5789, n_4866, n_4867);
  not g10319 (n_4868, n5789);
  and g10320 (n5790, n5767, n_4868);
  not g10321 (n_4869, n5767);
  and g10322 (n5791, n_4869, n5789);
  not g10323 (n_4870, n5790);
  not g10324 (n_4871, n5791);
  and g10325 (n5792, n_4870, n_4871);
  not g10326 (n_4872, n5756);
  and g10327 (n5793, n_4872, n5792);
  not g10328 (n_4873, n5792);
  and g10329 (n5794, n5756, n_4873);
  not g10330 (n_4874, n5793);
  not g10331 (n_4875, n5794);
  and g10332 (n5795, n_4874, n_4875);
  not g10333 (n_4876, n5754);
  and g10334 (n5796, n_4876, n5795);
  not g10335 (n_4877, n5796);
  and g10336 (n5797, n5795, n_4877);
  and g10337 (n5798, n_4876, n_4877);
  not g10338 (n_4878, n5797);
  not g10339 (n_4879, n5798);
  and g10340 (n5799, n_4878, n_4879);
  and g10341 (n5800, n_4644, n_4651);
  and g10342 (n5801, n5799, n5800);
  not g10343 (n_4880, n5799);
  not g10344 (n_4881, n5800);
  and g10345 (n5802, n_4880, n_4881);
  not g10346 (n_4882, n5801);
  not g10347 (n_4883, n5802);
  and g10348 (n5803, n_4882, n_4883);
  and g10349 (n5804, \b[10] , n3638);
  and g10350 (n5805, \b[8] , n3843);
  and g10351 (n5806, \b[9] , n3633);
  and g10357 (n5809, n738, n3641);
  not g10360 (n_4888, n5810);
  and g10361 (n5811, \a[32] , n_4888);
  not g10362 (n_4889, n5811);
  and g10363 (n5812, \a[32] , n_4889);
  and g10364 (n5813, n_4888, n_4889);
  not g10365 (n_4890, n5812);
  not g10366 (n_4891, n5813);
  and g10367 (n5814, n_4890, n_4891);
  not g10368 (n_4892, n5814);
  and g10369 (n5815, n5803, n_4892);
  not g10370 (n_4893, n5803);
  and g10371 (n5816, n_4893, n5814);
  not g10372 (n_4894, n5743);
  not g10373 (n_4895, n5816);
  and g10374 (n5817, n_4894, n_4895);
  not g10375 (n_4896, n5815);
  and g10376 (n5818, n_4896, n5817);
  not g10377 (n_4897, n5818);
  and g10378 (n5819, n_4894, n_4897);
  and g10379 (n5820, n_4896, n_4897);
  and g10380 (n5821, n_4895, n5820);
  not g10381 (n_4898, n5819);
  not g10382 (n_4899, n5821);
  and g10383 (n5822, n_4898, n_4899);
  and g10384 (n5823, \b[13] , n3050);
  and g10385 (n5824, \b[11] , n3243);
  and g10386 (n5825, \b[12] , n3045);
  and g10392 (n5828, n1008, n3053);
  not g10395 (n_4904, n5829);
  and g10396 (n5830, \a[29] , n_4904);
  not g10397 (n_4905, n5830);
  and g10398 (n5831, \a[29] , n_4905);
  and g10399 (n5832, n_4904, n_4905);
  not g10400 (n_4906, n5831);
  not g10401 (n_4907, n5832);
  and g10402 (n5833, n_4906, n_4907);
  and g10403 (n5834, n5822, n5833);
  not g10404 (n_4908, n5822);
  not g10405 (n_4909, n5833);
  and g10406 (n5835, n_4908, n_4909);
  not g10407 (n_4910, n5834);
  not g10408 (n_4911, n5835);
  and g10409 (n5836, n_4910, n_4911);
  not g10410 (n_4912, n5742);
  and g10411 (n5837, n_4912, n5836);
  not g10412 (n_4913, n5836);
  and g10413 (n5838, n5742, n_4913);
  not g10414 (n_4914, n5837);
  not g10415 (n_4915, n5838);
  and g10416 (n5839, n_4914, n_4915);
  not g10417 (n_4916, n5741);
  and g10418 (n5840, n_4916, n5839);
  not g10419 (n_4917, n5840);
  and g10420 (n5841, n5839, n_4917);
  and g10421 (n5842, n_4916, n_4917);
  not g10422 (n_4918, n5841);
  not g10423 (n_4919, n5842);
  and g10424 (n5843, n_4918, n_4919);
  and g10425 (n5844, n_4688, n_4689);
  not g10426 (n_4920, n5844);
  and g10427 (n5845, n_4685, n_4920);
  and g10428 (n5846, n5843, n5845);
  not g10429 (n_4921, n5843);
  not g10430 (n_4922, n5845);
  and g10431 (n5847, n_4921, n_4922);
  not g10432 (n_4923, n5846);
  not g10433 (n_4924, n5847);
  and g10434 (n5848, n_4923, n_4924);
  and g10435 (n5849, \b[19] , n2048);
  and g10436 (n5850, \b[17] , n2198);
  and g10437 (n5851, \b[18] , n2043);
  and g10443 (n5854, n1708, n2051);
  not g10446 (n_4929, n5855);
  and g10447 (n5856, \a[23] , n_4929);
  not g10448 (n_4930, n5856);
  and g10449 (n5857, \a[23] , n_4930);
  and g10450 (n5858, n_4929, n_4930);
  not g10451 (n_4931, n5857);
  not g10452 (n_4932, n5858);
  and g10453 (n5859, n_4931, n_4932);
  not g10454 (n_4933, n5859);
  and g10455 (n5860, n5848, n_4933);
  not g10456 (n_4934, n5860);
  and g10457 (n5861, n5848, n_4934);
  and g10458 (n5862, n_4933, n_4934);
  not g10459 (n_4935, n5861);
  not g10460 (n_4936, n5862);
  and g10461 (n5863, n_4935, n_4936);
  and g10462 (n5864, n_4702, n_4707);
  and g10463 (n5865, n5863, n5864);
  not g10464 (n_4937, n5863);
  not g10465 (n_4938, n5864);
  and g10466 (n5866, n_4937, n_4938);
  not g10467 (n_4939, n5865);
  not g10468 (n_4940, n5866);
  and g10469 (n5867, n_4939, n_4940);
  and g10470 (n5868, \b[22] , n1627);
  and g10471 (n5869, \b[20] , n1763);
  and g10472 (n5870, \b[21] , n1622);
  and g10478 (n5873, n1630, n2145);
  not g10481 (n_4945, n5874);
  and g10482 (n5875, \a[20] , n_4945);
  not g10483 (n_4946, n5875);
  and g10484 (n5876, \a[20] , n_4946);
  and g10485 (n5877, n_4945, n_4946);
  not g10486 (n_4947, n5876);
  not g10487 (n_4948, n5877);
  and g10488 (n5878, n_4947, n_4948);
  not g10489 (n_4949, n5878);
  and g10490 (n5879, n5867, n_4949);
  not g10491 (n_4950, n5879);
  and g10492 (n5880, n5867, n_4950);
  and g10493 (n5881, n_4949, n_4950);
  not g10494 (n_4951, n5880);
  not g10495 (n_4952, n5881);
  and g10496 (n5882, n_4951, n_4952);
  and g10497 (n5883, n_4717, n_4723);
  and g10498 (n5884, n5882, n5883);
  not g10499 (n_4953, n5882);
  not g10500 (n_4954, n5883);
  and g10501 (n5885, n_4953, n_4954);
  not g10502 (n_4955, n5884);
  not g10503 (n_4956, n5885);
  and g10504 (n5886, n_4955, n_4956);
  and g10505 (n5887, \b[25] , n1302);
  and g10506 (n5888, \b[23] , n1391);
  and g10507 (n5889, \b[24] , n1297);
  and g10513 (n5892, n1305, n2485);
  not g10516 (n_4961, n5893);
  and g10517 (n5894, \a[17] , n_4961);
  not g10518 (n_4962, n5894);
  and g10519 (n5895, \a[17] , n_4962);
  and g10520 (n5896, n_4961, n_4962);
  not g10521 (n_4963, n5895);
  not g10522 (n_4964, n5896);
  and g10523 (n5897, n_4963, n_4964);
  not g10524 (n_4965, n5897);
  and g10525 (n5898, n5886, n_4965);
  not g10526 (n_4966, n5898);
  and g10527 (n5899, n5886, n_4966);
  and g10528 (n5900, n_4965, n_4966);
  not g10529 (n_4967, n5899);
  not g10530 (n_4968, n5900);
  and g10531 (n5901, n_4967, n_4968);
  and g10532 (n5902, n_4735, n_4738);
  not g10533 (n_4969, n5901);
  not g10534 (n_4970, n5902);
  and g10535 (n5903, n_4969, n_4970);
  and g10536 (n5904, n5901, n5902);
  not g10537 (n_4971, n5903);
  not g10538 (n_4972, n5904);
  and g10539 (n5905, n_4971, n_4972);
  not g10540 (n_4973, n5730);
  and g10541 (n5906, n_4973, n5905);
  not g10542 (n_4974, n5906);
  and g10543 (n5907, n_4973, n_4974);
  and g10544 (n5908, n5905, n_4974);
  not g10545 (n_4975, n5907);
  not g10546 (n_4976, n5908);
  and g10547 (n5909, n_4975, n_4976);
  not g10548 (n_4977, n5719);
  not g10549 (n_4978, n5909);
  and g10550 (n5910, n_4977, n_4978);
  not g10551 (n_4979, n5910);
  and g10552 (n5911, n_4977, n_4979);
  and g10553 (n5912, n_4978, n_4979);
  not g10554 (n_4980, n5911);
  not g10555 (n_4981, n5912);
  and g10556 (n5913, n_4980, n_4981);
  and g10557 (n5914, \b[31] , n700);
  and g10558 (n5915, \b[29] , n767);
  and g10559 (n5916, \b[30] , n695);
  and g10565 (n5919, n703, n3796);
  not g10568 (n_4986, n5920);
  and g10569 (n5921, \a[11] , n_4986);
  not g10570 (n_4987, n5921);
  and g10571 (n5922, \a[11] , n_4987);
  and g10572 (n5923, n_4986, n_4987);
  not g10573 (n_4988, n5922);
  not g10574 (n_4989, n5923);
  and g10575 (n5924, n_4988, n_4989);
  and g10576 (n5925, n5913, n5924);
  not g10577 (n_4990, n5913);
  not g10578 (n_4991, n5924);
  and g10579 (n5926, n_4990, n_4991);
  not g10580 (n_4992, n5925);
  not g10581 (n_4993, n5926);
  and g10582 (n5927, n_4992, n_4993);
  not g10583 (n_4994, n5717);
  and g10584 (n5928, n_4994, n5927);
  not g10585 (n_4995, n5927);
  and g10586 (n5929, n5717, n_4995);
  not g10587 (n_4996, n5928);
  not g10588 (n_4997, n5929);
  and g10589 (n5930, n_4996, n_4997);
  not g10590 (n_4998, n5930);
  and g10591 (n5931, n5716, n_4998);
  not g10592 (n_4999, n5716);
  and g10593 (n5932, n_4999, n5930);
  not g10594 (n_5000, n5931);
  not g10595 (n_5001, n5932);
  and g10596 (n5933, n_5000, n_5001);
  not g10597 (n_5002, n5705);
  and g10598 (n5934, n_5002, n5933);
  not g10599 (n_5003, n5933);
  and g10600 (n5935, n5705, n_5003);
  not g10601 (n_5004, n5934);
  not g10602 (n_5005, n5935);
  and g10603 (n5936, n_5004, n_5005);
  not g10604 (n_5006, n5703);
  and g10605 (n5937, n_5006, n5936);
  not g10606 (n_5007, n5937);
  and g10607 (n5938, n5936, n_5007);
  and g10608 (n5939, n_5006, n_5007);
  not g10609 (n_5008, n5938);
  not g10610 (n_5009, n5939);
  and g10611 (n5940, n_5008, n_5009);
  not g10612 (n_5010, n5692);
  and g10613 (n5941, n_5010, n5940);
  not g10614 (n_5011, n5940);
  and g10615 (n5942, n5692, n_5011);
  not g10616 (n_5012, n5941);
  not g10617 (n_5013, n5942);
  and g10618 (n5943, n_5012, n_5013);
  and g10619 (n5944, \b[40] , n266);
  and g10620 (n5945, \b[38] , n284);
  and g10621 (n5946, \b[39] , n261);
  and g10627 (n5949, n_4581, n_4584);
  not g10628 (n_5018, \b[40] );
  and g10629 (n5950, n_4579, n_5018);
  and g10630 (n5951, \b[39] , \b[40] );
  not g10631 (n_5019, n5950);
  not g10632 (n_5020, n5951);
  and g10633 (n5952, n_5019, n_5020);
  not g10634 (n_5021, n5949);
  and g10635 (n5953, n_5021, n5952);
  not g10636 (n_5022, n5952);
  and g10637 (n5954, n5949, n_5022);
  not g10638 (n_5023, n5953);
  not g10639 (n_5024, n5954);
  and g10640 (n5955, n_5023, n_5024);
  and g10641 (n5956, n269, n5955);
  not g10644 (n_5026, n5957);
  and g10645 (n5958, \a[2] , n_5026);
  not g10646 (n_5027, n5958);
  and g10647 (n5959, \a[2] , n_5027);
  and g10648 (n5960, n_5026, n_5027);
  not g10649 (n_5028, n5959);
  not g10650 (n_5029, n5960);
  and g10651 (n5961, n_5028, n_5029);
  not g10652 (n_5030, n5943);
  not g10653 (n_5031, n5961);
  and g10654 (n5962, n_5030, n_5031);
  and g10655 (n5963, n5943, n5961);
  not g10656 (n_5032, n5962);
  not g10657 (n_5033, n5963);
  and g10658 (n5964, n_5032, n_5033);
  not g10659 (n_5034, n5691);
  and g10660 (n5965, n_5034, n5964);
  not g10661 (n_5035, n5964);
  and g10662 (n5966, n5691, n_5035);
  not g10663 (n_5036, n5965);
  not g10664 (n_5037, n5966);
  and g10665 (\f[40] , n_5036, n_5037);
  and g10666 (n5968, n_5032, n_5036);
  and g10667 (n5969, n_5010, n_5011);
  not g10668 (n_5038, n5969);
  and g10669 (n5970, n_5007, n_5038);
  and g10670 (n5971, n_5001, n_5004);
  and g10671 (n5972, \b[35] , n511);
  and g10672 (n5973, \b[33] , n541);
  and g10673 (n5974, \b[34] , n506);
  and g10679 (n5977, n514, n4696);
  not g10682 (n_5043, n5978);
  and g10683 (n5979, \a[8] , n_5043);
  not g10684 (n_5044, n5979);
  and g10685 (n5980, \a[8] , n_5044);
  and g10686 (n5981, n_5043, n_5044);
  not g10687 (n_5045, n5980);
  not g10688 (n_5046, n5981);
  and g10689 (n5982, n_5045, n_5046);
  and g10690 (n5983, n_4993, n_4996);
  and g10691 (n5984, \b[32] , n700);
  and g10692 (n5985, \b[30] , n767);
  and g10693 (n5986, \b[31] , n695);
  and g10699 (n5989, n703, n4013);
  not g10702 (n_5051, n5990);
  and g10703 (n5991, \a[11] , n_5051);
  not g10704 (n_5052, n5991);
  and g10705 (n5992, \a[11] , n_5052);
  and g10706 (n5993, n_5051, n_5052);
  not g10707 (n_5053, n5992);
  not g10708 (n_5054, n5993);
  and g10709 (n5994, n_5053, n_5054);
  and g10710 (n5995, n_4974, n_4979);
  and g10711 (n5996, \b[29] , n951);
  and g10712 (n5997, \b[27] , n1056);
  and g10713 (n5998, \b[28] , n946);
  and g10719 (n6001, n954, n3383);
  not g10722 (n_5059, n6002);
  and g10723 (n6003, \a[14] , n_5059);
  not g10724 (n_5060, n6003);
  and g10725 (n6004, \a[14] , n_5060);
  and g10726 (n6005, n_5059, n_5060);
  not g10727 (n_5061, n6004);
  not g10728 (n_5062, n6005);
  and g10729 (n6006, n_5061, n_5062);
  and g10730 (n6007, n_4966, n_4971);
  and g10731 (n6008, n_4950, n_4956);
  and g10732 (n6009, \b[20] , n2048);
  and g10733 (n6010, \b[18] , n2198);
  and g10734 (n6011, \b[19] , n2043);
  and g10740 (n6014, n1846, n2051);
  not g10743 (n_5067, n6015);
  and g10744 (n6016, \a[23] , n_5067);
  not g10745 (n_5068, n6016);
  and g10746 (n6017, \a[23] , n_5068);
  and g10747 (n6018, n_5067, n_5068);
  not g10748 (n_5069, n6017);
  not g10749 (n_5070, n6018);
  and g10750 (n6019, n_5069, n_5070);
  and g10751 (n6020, n_4917, n_4924);
  and g10752 (n6021, \b[17] , n2539);
  and g10753 (n6022, \b[15] , n2685);
  and g10754 (n6023, \b[16] , n2534);
  and g10760 (n6026, n1356, n2542);
  not g10763 (n_5075, n6027);
  and g10764 (n6028, \a[26] , n_5075);
  not g10765 (n_5076, n6028);
  and g10766 (n6029, \a[26] , n_5076);
  and g10767 (n6030, n_5075, n_5076);
  not g10768 (n_5077, n6029);
  not g10769 (n_5078, n6030);
  and g10770 (n6031, n_5077, n_5078);
  and g10771 (n6032, n_4911, n_4914);
  and g10772 (n6033, \b[14] , n3050);
  and g10773 (n6034, \b[12] , n3243);
  and g10774 (n6035, \b[13] , n3045);
  and g10780 (n6038, n1034, n3053);
  not g10783 (n_5083, n6039);
  and g10784 (n6040, \a[29] , n_5083);
  not g10785 (n_5084, n6040);
  and g10786 (n6041, \a[29] , n_5084);
  and g10787 (n6042, n_5083, n_5084);
  not g10788 (n_5085, n6041);
  not g10789 (n_5086, n6042);
  and g10790 (n6043, n_5085, n_5086);
  and g10791 (n6044, n_4877, n_4883);
  and g10792 (n6045, \b[8] , n4287);
  and g10793 (n6046, \b[6] , n4532);
  and g10794 (n6047, \b[7] , n4282);
  and g10800 (n6050, n585, n4290);
  not g10803 (n_5091, n6051);
  and g10804 (n6052, \a[35] , n_5091);
  not g10805 (n_5092, n6052);
  and g10806 (n6053, \a[35] , n_5092);
  and g10807 (n6054, n_5091, n_5092);
  not g10808 (n_5093, n6053);
  not g10809 (n_5094, n6054);
  and g10810 (n6055, n_5093, n_5094);
  and g10811 (n6056, n_4871, n_4874);
  and g10812 (n6057, \b[2] , n5777);
  and g10813 (n6058, n5510, n_4858);
  and g10814 (n6059, n5771, n6058);
  and g10815 (n6060, \b[0] , n6059);
  and g10816 (n6061, \b[1] , n5772);
  and g10822 (n6064, n296, n5780);
  not g10825 (n_5099, n6065);
  and g10826 (n6066, \a[41] , n_5099);
  not g10827 (n_5100, n6066);
  and g10828 (n6067, \a[41] , n_5100);
  and g10829 (n6068, n_5099, n_5100);
  not g10830 (n_5101, n6067);
  not g10831 (n_5102, n6068);
  and g10832 (n6069, n_5101, n_5102);
  and g10833 (n6070, n_4866, n6069);
  not g10834 (n_5103, n6069);
  and g10835 (n6071, n5787, n_5103);
  not g10836 (n_5104, n6070);
  not g10837 (n_5105, n6071);
  and g10838 (n6072, n_5104, n_5105);
  and g10839 (n6073, \b[5] , n5035);
  and g10840 (n6074, \b[3] , n5277);
  and g10841 (n6075, \b[4] , n5030);
  and g10847 (n6078, n394, n5038);
  not g10850 (n_5110, n6079);
  and g10851 (n6080, \a[38] , n_5110);
  not g10852 (n_5111, n6080);
  and g10853 (n6081, \a[38] , n_5111);
  and g10854 (n6082, n_5110, n_5111);
  not g10855 (n_5112, n6081);
  not g10856 (n_5113, n6082);
  and g10857 (n6083, n_5112, n_5113);
  not g10858 (n_5114, n6083);
  and g10859 (n6084, n6072, n_5114);
  not g10860 (n_5115, n6084);
  and g10861 (n6085, n6072, n_5115);
  and g10862 (n6086, n_5114, n_5115);
  not g10863 (n_5116, n6085);
  not g10864 (n_5117, n6086);
  and g10865 (n6087, n_5116, n_5117);
  not g10866 (n_5118, n6056);
  not g10867 (n_5119, n6087);
  and g10868 (n6088, n_5118, n_5119);
  and g10869 (n6089, n6056, n6087);
  not g10870 (n_5120, n6088);
  not g10871 (n_5121, n6089);
  and g10872 (n6090, n_5120, n_5121);
  not g10873 (n_5122, n6055);
  and g10874 (n6091, n_5122, n6090);
  not g10875 (n_5123, n6091);
  and g10876 (n6092, n_5122, n_5123);
  and g10877 (n6093, n6090, n_5123);
  not g10878 (n_5124, n6092);
  not g10879 (n_5125, n6093);
  and g10880 (n6094, n_5124, n_5125);
  not g10881 (n_5126, n6044);
  not g10882 (n_5127, n6094);
  and g10883 (n6095, n_5126, n_5127);
  not g10884 (n_5128, n6095);
  and g10885 (n6096, n_5126, n_5128);
  and g10886 (n6097, n_5127, n_5128);
  not g10887 (n_5129, n6096);
  not g10888 (n_5130, n6097);
  and g10889 (n6098, n_5129, n_5130);
  and g10890 (n6099, \b[11] , n3638);
  and g10891 (n6100, \b[9] , n3843);
  and g10892 (n6101, \b[10] , n3633);
  and g10898 (n6104, n818, n3641);
  not g10901 (n_5135, n6105);
  and g10902 (n6106, \a[32] , n_5135);
  not g10903 (n_5136, n6106);
  and g10904 (n6107, \a[32] , n_5136);
  and g10905 (n6108, n_5135, n_5136);
  not g10906 (n_5137, n6107);
  not g10907 (n_5138, n6108);
  and g10908 (n6109, n_5137, n_5138);
  and g10909 (n6110, n6098, n6109);
  not g10910 (n_5139, n6098);
  not g10911 (n_5140, n6109);
  and g10912 (n6111, n_5139, n_5140);
  not g10913 (n_5141, n6110);
  not g10914 (n_5142, n6111);
  and g10915 (n6112, n_5141, n_5142);
  not g10916 (n_5143, n5820);
  and g10917 (n6113, n_5143, n6112);
  not g10918 (n_5144, n6112);
  and g10919 (n6114, n5820, n_5144);
  not g10920 (n_5145, n6113);
  not g10921 (n_5146, n6114);
  and g10922 (n6115, n_5145, n_5146);
  not g10923 (n_5147, n6115);
  and g10924 (n6116, n6043, n_5147);
  not g10925 (n_5148, n6043);
  and g10926 (n6117, n_5148, n6115);
  not g10927 (n_5149, n6116);
  not g10928 (n_5150, n6117);
  and g10929 (n6118, n_5149, n_5150);
  not g10930 (n_5151, n6032);
  and g10931 (n6119, n_5151, n6118);
  not g10932 (n_5152, n6118);
  and g10933 (n6120, n6032, n_5152);
  not g10934 (n_5153, n6119);
  not g10935 (n_5154, n6120);
  and g10936 (n6121, n_5153, n_5154);
  not g10937 (n_5155, n6121);
  and g10938 (n6122, n6031, n_5155);
  not g10939 (n_5156, n6031);
  and g10940 (n6123, n_5156, n6121);
  not g10941 (n_5157, n6122);
  not g10942 (n_5158, n6123);
  and g10943 (n6124, n_5157, n_5158);
  not g10944 (n_5159, n6020);
  and g10945 (n6125, n_5159, n6124);
  not g10946 (n_5160, n6124);
  and g10947 (n6126, n6020, n_5160);
  not g10948 (n_5161, n6125);
  not g10949 (n_5162, n6126);
  and g10950 (n6127, n_5161, n_5162);
  not g10951 (n_5163, n6019);
  and g10952 (n6128, n_5163, n6127);
  not g10953 (n_5164, n6128);
  and g10954 (n6129, n6127, n_5164);
  and g10955 (n6130, n_5163, n_5164);
  not g10956 (n_5165, n6129);
  not g10957 (n_5166, n6130);
  and g10958 (n6131, n_5165, n_5166);
  and g10959 (n6132, n_4934, n_4940);
  and g10960 (n6133, n6131, n6132);
  not g10961 (n_5167, n6131);
  not g10962 (n_5168, n6132);
  and g10963 (n6134, n_5167, n_5168);
  not g10964 (n_5169, n6133);
  not g10965 (n_5170, n6134);
  and g10966 (n6135, n_5169, n_5170);
  and g10967 (n6136, \b[23] , n1627);
  and g10968 (n6137, \b[21] , n1763);
  and g10969 (n6138, \b[22] , n1622);
  and g10975 (n6141, n1630, n2300);
  not g10978 (n_5175, n6142);
  and g10979 (n6143, \a[20] , n_5175);
  not g10980 (n_5176, n6143);
  and g10981 (n6144, \a[20] , n_5176);
  and g10982 (n6145, n_5175, n_5176);
  not g10983 (n_5177, n6144);
  not g10984 (n_5178, n6145);
  and g10985 (n6146, n_5177, n_5178);
  not g10986 (n_5179, n6146);
  and g10987 (n6147, n6135, n_5179);
  not g10988 (n_5180, n6135);
  and g10989 (n6148, n_5180, n6146);
  not g10990 (n_5181, n6008);
  not g10991 (n_5182, n6148);
  and g10992 (n6149, n_5181, n_5182);
  not g10993 (n_5183, n6147);
  and g10994 (n6150, n_5183, n6149);
  not g10995 (n_5184, n6150);
  and g10996 (n6151, n_5181, n_5184);
  and g10997 (n6152, n_5183, n_5184);
  and g10998 (n6153, n_5182, n6152);
  not g10999 (n_5185, n6151);
  not g11000 (n_5186, n6153);
  and g11001 (n6154, n_5185, n_5186);
  and g11002 (n6155, \b[26] , n1302);
  and g11003 (n6156, \b[24] , n1391);
  and g11004 (n6157, \b[25] , n1297);
  and g11010 (n6160, n1305, n2813);
  not g11013 (n_5191, n6161);
  and g11014 (n6162, \a[17] , n_5191);
  not g11015 (n_5192, n6162);
  and g11016 (n6163, \a[17] , n_5192);
  and g11017 (n6164, n_5191, n_5192);
  not g11018 (n_5193, n6163);
  not g11019 (n_5194, n6164);
  and g11020 (n6165, n_5193, n_5194);
  and g11021 (n6166, n6154, n6165);
  not g11022 (n_5195, n6154);
  not g11023 (n_5196, n6165);
  and g11024 (n6167, n_5195, n_5196);
  not g11025 (n_5197, n6166);
  not g11026 (n_5198, n6167);
  and g11027 (n6168, n_5197, n_5198);
  not g11028 (n_5199, n6007);
  and g11029 (n6169, n_5199, n6168);
  not g11030 (n_5200, n6168);
  and g11031 (n6170, n6007, n_5200);
  not g11032 (n_5201, n6169);
  not g11033 (n_5202, n6170);
  and g11034 (n6171, n_5201, n_5202);
  not g11035 (n_5203, n6171);
  and g11036 (n6172, n6006, n_5203);
  not g11037 (n_5204, n6006);
  and g11038 (n6173, n_5204, n6171);
  not g11039 (n_5205, n6172);
  not g11040 (n_5206, n6173);
  and g11041 (n6174, n_5205, n_5206);
  not g11042 (n_5207, n5995);
  and g11043 (n6175, n_5207, n6174);
  not g11044 (n_5208, n6174);
  and g11045 (n6176, n5995, n_5208);
  not g11046 (n_5209, n6175);
  not g11047 (n_5210, n6176);
  and g11048 (n6177, n_5209, n_5210);
  not g11049 (n_5211, n6177);
  and g11050 (n6178, n5994, n_5211);
  not g11051 (n_5212, n5994);
  and g11052 (n6179, n_5212, n6177);
  not g11053 (n_5213, n6178);
  not g11054 (n_5214, n6179);
  and g11055 (n6180, n_5213, n_5214);
  not g11056 (n_5215, n5983);
  and g11057 (n6181, n_5215, n6180);
  not g11058 (n_5216, n6180);
  and g11059 (n6182, n5983, n_5216);
  not g11060 (n_5217, n6181);
  not g11061 (n_5218, n6182);
  and g11062 (n6183, n_5217, n_5218);
  not g11063 (n_5219, n5982);
  and g11064 (n6184, n_5219, n6183);
  not g11065 (n_5220, n6184);
  and g11066 (n6185, n6183, n_5220);
  and g11067 (n6186, n_5219, n_5220);
  not g11068 (n_5221, n6185);
  not g11069 (n_5222, n6186);
  and g11070 (n6187, n_5221, n_5222);
  not g11071 (n_5223, n5971);
  and g11072 (n6188, n_5223, n6187);
  not g11073 (n_5224, n6187);
  and g11074 (n6189, n5971, n_5224);
  not g11075 (n_5225, n6188);
  not g11076 (n_5226, n6189);
  and g11077 (n6190, n_5225, n_5226);
  and g11078 (n6191, \b[38] , n362);
  and g11079 (n6192, \b[36] , n403);
  and g11080 (n6193, \b[37] , n357);
  and g11086 (n6196, n365, n5205);
  not g11089 (n_5231, n6197);
  and g11090 (n6198, \a[5] , n_5231);
  not g11091 (n_5232, n6198);
  and g11092 (n6199, \a[5] , n_5232);
  and g11093 (n6200, n_5231, n_5232);
  not g11094 (n_5233, n6199);
  not g11095 (n_5234, n6200);
  and g11096 (n6201, n_5233, n_5234);
  not g11097 (n_5235, n6190);
  not g11098 (n_5236, n6201);
  and g11099 (n6202, n_5235, n_5236);
  and g11100 (n6203, n6190, n6201);
  not g11101 (n_5237, n6202);
  not g11102 (n_5238, n6203);
  and g11103 (n6204, n_5237, n_5238);
  not g11104 (n_5239, n6204);
  and g11105 (n6205, n5970, n_5239);
  not g11106 (n_5240, n5970);
  and g11107 (n6206, n_5240, n6204);
  not g11108 (n_5241, n6205);
  not g11109 (n_5242, n6206);
  and g11110 (n6207, n_5241, n_5242);
  and g11111 (n6208, \b[41] , n266);
  and g11112 (n6209, \b[39] , n284);
  and g11113 (n6210, \b[40] , n261);
  and g11119 (n6213, n_5020, n_5023);
  not g11120 (n_5247, \b[41] );
  and g11121 (n6214, n_5018, n_5247);
  and g11122 (n6215, \b[40] , \b[41] );
  not g11123 (n_5248, n6214);
  not g11124 (n_5249, n6215);
  and g11125 (n6216, n_5248, n_5249);
  not g11126 (n_5250, n6213);
  and g11127 (n6217, n_5250, n6216);
  not g11128 (n_5251, n6216);
  and g11129 (n6218, n6213, n_5251);
  not g11130 (n_5252, n6217);
  not g11131 (n_5253, n6218);
  and g11132 (n6219, n_5252, n_5253);
  and g11133 (n6220, n269, n6219);
  not g11136 (n_5255, n6221);
  and g11137 (n6222, \a[2] , n_5255);
  not g11138 (n_5256, n6222);
  and g11139 (n6223, \a[2] , n_5256);
  and g11140 (n6224, n_5255, n_5256);
  not g11141 (n_5257, n6223);
  not g11142 (n_5258, n6224);
  and g11143 (n6225, n_5257, n_5258);
  not g11144 (n_5259, n6207);
  and g11145 (n6226, n_5259, n6225);
  not g11146 (n_5260, n6225);
  and g11147 (n6227, n6207, n_5260);
  not g11148 (n_5261, n6226);
  not g11149 (n_5262, n6227);
  and g11150 (n6228, n_5261, n_5262);
  not g11151 (n_5263, n5968);
  and g11152 (n6229, n_5263, n6228);
  not g11153 (n_5264, n6228);
  and g11154 (n6230, n5968, n_5264);
  not g11155 (n_5265, n6229);
  not g11156 (n_5266, n6230);
  and g11157 (\f[41] , n_5265, n_5266);
  and g11158 (n6232, n_5237, n_5242);
  and g11159 (n6233, \b[39] , n362);
  and g11160 (n6234, \b[37] , n403);
  and g11161 (n6235, \b[38] , n357);
  and g11167 (n6238, n365, n5451);
  not g11170 (n_5271, n6239);
  and g11171 (n6240, \a[5] , n_5271);
  not g11172 (n_5272, n6240);
  and g11173 (n6241, \a[5] , n_5272);
  and g11174 (n6242, n_5271, n_5272);
  not g11175 (n_5273, n6241);
  not g11176 (n_5274, n6242);
  and g11177 (n6243, n_5273, n_5274);
  and g11178 (n6244, n_5223, n_5224);
  not g11179 (n_5275, n6244);
  and g11180 (n6245, n_5220, n_5275);
  and g11181 (n6246, n_5214, n_5217);
  and g11182 (n6247, \b[33] , n700);
  and g11183 (n6248, \b[31] , n767);
  and g11184 (n6249, \b[32] , n695);
  and g11190 (n6252, n703, n4223);
  not g11193 (n_5280, n6253);
  and g11194 (n6254, \a[11] , n_5280);
  not g11195 (n_5281, n6254);
  and g11196 (n6255, \a[11] , n_5281);
  and g11197 (n6256, n_5280, n_5281);
  not g11198 (n_5282, n6255);
  not g11199 (n_5283, n6256);
  and g11200 (n6257, n_5282, n_5283);
  and g11201 (n6258, n_5206, n_5209);
  and g11202 (n6259, n_5198, n_5201);
  and g11203 (n6260, \b[27] , n1302);
  and g11204 (n6261, \b[25] , n1391);
  and g11205 (n6262, \b[26] , n1297);
  and g11211 (n6265, n1305, n2990);
  not g11214 (n_5288, n6266);
  and g11215 (n6267, \a[17] , n_5288);
  not g11216 (n_5289, n6267);
  and g11217 (n6268, \a[17] , n_5289);
  and g11218 (n6269, n_5288, n_5289);
  not g11219 (n_5290, n6268);
  not g11220 (n_5291, n6269);
  and g11221 (n6270, n_5290, n_5291);
  and g11222 (n6271, \b[21] , n2048);
  and g11223 (n6272, \b[19] , n2198);
  and g11224 (n6273, \b[20] , n2043);
  and g11230 (n6276, n1984, n2051);
  not g11233 (n_5296, n6277);
  and g11234 (n6278, \a[23] , n_5296);
  not g11235 (n_5297, n6278);
  and g11236 (n6279, \a[23] , n_5297);
  and g11237 (n6280, n_5296, n_5297);
  not g11238 (n_5298, n6279);
  not g11239 (n_5299, n6280);
  and g11240 (n6281, n_5298, n_5299);
  and g11241 (n6282, n_5158, n_5161);
  and g11242 (n6283, n_5150, n_5153);
  and g11243 (n6284, n_5142, n_5145);
  and g11244 (n6285, \b[12] , n3638);
  and g11245 (n6286, \b[10] , n3843);
  and g11246 (n6287, \b[11] , n3633);
  and g11252 (n6290, n842, n3641);
  not g11255 (n_5304, n6291);
  and g11256 (n6292, \a[32] , n_5304);
  not g11257 (n_5305, n6292);
  and g11258 (n6293, \a[32] , n_5305);
  and g11259 (n6294, n_5304, n_5305);
  not g11260 (n_5306, n6293);
  not g11261 (n_5307, n6294);
  and g11262 (n6295, n_5306, n_5307);
  and g11263 (n6296, n_5123, n_5128);
  and g11264 (n6297, \b[6] , n5035);
  and g11265 (n6298, \b[4] , n5277);
  and g11266 (n6299, \b[5] , n5030);
  and g11272 (n6302, n459, n5038);
  not g11275 (n_5312, n6303);
  and g11276 (n6304, \a[38] , n_5312);
  not g11277 (n_5313, n6304);
  and g11278 (n6305, \a[38] , n_5313);
  and g11279 (n6306, n_5312, n_5313);
  not g11280 (n_5314, n6305);
  not g11281 (n_5315, n6306);
  and g11282 (n6307, n_5314, n_5315);
  not g11283 (n_5317, \a[42] );
  and g11284 (n6308, \a[41] , n_5317);
  and g11285 (n6309, n_4853, \a[42] );
  not g11286 (n_5318, n6308);
  not g11287 (n_5319, n6309);
  and g11288 (n6310, n_5318, n_5319);
  not g11289 (n_5320, n6310);
  and g11290 (n6311, \b[0] , n_5320);
  and g11291 (n6312, n_5105, n6311);
  not g11292 (n_5321, n6311);
  and g11293 (n6313, n6071, n_5321);
  not g11294 (n_5322, n6312);
  not g11295 (n_5323, n6313);
  and g11296 (n6314, n_5322, n_5323);
  and g11297 (n6315, \b[3] , n5777);
  and g11298 (n6316, \b[1] , n6059);
  and g11299 (n6317, \b[2] , n5772);
  and g11305 (n6320, n318, n5780);
  not g11308 (n_5328, n6321);
  and g11309 (n6322, \a[41] , n_5328);
  not g11310 (n_5329, n6322);
  and g11311 (n6323, \a[41] , n_5329);
  and g11312 (n6324, n_5328, n_5329);
  not g11313 (n_5330, n6323);
  not g11314 (n_5331, n6324);
  and g11315 (n6325, n_5330, n_5331);
  not g11316 (n_5332, n6314);
  not g11317 (n_5333, n6325);
  and g11318 (n6326, n_5332, n_5333);
  and g11319 (n6327, n6314, n6325);
  not g11320 (n_5334, n6326);
  not g11321 (n_5335, n6327);
  and g11322 (n6328, n_5334, n_5335);
  not g11323 (n_5336, n6307);
  and g11324 (n6329, n_5336, n6328);
  not g11325 (n_5337, n6329);
  and g11326 (n6330, n6328, n_5337);
  and g11327 (n6331, n_5336, n_5337);
  not g11328 (n_5338, n6330);
  not g11329 (n_5339, n6331);
  and g11330 (n6332, n_5338, n_5339);
  and g11331 (n6333, n_5115, n_5120);
  and g11332 (n6334, n6332, n6333);
  not g11333 (n_5340, n6332);
  not g11334 (n_5341, n6333);
  and g11335 (n6335, n_5340, n_5341);
  not g11336 (n_5342, n6334);
  not g11337 (n_5343, n6335);
  and g11338 (n6336, n_5342, n_5343);
  and g11339 (n6337, \b[9] , n4287);
  and g11340 (n6338, \b[7] , n4532);
  and g11341 (n6339, \b[8] , n4282);
  and g11347 (n6342, n651, n4290);
  not g11350 (n_5348, n6343);
  and g11351 (n6344, \a[35] , n_5348);
  not g11352 (n_5349, n6344);
  and g11353 (n6345, \a[35] , n_5349);
  and g11354 (n6346, n_5348, n_5349);
  not g11355 (n_5350, n6345);
  not g11356 (n_5351, n6346);
  and g11357 (n6347, n_5350, n_5351);
  not g11358 (n_5352, n6336);
  and g11359 (n6348, n_5352, n6347);
  not g11360 (n_5353, n6347);
  and g11361 (n6349, n6336, n_5353);
  not g11362 (n_5354, n6348);
  not g11363 (n_5355, n6349);
  and g11364 (n6350, n_5354, n_5355);
  not g11365 (n_5356, n6296);
  and g11366 (n6351, n_5356, n6350);
  not g11367 (n_5357, n6350);
  and g11368 (n6352, n6296, n_5357);
  not g11369 (n_5358, n6351);
  not g11370 (n_5359, n6352);
  and g11371 (n6353, n_5358, n_5359);
  not g11372 (n_5360, n6295);
  and g11373 (n6354, n_5360, n6353);
  not g11374 (n_5361, n6354);
  and g11375 (n6355, n_5360, n_5361);
  and g11376 (n6356, n6353, n_5361);
  not g11377 (n_5362, n6355);
  not g11378 (n_5363, n6356);
  and g11379 (n6357, n_5362, n_5363);
  not g11380 (n_5364, n6284);
  not g11381 (n_5365, n6357);
  and g11382 (n6358, n_5364, n_5365);
  not g11383 (n_5366, n6358);
  and g11384 (n6359, n_5364, n_5366);
  and g11385 (n6360, n_5365, n_5366);
  not g11386 (n_5367, n6359);
  not g11387 (n_5368, n6360);
  and g11388 (n6361, n_5367, n_5368);
  and g11389 (n6362, \b[15] , n3050);
  and g11390 (n6363, \b[13] , n3243);
  and g11391 (n6364, \b[14] , n3045);
  and g11397 (n6367, n1131, n3053);
  not g11400 (n_5373, n6368);
  and g11401 (n6369, \a[29] , n_5373);
  not g11402 (n_5374, n6369);
  and g11403 (n6370, \a[29] , n_5374);
  and g11404 (n6371, n_5373, n_5374);
  not g11405 (n_5375, n6370);
  not g11406 (n_5376, n6371);
  and g11407 (n6372, n_5375, n_5376);
  not g11408 (n_5377, n6361);
  not g11409 (n_5378, n6372);
  and g11410 (n6373, n_5377, n_5378);
  not g11411 (n_5379, n6373);
  and g11412 (n6374, n_5377, n_5379);
  and g11413 (n6375, n_5378, n_5379);
  not g11414 (n_5380, n6374);
  not g11415 (n_5381, n6375);
  and g11416 (n6376, n_5380, n_5381);
  not g11417 (n_5382, n6283);
  and g11418 (n6377, n_5382, n6376);
  not g11419 (n_5383, n6376);
  and g11420 (n6378, n6283, n_5383);
  not g11421 (n_5384, n6377);
  not g11422 (n_5385, n6378);
  and g11423 (n6379, n_5384, n_5385);
  and g11424 (n6380, \b[18] , n2539);
  and g11425 (n6381, \b[16] , n2685);
  and g11426 (n6382, \b[17] , n2534);
  and g11432 (n6385, n1566, n2542);
  not g11435 (n_5390, n6386);
  and g11436 (n6387, \a[26] , n_5390);
  not g11437 (n_5391, n6387);
  and g11438 (n6388, \a[26] , n_5391);
  and g11439 (n6389, n_5390, n_5391);
  not g11440 (n_5392, n6388);
  not g11441 (n_5393, n6389);
  and g11442 (n6390, n_5392, n_5393);
  not g11443 (n_5394, n6379);
  not g11444 (n_5395, n6390);
  and g11445 (n6391, n_5394, n_5395);
  and g11446 (n6392, n6379, n6390);
  not g11447 (n_5396, n6391);
  not g11448 (n_5397, n6392);
  and g11449 (n6393, n_5396, n_5397);
  not g11450 (n_5398, n6282);
  and g11451 (n6394, n_5398, n6393);
  not g11452 (n_5399, n6393);
  and g11453 (n6395, n6282, n_5399);
  not g11454 (n_5400, n6394);
  not g11455 (n_5401, n6395);
  and g11456 (n6396, n_5400, n_5401);
  not g11457 (n_5402, n6281);
  and g11458 (n6397, n_5402, n6396);
  not g11459 (n_5403, n6397);
  and g11460 (n6398, n6396, n_5403);
  and g11461 (n6399, n_5402, n_5403);
  not g11462 (n_5404, n6398);
  not g11463 (n_5405, n6399);
  and g11464 (n6400, n_5404, n_5405);
  and g11465 (n6401, n_5164, n_5170);
  and g11466 (n6402, n6400, n6401);
  not g11467 (n_5406, n6400);
  not g11468 (n_5407, n6401);
  and g11469 (n6403, n_5406, n_5407);
  not g11470 (n_5408, n6402);
  not g11471 (n_5409, n6403);
  and g11472 (n6404, n_5408, n_5409);
  and g11473 (n6405, \b[24] , n1627);
  and g11474 (n6406, \b[22] , n1763);
  and g11475 (n6407, \b[23] , n1622);
  and g11481 (n6410, n1630, n2458);
  not g11484 (n_5414, n6411);
  and g11485 (n6412, \a[20] , n_5414);
  not g11486 (n_5415, n6412);
  and g11487 (n6413, \a[20] , n_5415);
  and g11488 (n6414, n_5414, n_5415);
  not g11489 (n_5416, n6413);
  not g11490 (n_5417, n6414);
  and g11491 (n6415, n_5416, n_5417);
  not g11492 (n_5418, n6404);
  and g11493 (n6416, n_5418, n6415);
  not g11494 (n_5419, n6415);
  and g11495 (n6417, n6404, n_5419);
  not g11496 (n_5420, n6416);
  not g11497 (n_5421, n6417);
  and g11498 (n6418, n_5420, n_5421);
  not g11499 (n_5422, n6152);
  and g11500 (n6419, n_5422, n6418);
  not g11501 (n_5423, n6418);
  and g11502 (n6420, n6152, n_5423);
  not g11503 (n_5424, n6419);
  not g11504 (n_5425, n6420);
  and g11505 (n6421, n_5424, n_5425);
  not g11506 (n_5426, n6270);
  and g11507 (n6422, n_5426, n6421);
  not g11508 (n_5427, n6422);
  and g11509 (n6423, n6421, n_5427);
  and g11510 (n6424, n_5426, n_5427);
  not g11511 (n_5428, n6423);
  not g11512 (n_5429, n6424);
  and g11513 (n6425, n_5428, n_5429);
  not g11514 (n_5430, n6259);
  and g11515 (n6426, n_5430, n6425);
  not g11516 (n_5431, n6425);
  and g11517 (n6427, n6259, n_5431);
  not g11518 (n_5432, n6426);
  not g11519 (n_5433, n6427);
  and g11520 (n6428, n_5432, n_5433);
  and g11521 (n6429, \b[30] , n951);
  and g11522 (n6430, \b[28] , n1056);
  and g11523 (n6431, \b[29] , n946);
  and g11529 (n6434, n954, n3577);
  not g11532 (n_5438, n6435);
  and g11533 (n6436, \a[14] , n_5438);
  not g11534 (n_5439, n6436);
  and g11535 (n6437, \a[14] , n_5439);
  and g11536 (n6438, n_5438, n_5439);
  not g11537 (n_5440, n6437);
  not g11538 (n_5441, n6438);
  and g11539 (n6439, n_5440, n_5441);
  not g11540 (n_5442, n6428);
  not g11541 (n_5443, n6439);
  and g11542 (n6440, n_5442, n_5443);
  and g11543 (n6441, n6428, n6439);
  not g11544 (n_5444, n6440);
  not g11545 (n_5445, n6441);
  and g11546 (n6442, n_5444, n_5445);
  not g11547 (n_5446, n6258);
  and g11548 (n6443, n_5446, n6442);
  not g11549 (n_5447, n6442);
  and g11550 (n6444, n6258, n_5447);
  not g11551 (n_5448, n6443);
  not g11552 (n_5449, n6444);
  and g11553 (n6445, n_5448, n_5449);
  not g11554 (n_5450, n6257);
  and g11555 (n6446, n_5450, n6445);
  not g11556 (n_5451, n6446);
  and g11557 (n6447, n6445, n_5451);
  and g11558 (n6448, n_5450, n_5451);
  not g11559 (n_5452, n6447);
  not g11560 (n_5453, n6448);
  and g11561 (n6449, n_5452, n_5453);
  not g11562 (n_5454, n6246);
  and g11563 (n6450, n_5454, n6449);
  not g11564 (n_5455, n6449);
  and g11565 (n6451, n6246, n_5455);
  not g11566 (n_5456, n6450);
  not g11567 (n_5457, n6451);
  and g11568 (n6452, n_5456, n_5457);
  and g11569 (n6453, \b[36] , n511);
  and g11570 (n6454, \b[34] , n541);
  and g11571 (n6455, \b[35] , n506);
  and g11577 (n6458, n514, n4922);
  not g11580 (n_5462, n6459);
  and g11581 (n6460, \a[8] , n_5462);
  not g11582 (n_5463, n6460);
  and g11583 (n6461, \a[8] , n_5463);
  and g11584 (n6462, n_5462, n_5463);
  not g11585 (n_5464, n6461);
  not g11586 (n_5465, n6462);
  and g11587 (n6463, n_5464, n_5465);
  and g11588 (n6464, n6452, n6463);
  not g11589 (n_5466, n6452);
  not g11590 (n_5467, n6463);
  and g11591 (n6465, n_5466, n_5467);
  not g11592 (n_5468, n6464);
  not g11593 (n_5469, n6465);
  and g11594 (n6466, n_5468, n_5469);
  not g11595 (n_5470, n6245);
  and g11596 (n6467, n_5470, n6466);
  not g11597 (n_5471, n6466);
  and g11598 (n6468, n6245, n_5471);
  not g11599 (n_5472, n6467);
  not g11600 (n_5473, n6468);
  and g11601 (n6469, n_5472, n_5473);
  not g11602 (n_5474, n6243);
  and g11603 (n6470, n_5474, n6469);
  not g11604 (n_5475, n6470);
  and g11605 (n6471, n_5474, n_5475);
  and g11606 (n6472, n6469, n_5475);
  not g11607 (n_5476, n6471);
  not g11608 (n_5477, n6472);
  and g11609 (n6473, n_5476, n_5477);
  not g11610 (n_5478, n6232);
  not g11611 (n_5479, n6473);
  and g11612 (n6474, n_5478, n_5479);
  not g11613 (n_5480, n6474);
  and g11614 (n6475, n_5478, n_5480);
  and g11615 (n6476, n_5479, n_5480);
  not g11616 (n_5481, n6475);
  not g11617 (n_5482, n6476);
  and g11618 (n6477, n_5481, n_5482);
  and g11619 (n6478, \b[42] , n266);
  and g11620 (n6479, \b[40] , n284);
  and g11621 (n6480, \b[41] , n261);
  and g11627 (n6483, n_5249, n_5252);
  not g11628 (n_5487, \b[42] );
  and g11629 (n6484, n_5247, n_5487);
  and g11630 (n6485, \b[41] , \b[42] );
  not g11631 (n_5488, n6484);
  not g11632 (n_5489, n6485);
  and g11633 (n6486, n_5488, n_5489);
  not g11634 (n_5490, n6483);
  and g11635 (n6487, n_5490, n6486);
  not g11636 (n_5491, n6486);
  and g11637 (n6488, n6483, n_5491);
  not g11638 (n_5492, n6487);
  not g11639 (n_5493, n6488);
  and g11640 (n6489, n_5492, n_5493);
  and g11641 (n6490, n269, n6489);
  not g11644 (n_5495, n6491);
  and g11645 (n6492, \a[2] , n_5495);
  not g11646 (n_5496, n6492);
  and g11647 (n6493, \a[2] , n_5496);
  and g11648 (n6494, n_5495, n_5496);
  not g11649 (n_5497, n6493);
  not g11650 (n_5498, n6494);
  and g11651 (n6495, n_5497, n_5498);
  not g11652 (n_5499, n6477);
  not g11653 (n_5500, n6495);
  and g11654 (n6496, n_5499, n_5500);
  not g11655 (n_5501, n6496);
  and g11656 (n6497, n_5499, n_5501);
  and g11657 (n6498, n_5500, n_5501);
  not g11658 (n_5502, n6497);
  not g11659 (n_5503, n6498);
  and g11660 (n6499, n_5502, n_5503);
  and g11661 (n6500, n_5262, n_5265);
  not g11662 (n_5504, n6499);
  not g11663 (n_5505, n6500);
  and g11664 (n6501, n_5504, n_5505);
  and g11665 (n6502, n6499, n6500);
  not g11666 (n_5506, n6501);
  not g11667 (n_5507, n6502);
  and g11668 (\f[42] , n_5506, n_5507);
  and g11669 (n6504, \b[43] , n266);
  and g11670 (n6505, \b[41] , n284);
  and g11671 (n6506, \b[42] , n261);
  and g11677 (n6509, n_5489, n_5492);
  not g11678 (n_5512, \b[43] );
  and g11679 (n6510, n_5487, n_5512);
  and g11680 (n6511, \b[42] , \b[43] );
  not g11681 (n_5513, n6510);
  not g11682 (n_5514, n6511);
  and g11683 (n6512, n_5513, n_5514);
  not g11684 (n_5515, n6509);
  and g11685 (n6513, n_5515, n6512);
  not g11686 (n_5516, n6512);
  and g11687 (n6514, n6509, n_5516);
  not g11688 (n_5517, n6513);
  not g11689 (n_5518, n6514);
  and g11690 (n6515, n_5517, n_5518);
  and g11691 (n6516, n269, n6515);
  not g11694 (n_5520, n6517);
  and g11695 (n6518, \a[2] , n_5520);
  not g11696 (n_5521, n6518);
  and g11697 (n6519, \a[2] , n_5521);
  and g11698 (n6520, n_5520, n_5521);
  not g11699 (n_5522, n6519);
  not g11700 (n_5523, n6520);
  and g11701 (n6521, n_5522, n_5523);
  and g11702 (n6522, n_5475, n_5480);
  and g11703 (n6523, n_5469, n_5472);
  and g11704 (n6524, \b[34] , n700);
  and g11705 (n6525, \b[32] , n767);
  and g11706 (n6526, \b[33] , n695);
  and g11712 (n6529, n703, n4466);
  not g11715 (n_5528, n6530);
  and g11716 (n6531, \a[11] , n_5528);
  not g11717 (n_5529, n6531);
  and g11718 (n6532, \a[11] , n_5529);
  and g11719 (n6533, n_5528, n_5529);
  not g11720 (n_5530, n6532);
  not g11721 (n_5531, n6533);
  and g11722 (n6534, n_5530, n_5531);
  and g11723 (n6535, n_5444, n_5448);
  and g11724 (n6536, n_5430, n_5431);
  not g11725 (n_5532, n6536);
  and g11726 (n6537, n_5427, n_5532);
  and g11727 (n6538, \b[28] , n1302);
  and g11728 (n6539, \b[26] , n1391);
  and g11729 (n6540, \b[27] , n1297);
  and g11735 (n6543, n1305, n3189);
  not g11738 (n_5537, n6544);
  and g11739 (n6545, \a[17] , n_5537);
  not g11740 (n_5538, n6545);
  and g11741 (n6546, \a[17] , n_5538);
  and g11742 (n6547, n_5537, n_5538);
  not g11743 (n_5539, n6546);
  not g11744 (n_5540, n6547);
  and g11745 (n6548, n_5539, n_5540);
  and g11746 (n6549, \b[16] , n3050);
  and g11747 (n6550, \b[14] , n3243);
  and g11748 (n6551, \b[15] , n3045);
  and g11754 (n6554, n1237, n3053);
  not g11757 (n_5545, n6555);
  and g11758 (n6556, \a[29] , n_5545);
  not g11759 (n_5546, n6556);
  and g11760 (n6557, \a[29] , n_5546);
  and g11761 (n6558, n_5545, n_5546);
  not g11762 (n_5547, n6557);
  not g11763 (n_5548, n6558);
  and g11764 (n6559, n_5547, n_5548);
  and g11765 (n6560, n_5361, n_5366);
  and g11766 (n6561, n_5355, n_5358);
  and g11767 (n6562, \b[7] , n5035);
  and g11768 (n6563, \b[5] , n5277);
  and g11769 (n6564, \b[6] , n5030);
  and g11775 (n6567, n484, n5038);
  not g11778 (n_5553, n6568);
  and g11779 (n6569, \a[38] , n_5553);
  not g11780 (n_5554, n6569);
  and g11781 (n6570, \a[38] , n_5554);
  and g11782 (n6571, n_5553, n_5554);
  not g11783 (n_5555, n6570);
  not g11784 (n_5556, n6571);
  and g11785 (n6572, n_5555, n_5556);
  and g11786 (n6573, n6071, n6311);
  not g11787 (n_5557, n6573);
  and g11788 (n6574, n_5334, n_5557);
  and g11789 (n6575, \b[4] , n5777);
  and g11790 (n6576, \b[2] , n6059);
  and g11791 (n6577, \b[3] , n5772);
  and g11797 (n6580, n346, n5780);
  not g11800 (n_5562, n6581);
  and g11801 (n6582, \a[41] , n_5562);
  not g11802 (n_5563, n6582);
  and g11803 (n6583, \a[41] , n_5563);
  and g11804 (n6584, n_5562, n_5563);
  not g11805 (n_5564, n6583);
  not g11806 (n_5565, n6584);
  and g11807 (n6585, n_5564, n_5565);
  and g11808 (n6586, \a[44] , n_5321);
  and g11809 (n6587, n_5317, \a[43] );
  not g11810 (n_5568, \a[43] );
  and g11811 (n6588, \a[42] , n_5568);
  not g11812 (n_5569, n6587);
  not g11813 (n_5570, n6588);
  and g11814 (n6589, n_5569, n_5570);
  not g11815 (n_5571, n6589);
  and g11816 (n6590, n6310, n_5571);
  and g11817 (n6591, \b[0] , n6590);
  and g11818 (n6592, n_5568, \a[44] );
  not g11819 (n_5572, \a[44] );
  and g11820 (n6593, \a[43] , n_5572);
  not g11821 (n_5573, n6592);
  not g11822 (n_5574, n6593);
  and g11823 (n6594, n_5573, n_5574);
  and g11824 (n6595, n_5320, n6594);
  and g11825 (n6596, \b[1] , n6595);
  not g11826 (n_5575, n6591);
  not g11827 (n_5576, n6596);
  and g11828 (n6597, n_5575, n_5576);
  not g11829 (n_5577, n6594);
  and g11830 (n6598, n_5320, n_5577);
  and g11831 (n6599, n_21, n6598);
  not g11832 (n_5578, n6599);
  and g11833 (n6600, n6597, n_5578);
  not g11834 (n_5579, n6600);
  and g11835 (n6601, \a[44] , n_5579);
  not g11836 (n_5580, n6601);
  and g11837 (n6602, \a[44] , n_5580);
  and g11838 (n6603, n_5579, n_5580);
  not g11839 (n_5581, n6602);
  not g11840 (n_5582, n6603);
  and g11841 (n6604, n_5581, n_5582);
  not g11842 (n_5583, n6604);
  and g11843 (n6605, n6586, n_5583);
  not g11844 (n_5584, n6586);
  and g11845 (n6606, n_5584, n6604);
  not g11846 (n_5585, n6605);
  not g11847 (n_5586, n6606);
  and g11848 (n6607, n_5585, n_5586);
  not g11849 (n_5587, n6607);
  and g11850 (n6608, n6585, n_5587);
  not g11851 (n_5588, n6585);
  and g11852 (n6609, n_5588, n6607);
  not g11853 (n_5589, n6608);
  not g11854 (n_5590, n6609);
  and g11855 (n6610, n_5589, n_5590);
  not g11856 (n_5591, n6574);
  and g11857 (n6611, n_5591, n6610);
  not g11858 (n_5592, n6610);
  and g11859 (n6612, n6574, n_5592);
  not g11860 (n_5593, n6611);
  not g11861 (n_5594, n6612);
  and g11862 (n6613, n_5593, n_5594);
  not g11863 (n_5595, n6572);
  and g11864 (n6614, n_5595, n6613);
  not g11865 (n_5596, n6614);
  and g11866 (n6615, n6613, n_5596);
  and g11867 (n6616, n_5595, n_5596);
  not g11868 (n_5597, n6615);
  not g11869 (n_5598, n6616);
  and g11870 (n6617, n_5597, n_5598);
  and g11871 (n6618, n_5337, n_5343);
  and g11872 (n6619, n6617, n6618);
  not g11873 (n_5599, n6617);
  not g11874 (n_5600, n6618);
  and g11875 (n6620, n_5599, n_5600);
  not g11876 (n_5601, n6619);
  not g11877 (n_5602, n6620);
  and g11878 (n6621, n_5601, n_5602);
  and g11879 (n6622, \b[10] , n4287);
  and g11880 (n6623, \b[8] , n4532);
  and g11881 (n6624, \b[9] , n4282);
  and g11887 (n6627, n738, n4290);
  not g11890 (n_5607, n6628);
  and g11891 (n6629, \a[35] , n_5607);
  not g11892 (n_5608, n6629);
  and g11893 (n6630, \a[35] , n_5608);
  and g11894 (n6631, n_5607, n_5608);
  not g11895 (n_5609, n6630);
  not g11896 (n_5610, n6631);
  and g11897 (n6632, n_5609, n_5610);
  not g11898 (n_5611, n6632);
  and g11899 (n6633, n6621, n_5611);
  not g11900 (n_5612, n6621);
  and g11901 (n6634, n_5612, n6632);
  not g11902 (n_5613, n6561);
  not g11903 (n_5614, n6634);
  and g11904 (n6635, n_5613, n_5614);
  not g11905 (n_5615, n6633);
  and g11906 (n6636, n_5615, n6635);
  not g11907 (n_5616, n6636);
  and g11908 (n6637, n_5613, n_5616);
  and g11909 (n6638, n_5615, n_5616);
  and g11910 (n6639, n_5614, n6638);
  not g11911 (n_5617, n6637);
  not g11912 (n_5618, n6639);
  and g11913 (n6640, n_5617, n_5618);
  and g11914 (n6641, \b[13] , n3638);
  and g11915 (n6642, \b[11] , n3843);
  and g11916 (n6643, \b[12] , n3633);
  and g11922 (n6646, n1008, n3641);
  not g11925 (n_5623, n6647);
  and g11926 (n6648, \a[32] , n_5623);
  not g11927 (n_5624, n6648);
  and g11928 (n6649, \a[32] , n_5624);
  and g11929 (n6650, n_5623, n_5624);
  not g11930 (n_5625, n6649);
  not g11931 (n_5626, n6650);
  and g11932 (n6651, n_5625, n_5626);
  and g11933 (n6652, n6640, n6651);
  not g11934 (n_5627, n6640);
  not g11935 (n_5628, n6651);
  and g11936 (n6653, n_5627, n_5628);
  not g11937 (n_5629, n6652);
  not g11938 (n_5630, n6653);
  and g11939 (n6654, n_5629, n_5630);
  not g11940 (n_5631, n6560);
  and g11941 (n6655, n_5631, n6654);
  not g11942 (n_5632, n6654);
  and g11943 (n6656, n6560, n_5632);
  not g11944 (n_5633, n6655);
  not g11945 (n_5634, n6656);
  and g11946 (n6657, n_5633, n_5634);
  not g11947 (n_5635, n6559);
  and g11948 (n6658, n_5635, n6657);
  not g11949 (n_5636, n6658);
  and g11950 (n6659, n6657, n_5636);
  and g11951 (n6660, n_5635, n_5636);
  not g11952 (n_5637, n6659);
  not g11953 (n_5638, n6660);
  and g11954 (n6661, n_5637, n_5638);
  and g11955 (n6662, n_5382, n_5383);
  not g11956 (n_5639, n6662);
  and g11957 (n6663, n_5379, n_5639);
  and g11958 (n6664, n6661, n6663);
  not g11959 (n_5640, n6661);
  not g11960 (n_5641, n6663);
  and g11961 (n6665, n_5640, n_5641);
  not g11962 (n_5642, n6664);
  not g11963 (n_5643, n6665);
  and g11964 (n6666, n_5642, n_5643);
  and g11965 (n6667, \b[19] , n2539);
  and g11966 (n6668, \b[17] , n2685);
  and g11967 (n6669, \b[18] , n2534);
  and g11973 (n6672, n1708, n2542);
  not g11976 (n_5648, n6673);
  and g11977 (n6674, \a[26] , n_5648);
  not g11978 (n_5649, n6674);
  and g11979 (n6675, \a[26] , n_5649);
  and g11980 (n6676, n_5648, n_5649);
  not g11981 (n_5650, n6675);
  not g11982 (n_5651, n6676);
  and g11983 (n6677, n_5650, n_5651);
  not g11984 (n_5652, n6677);
  and g11985 (n6678, n6666, n_5652);
  not g11986 (n_5653, n6678);
  and g11987 (n6679, n6666, n_5653);
  and g11988 (n6680, n_5652, n_5653);
  not g11989 (n_5654, n6679);
  not g11990 (n_5655, n6680);
  and g11991 (n6681, n_5654, n_5655);
  and g11992 (n6682, n_5396, n_5400);
  and g11993 (n6683, n6681, n6682);
  not g11994 (n_5656, n6681);
  not g11995 (n_5657, n6682);
  and g11996 (n6684, n_5656, n_5657);
  not g11997 (n_5658, n6683);
  not g11998 (n_5659, n6684);
  and g11999 (n6685, n_5658, n_5659);
  and g12000 (n6686, \b[22] , n2048);
  and g12001 (n6687, \b[20] , n2198);
  and g12002 (n6688, \b[21] , n2043);
  and g12008 (n6691, n2051, n2145);
  not g12011 (n_5664, n6692);
  and g12012 (n6693, \a[23] , n_5664);
  not g12013 (n_5665, n6693);
  and g12014 (n6694, \a[23] , n_5665);
  and g12015 (n6695, n_5664, n_5665);
  not g12016 (n_5666, n6694);
  not g12017 (n_5667, n6695);
  and g12018 (n6696, n_5666, n_5667);
  not g12019 (n_5668, n6696);
  and g12020 (n6697, n6685, n_5668);
  not g12021 (n_5669, n6697);
  and g12022 (n6698, n6685, n_5669);
  and g12023 (n6699, n_5668, n_5669);
  not g12024 (n_5670, n6698);
  not g12025 (n_5671, n6699);
  and g12026 (n6700, n_5670, n_5671);
  and g12027 (n6701, n_5403, n_5409);
  and g12028 (n6702, n6700, n6701);
  not g12029 (n_5672, n6700);
  not g12030 (n_5673, n6701);
  and g12031 (n6703, n_5672, n_5673);
  not g12032 (n_5674, n6702);
  not g12033 (n_5675, n6703);
  and g12034 (n6704, n_5674, n_5675);
  and g12035 (n6705, \b[25] , n1627);
  and g12036 (n6706, \b[23] , n1763);
  and g12037 (n6707, \b[24] , n1622);
  and g12043 (n6710, n1630, n2485);
  not g12046 (n_5680, n6711);
  and g12047 (n6712, \a[20] , n_5680);
  not g12048 (n_5681, n6712);
  and g12049 (n6713, \a[20] , n_5681);
  and g12050 (n6714, n_5680, n_5681);
  not g12051 (n_5682, n6713);
  not g12052 (n_5683, n6714);
  and g12053 (n6715, n_5682, n_5683);
  not g12054 (n_5684, n6715);
  and g12055 (n6716, n6704, n_5684);
  not g12056 (n_5685, n6716);
  and g12057 (n6717, n6704, n_5685);
  and g12058 (n6718, n_5684, n_5685);
  not g12059 (n_5686, n6717);
  not g12060 (n_5687, n6718);
  and g12061 (n6719, n_5686, n_5687);
  and g12062 (n6720, n_5421, n_5424);
  not g12063 (n_5688, n6719);
  not g12064 (n_5689, n6720);
  and g12065 (n6721, n_5688, n_5689);
  and g12066 (n6722, n6719, n6720);
  not g12067 (n_5690, n6721);
  not g12068 (n_5691, n6722);
  and g12069 (n6723, n_5690, n_5691);
  not g12070 (n_5692, n6548);
  and g12071 (n6724, n_5692, n6723);
  not g12072 (n_5693, n6724);
  and g12073 (n6725, n_5692, n_5693);
  and g12074 (n6726, n6723, n_5693);
  not g12075 (n_5694, n6725);
  not g12076 (n_5695, n6726);
  and g12077 (n6727, n_5694, n_5695);
  not g12078 (n_5696, n6537);
  not g12079 (n_5697, n6727);
  and g12080 (n6728, n_5696, n_5697);
  not g12081 (n_5698, n6728);
  and g12082 (n6729, n_5696, n_5698);
  and g12083 (n6730, n_5697, n_5698);
  not g12084 (n_5699, n6729);
  not g12085 (n_5700, n6730);
  and g12086 (n6731, n_5699, n_5700);
  and g12087 (n6732, \b[31] , n951);
  and g12088 (n6733, \b[29] , n1056);
  and g12089 (n6734, \b[30] , n946);
  and g12095 (n6737, n954, n3796);
  not g12098 (n_5705, n6738);
  and g12099 (n6739, \a[14] , n_5705);
  not g12100 (n_5706, n6739);
  and g12101 (n6740, \a[14] , n_5706);
  and g12102 (n6741, n_5705, n_5706);
  not g12103 (n_5707, n6740);
  not g12104 (n_5708, n6741);
  and g12105 (n6742, n_5707, n_5708);
  and g12106 (n6743, n6731, n6742);
  not g12107 (n_5709, n6731);
  not g12108 (n_5710, n6742);
  and g12109 (n6744, n_5709, n_5710);
  not g12110 (n_5711, n6743);
  not g12111 (n_5712, n6744);
  and g12112 (n6745, n_5711, n_5712);
  not g12113 (n_5713, n6535);
  and g12114 (n6746, n_5713, n6745);
  not g12115 (n_5714, n6745);
  and g12116 (n6747, n6535, n_5714);
  not g12117 (n_5715, n6746);
  not g12118 (n_5716, n6747);
  and g12119 (n6748, n_5715, n_5716);
  not g12120 (n_5717, n6534);
  and g12121 (n6749, n_5717, n6748);
  not g12122 (n_5718, n6749);
  and g12123 (n6750, n6748, n_5718);
  and g12124 (n6751, n_5717, n_5718);
  not g12125 (n_5719, n6750);
  not g12126 (n_5720, n6751);
  and g12127 (n6752, n_5719, n_5720);
  and g12128 (n6753, n_5454, n_5455);
  not g12129 (n_5721, n6753);
  and g12130 (n6754, n_5451, n_5721);
  and g12131 (n6755, n6752, n6754);
  not g12132 (n_5722, n6752);
  not g12133 (n_5723, n6754);
  and g12134 (n6756, n_5722, n_5723);
  not g12135 (n_5724, n6755);
  not g12136 (n_5725, n6756);
  and g12137 (n6757, n_5724, n_5725);
  and g12138 (n6758, \b[37] , n511);
  and g12139 (n6759, \b[35] , n541);
  and g12140 (n6760, \b[36] , n506);
  and g12146 (n6763, n514, n5181);
  not g12149 (n_5730, n6764);
  and g12150 (n6765, \a[8] , n_5730);
  not g12151 (n_5731, n6765);
  and g12152 (n6766, \a[8] , n_5731);
  and g12153 (n6767, n_5730, n_5731);
  not g12154 (n_5732, n6766);
  not g12155 (n_5733, n6767);
  and g12156 (n6768, n_5732, n_5733);
  not g12157 (n_5734, n6768);
  and g12158 (n6769, n6757, n_5734);
  not g12159 (n_5735, n6757);
  and g12160 (n6770, n_5735, n6768);
  not g12161 (n_5736, n6523);
  not g12162 (n_5737, n6770);
  and g12163 (n6771, n_5736, n_5737);
  not g12164 (n_5738, n6769);
  and g12165 (n6772, n_5738, n6771);
  not g12166 (n_5739, n6772);
  and g12167 (n6773, n_5736, n_5739);
  and g12168 (n6774, n_5738, n_5739);
  and g12169 (n6775, n_5737, n6774);
  not g12170 (n_5740, n6773);
  not g12171 (n_5741, n6775);
  and g12172 (n6776, n_5740, n_5741);
  and g12173 (n6777, \b[40] , n362);
  and g12174 (n6778, \b[38] , n403);
  and g12175 (n6779, \b[39] , n357);
  and g12181 (n6782, n365, n5955);
  not g12184 (n_5746, n6783);
  and g12185 (n6784, \a[5] , n_5746);
  not g12186 (n_5747, n6784);
  and g12187 (n6785, \a[5] , n_5747);
  and g12188 (n6786, n_5746, n_5747);
  not g12189 (n_5748, n6785);
  not g12190 (n_5749, n6786);
  and g12191 (n6787, n_5748, n_5749);
  and g12192 (n6788, n6776, n6787);
  not g12193 (n_5750, n6776);
  not g12194 (n_5751, n6787);
  and g12195 (n6789, n_5750, n_5751);
  not g12196 (n_5752, n6788);
  not g12197 (n_5753, n6789);
  and g12198 (n6790, n_5752, n_5753);
  not g12199 (n_5754, n6522);
  and g12200 (n6791, n_5754, n6790);
  not g12201 (n_5755, n6790);
  and g12202 (n6792, n6522, n_5755);
  not g12203 (n_5756, n6791);
  not g12204 (n_5757, n6792);
  and g12205 (n6793, n_5756, n_5757);
  not g12206 (n_5758, n6521);
  and g12207 (n6794, n_5758, n6793);
  not g12208 (n_5759, n6794);
  and g12209 (n6795, n6793, n_5759);
  and g12210 (n6796, n_5758, n_5759);
  not g12211 (n_5760, n6795);
  not g12212 (n_5761, n6796);
  and g12213 (n6797, n_5760, n_5761);
  and g12214 (n6798, n_5501, n_5506);
  not g12215 (n_5762, n6797);
  not g12216 (n_5763, n6798);
  and g12217 (n6799, n_5762, n_5763);
  and g12218 (n6800, n6797, n6798);
  not g12219 (n_5764, n6799);
  not g12220 (n_5765, n6800);
  and g12221 (\f[43] , n_5764, n_5765);
  and g12222 (n6802, n_5759, n_5764);
  and g12223 (n6803, n_5753, n_5756);
  and g12224 (n6804, \b[41] , n362);
  and g12225 (n6805, \b[39] , n403);
  and g12226 (n6806, \b[40] , n357);
  and g12232 (n6809, n365, n6219);
  not g12235 (n_5770, n6810);
  and g12236 (n6811, \a[5] , n_5770);
  not g12237 (n_5771, n6811);
  and g12238 (n6812, \a[5] , n_5771);
  and g12239 (n6813, n_5770, n_5771);
  not g12240 (n_5772, n6812);
  not g12241 (n_5773, n6813);
  and g12242 (n6814, n_5772, n_5773);
  and g12243 (n6815, \b[35] , n700);
  and g12244 (n6816, \b[33] , n767);
  and g12245 (n6817, \b[34] , n695);
  and g12251 (n6820, n703, n4696);
  not g12254 (n_5778, n6821);
  and g12255 (n6822, \a[11] , n_5778);
  not g12256 (n_5779, n6822);
  and g12257 (n6823, \a[11] , n_5779);
  and g12258 (n6824, n_5778, n_5779);
  not g12259 (n_5780, n6823);
  not g12260 (n_5781, n6824);
  and g12261 (n6825, n_5780, n_5781);
  and g12262 (n6826, n_5712, n_5715);
  and g12263 (n6827, \b[32] , n951);
  and g12264 (n6828, \b[30] , n1056);
  and g12265 (n6829, \b[31] , n946);
  and g12271 (n6832, n954, n4013);
  not g12274 (n_5786, n6833);
  and g12275 (n6834, \a[14] , n_5786);
  not g12276 (n_5787, n6834);
  and g12277 (n6835, \a[14] , n_5787);
  and g12278 (n6836, n_5786, n_5787);
  not g12279 (n_5788, n6835);
  not g12280 (n_5789, n6836);
  and g12281 (n6837, n_5788, n_5789);
  and g12282 (n6838, n_5693, n_5698);
  and g12283 (n6839, \b[29] , n1302);
  and g12284 (n6840, \b[27] , n1391);
  and g12285 (n6841, \b[28] , n1297);
  and g12291 (n6844, n1305, n3383);
  not g12294 (n_5794, n6845);
  and g12295 (n6846, \a[17] , n_5794);
  not g12296 (n_5795, n6846);
  and g12297 (n6847, \a[17] , n_5795);
  and g12298 (n6848, n_5794, n_5795);
  not g12299 (n_5796, n6847);
  not g12300 (n_5797, n6848);
  and g12301 (n6849, n_5796, n_5797);
  and g12302 (n6850, n_5685, n_5690);
  and g12303 (n6851, n_5669, n_5675);
  and g12304 (n6852, \b[20] , n2539);
  and g12305 (n6853, \b[18] , n2685);
  and g12306 (n6854, \b[19] , n2534);
  and g12312 (n6857, n1846, n2542);
  not g12315 (n_5802, n6858);
  and g12316 (n6859, \a[26] , n_5802);
  not g12317 (n_5803, n6859);
  and g12318 (n6860, \a[26] , n_5803);
  and g12319 (n6861, n_5802, n_5803);
  not g12320 (n_5804, n6860);
  not g12321 (n_5805, n6861);
  and g12322 (n6862, n_5804, n_5805);
  and g12323 (n6863, n_5636, n_5643);
  and g12324 (n6864, \b[17] , n3050);
  and g12325 (n6865, \b[15] , n3243);
  and g12326 (n6866, \b[16] , n3045);
  and g12332 (n6869, n1356, n3053);
  not g12335 (n_5810, n6870);
  and g12336 (n6871, \a[29] , n_5810);
  not g12337 (n_5811, n6871);
  and g12338 (n6872, \a[29] , n_5811);
  and g12339 (n6873, n_5810, n_5811);
  not g12340 (n_5812, n6872);
  not g12341 (n_5813, n6873);
  and g12342 (n6874, n_5812, n_5813);
  and g12343 (n6875, n_5630, n_5633);
  and g12344 (n6876, \b[14] , n3638);
  and g12345 (n6877, \b[12] , n3843);
  and g12346 (n6878, \b[13] , n3633);
  and g12352 (n6881, n1034, n3641);
  not g12355 (n_5818, n6882);
  and g12356 (n6883, \a[32] , n_5818);
  not g12357 (n_5819, n6883);
  and g12358 (n6884, \a[32] , n_5819);
  and g12359 (n6885, n_5818, n_5819);
  not g12360 (n_5820, n6884);
  not g12361 (n_5821, n6885);
  and g12362 (n6886, n_5820, n_5821);
  and g12363 (n6887, n_5596, n_5602);
  and g12364 (n6888, \b[8] , n5035);
  and g12365 (n6889, \b[6] , n5277);
  and g12366 (n6890, \b[7] , n5030);
  and g12372 (n6893, n585, n5038);
  not g12375 (n_5826, n6894);
  and g12376 (n6895, \a[38] , n_5826);
  not g12377 (n_5827, n6895);
  and g12378 (n6896, \a[38] , n_5827);
  and g12379 (n6897, n_5826, n_5827);
  not g12380 (n_5828, n6896);
  not g12381 (n_5829, n6897);
  and g12382 (n6898, n_5828, n_5829);
  and g12383 (n6899, n_5590, n_5593);
  and g12384 (n6900, \b[2] , n6595);
  and g12385 (n6901, n6310, n_5577);
  and g12386 (n6902, n6589, n6901);
  and g12387 (n6903, \b[0] , n6902);
  and g12388 (n6904, \b[1] , n6590);
  and g12394 (n6907, n296, n6598);
  not g12397 (n_5834, n6908);
  and g12398 (n6909, \a[44] , n_5834);
  not g12399 (n_5835, n6909);
  and g12400 (n6910, \a[44] , n_5835);
  and g12401 (n6911, n_5834, n_5835);
  not g12402 (n_5836, n6910);
  not g12403 (n_5837, n6911);
  and g12404 (n6912, n_5836, n_5837);
  and g12405 (n6913, n_5585, n6912);
  not g12406 (n_5838, n6912);
  and g12407 (n6914, n6605, n_5838);
  not g12408 (n_5839, n6913);
  not g12409 (n_5840, n6914);
  and g12410 (n6915, n_5839, n_5840);
  and g12411 (n6916, \b[5] , n5777);
  and g12412 (n6917, \b[3] , n6059);
  and g12413 (n6918, \b[4] , n5772);
  and g12419 (n6921, n394, n5780);
  not g12422 (n_5845, n6922);
  and g12423 (n6923, \a[41] , n_5845);
  not g12424 (n_5846, n6923);
  and g12425 (n6924, \a[41] , n_5846);
  and g12426 (n6925, n_5845, n_5846);
  not g12427 (n_5847, n6924);
  not g12428 (n_5848, n6925);
  and g12429 (n6926, n_5847, n_5848);
  not g12430 (n_5849, n6926);
  and g12431 (n6927, n6915, n_5849);
  not g12432 (n_5850, n6927);
  and g12433 (n6928, n6915, n_5850);
  and g12434 (n6929, n_5849, n_5850);
  not g12435 (n_5851, n6928);
  not g12436 (n_5852, n6929);
  and g12437 (n6930, n_5851, n_5852);
  not g12438 (n_5853, n6899);
  not g12439 (n_5854, n6930);
  and g12440 (n6931, n_5853, n_5854);
  and g12441 (n6932, n6899, n6930);
  not g12442 (n_5855, n6931);
  not g12443 (n_5856, n6932);
  and g12444 (n6933, n_5855, n_5856);
  not g12445 (n_5857, n6898);
  and g12446 (n6934, n_5857, n6933);
  not g12447 (n_5858, n6934);
  and g12448 (n6935, n_5857, n_5858);
  and g12449 (n6936, n6933, n_5858);
  not g12450 (n_5859, n6935);
  not g12451 (n_5860, n6936);
  and g12452 (n6937, n_5859, n_5860);
  not g12453 (n_5861, n6887);
  not g12454 (n_5862, n6937);
  and g12455 (n6938, n_5861, n_5862);
  not g12456 (n_5863, n6938);
  and g12457 (n6939, n_5861, n_5863);
  and g12458 (n6940, n_5862, n_5863);
  not g12459 (n_5864, n6939);
  not g12460 (n_5865, n6940);
  and g12461 (n6941, n_5864, n_5865);
  and g12462 (n6942, \b[11] , n4287);
  and g12463 (n6943, \b[9] , n4532);
  and g12464 (n6944, \b[10] , n4282);
  and g12470 (n6947, n818, n4290);
  not g12473 (n_5870, n6948);
  and g12474 (n6949, \a[35] , n_5870);
  not g12475 (n_5871, n6949);
  and g12476 (n6950, \a[35] , n_5871);
  and g12477 (n6951, n_5870, n_5871);
  not g12478 (n_5872, n6950);
  not g12479 (n_5873, n6951);
  and g12480 (n6952, n_5872, n_5873);
  and g12481 (n6953, n6941, n6952);
  not g12482 (n_5874, n6941);
  not g12483 (n_5875, n6952);
  and g12484 (n6954, n_5874, n_5875);
  not g12485 (n_5876, n6953);
  not g12486 (n_5877, n6954);
  and g12487 (n6955, n_5876, n_5877);
  not g12488 (n_5878, n6638);
  and g12489 (n6956, n_5878, n6955);
  not g12490 (n_5879, n6955);
  and g12491 (n6957, n6638, n_5879);
  not g12492 (n_5880, n6956);
  not g12493 (n_5881, n6957);
  and g12494 (n6958, n_5880, n_5881);
  not g12495 (n_5882, n6958);
  and g12496 (n6959, n6886, n_5882);
  not g12497 (n_5883, n6886);
  and g12498 (n6960, n_5883, n6958);
  not g12499 (n_5884, n6959);
  not g12500 (n_5885, n6960);
  and g12501 (n6961, n_5884, n_5885);
  not g12502 (n_5886, n6875);
  and g12503 (n6962, n_5886, n6961);
  not g12504 (n_5887, n6961);
  and g12505 (n6963, n6875, n_5887);
  not g12506 (n_5888, n6962);
  not g12507 (n_5889, n6963);
  and g12508 (n6964, n_5888, n_5889);
  not g12509 (n_5890, n6964);
  and g12510 (n6965, n6874, n_5890);
  not g12511 (n_5891, n6874);
  and g12512 (n6966, n_5891, n6964);
  not g12513 (n_5892, n6965);
  not g12514 (n_5893, n6966);
  and g12515 (n6967, n_5892, n_5893);
  not g12516 (n_5894, n6863);
  and g12517 (n6968, n_5894, n6967);
  not g12518 (n_5895, n6967);
  and g12519 (n6969, n6863, n_5895);
  not g12520 (n_5896, n6968);
  not g12521 (n_5897, n6969);
  and g12522 (n6970, n_5896, n_5897);
  not g12523 (n_5898, n6862);
  and g12524 (n6971, n_5898, n6970);
  not g12525 (n_5899, n6971);
  and g12526 (n6972, n6970, n_5899);
  and g12527 (n6973, n_5898, n_5899);
  not g12528 (n_5900, n6972);
  not g12529 (n_5901, n6973);
  and g12530 (n6974, n_5900, n_5901);
  and g12531 (n6975, n_5653, n_5659);
  and g12532 (n6976, n6974, n6975);
  not g12533 (n_5902, n6974);
  not g12534 (n_5903, n6975);
  and g12535 (n6977, n_5902, n_5903);
  not g12536 (n_5904, n6976);
  not g12537 (n_5905, n6977);
  and g12538 (n6978, n_5904, n_5905);
  and g12539 (n6979, \b[23] , n2048);
  and g12540 (n6980, \b[21] , n2198);
  and g12541 (n6981, \b[22] , n2043);
  and g12547 (n6984, n2051, n2300);
  not g12550 (n_5910, n6985);
  and g12551 (n6986, \a[23] , n_5910);
  not g12552 (n_5911, n6986);
  and g12553 (n6987, \a[23] , n_5911);
  and g12554 (n6988, n_5910, n_5911);
  not g12555 (n_5912, n6987);
  not g12556 (n_5913, n6988);
  and g12557 (n6989, n_5912, n_5913);
  not g12558 (n_5914, n6989);
  and g12559 (n6990, n6978, n_5914);
  not g12560 (n_5915, n6978);
  and g12561 (n6991, n_5915, n6989);
  not g12562 (n_5916, n6851);
  not g12563 (n_5917, n6991);
  and g12564 (n6992, n_5916, n_5917);
  not g12565 (n_5918, n6990);
  and g12566 (n6993, n_5918, n6992);
  not g12567 (n_5919, n6993);
  and g12568 (n6994, n_5916, n_5919);
  and g12569 (n6995, n_5918, n_5919);
  and g12570 (n6996, n_5917, n6995);
  not g12571 (n_5920, n6994);
  not g12572 (n_5921, n6996);
  and g12573 (n6997, n_5920, n_5921);
  and g12574 (n6998, \b[26] , n1627);
  and g12575 (n6999, \b[24] , n1763);
  and g12576 (n7000, \b[25] , n1622);
  and g12582 (n7003, n1630, n2813);
  not g12585 (n_5926, n7004);
  and g12586 (n7005, \a[20] , n_5926);
  not g12587 (n_5927, n7005);
  and g12588 (n7006, \a[20] , n_5927);
  and g12589 (n7007, n_5926, n_5927);
  not g12590 (n_5928, n7006);
  not g12591 (n_5929, n7007);
  and g12592 (n7008, n_5928, n_5929);
  and g12593 (n7009, n6997, n7008);
  not g12594 (n_5930, n6997);
  not g12595 (n_5931, n7008);
  and g12596 (n7010, n_5930, n_5931);
  not g12597 (n_5932, n7009);
  not g12598 (n_5933, n7010);
  and g12599 (n7011, n_5932, n_5933);
  not g12600 (n_5934, n6850);
  and g12601 (n7012, n_5934, n7011);
  not g12602 (n_5935, n7011);
  and g12603 (n7013, n6850, n_5935);
  not g12604 (n_5936, n7012);
  not g12605 (n_5937, n7013);
  and g12606 (n7014, n_5936, n_5937);
  not g12607 (n_5938, n7014);
  and g12608 (n7015, n6849, n_5938);
  not g12609 (n_5939, n6849);
  and g12610 (n7016, n_5939, n7014);
  not g12611 (n_5940, n7015);
  not g12612 (n_5941, n7016);
  and g12613 (n7017, n_5940, n_5941);
  not g12614 (n_5942, n6838);
  and g12615 (n7018, n_5942, n7017);
  not g12616 (n_5943, n7017);
  and g12617 (n7019, n6838, n_5943);
  not g12618 (n_5944, n7018);
  not g12619 (n_5945, n7019);
  and g12620 (n7020, n_5944, n_5945);
  not g12621 (n_5946, n7020);
  and g12622 (n7021, n6837, n_5946);
  not g12623 (n_5947, n6837);
  and g12624 (n7022, n_5947, n7020);
  not g12625 (n_5948, n7021);
  not g12626 (n_5949, n7022);
  and g12627 (n7023, n_5948, n_5949);
  not g12628 (n_5950, n6826);
  and g12629 (n7024, n_5950, n7023);
  not g12630 (n_5951, n7023);
  and g12631 (n7025, n6826, n_5951);
  not g12632 (n_5952, n7024);
  not g12633 (n_5953, n7025);
  and g12634 (n7026, n_5952, n_5953);
  not g12635 (n_5954, n6825);
  and g12636 (n7027, n_5954, n7026);
  not g12637 (n_5955, n7027);
  and g12638 (n7028, n7026, n_5955);
  and g12639 (n7029, n_5954, n_5955);
  not g12640 (n_5956, n7028);
  not g12641 (n_5957, n7029);
  and g12642 (n7030, n_5956, n_5957);
  and g12643 (n7031, n_5718, n_5725);
  and g12644 (n7032, n7030, n7031);
  not g12645 (n_5958, n7030);
  not g12646 (n_5959, n7031);
  and g12647 (n7033, n_5958, n_5959);
  not g12648 (n_5960, n7032);
  not g12649 (n_5961, n7033);
  and g12650 (n7034, n_5960, n_5961);
  and g12651 (n7035, \b[38] , n511);
  and g12652 (n7036, \b[36] , n541);
  and g12653 (n7037, \b[37] , n506);
  and g12659 (n7040, n514, n5205);
  not g12662 (n_5966, n7041);
  and g12663 (n7042, \a[8] , n_5966);
  not g12664 (n_5967, n7042);
  and g12665 (n7043, \a[8] , n_5967);
  and g12666 (n7044, n_5966, n_5967);
  not g12667 (n_5968, n7043);
  not g12668 (n_5969, n7044);
  and g12669 (n7045, n_5968, n_5969);
  not g12670 (n_5970, n7045);
  and g12671 (n7046, n7034, n_5970);
  not g12672 (n_5971, n7046);
  and g12673 (n7047, n7034, n_5971);
  and g12674 (n7048, n_5970, n_5971);
  not g12675 (n_5972, n7047);
  not g12676 (n_5973, n7048);
  and g12677 (n7049, n_5972, n_5973);
  not g12678 (n_5974, n6774);
  not g12679 (n_5975, n7049);
  and g12680 (n7050, n_5974, n_5975);
  and g12681 (n7051, n6774, n7049);
  not g12682 (n_5976, n7050);
  not g12683 (n_5977, n7051);
  and g12684 (n7052, n_5976, n_5977);
  not g12685 (n_5978, n6814);
  and g12686 (n7053, n_5978, n7052);
  not g12687 (n_5979, n7053);
  and g12688 (n7054, n_5978, n_5979);
  and g12689 (n7055, n7052, n_5979);
  not g12690 (n_5980, n7054);
  not g12691 (n_5981, n7055);
  and g12692 (n7056, n_5980, n_5981);
  not g12693 (n_5982, n6803);
  not g12694 (n_5983, n7056);
  and g12695 (n7057, n_5982, n_5983);
  not g12696 (n_5984, n7057);
  and g12697 (n7058, n_5982, n_5984);
  and g12698 (n7059, n_5983, n_5984);
  not g12699 (n_5985, n7058);
  not g12700 (n_5986, n7059);
  and g12701 (n7060, n_5985, n_5986);
  and g12702 (n7061, \b[44] , n266);
  and g12703 (n7062, \b[42] , n284);
  and g12704 (n7063, \b[43] , n261);
  and g12710 (n7066, n_5514, n_5517);
  not g12711 (n_5991, \b[44] );
  and g12712 (n7067, n_5512, n_5991);
  and g12713 (n7068, \b[43] , \b[44] );
  not g12714 (n_5992, n7067);
  not g12715 (n_5993, n7068);
  and g12716 (n7069, n_5992, n_5993);
  not g12717 (n_5994, n7066);
  and g12718 (n7070, n_5994, n7069);
  not g12719 (n_5995, n7069);
  and g12720 (n7071, n7066, n_5995);
  not g12721 (n_5996, n7070);
  not g12722 (n_5997, n7071);
  and g12723 (n7072, n_5996, n_5997);
  and g12724 (n7073, n269, n7072);
  not g12727 (n_5999, n7074);
  and g12728 (n7075, \a[2] , n_5999);
  not g12729 (n_6000, n7075);
  and g12730 (n7076, \a[2] , n_6000);
  and g12731 (n7077, n_5999, n_6000);
  not g12732 (n_6001, n7076);
  not g12733 (n_6002, n7077);
  and g12734 (n7078, n_6001, n_6002);
  not g12735 (n_6003, n7060);
  and g12736 (n7079, n_6003, n7078);
  not g12737 (n_6004, n7078);
  and g12738 (n7080, n7060, n_6004);
  not g12739 (n_6005, n7079);
  not g12740 (n_6006, n7080);
  and g12741 (n7081, n_6005, n_6006);
  not g12742 (n_6007, n6802);
  not g12743 (n_6008, n7081);
  and g12744 (n7082, n_6007, n_6008);
  and g12745 (n7083, n6802, n7081);
  not g12746 (n_6009, n7082);
  not g12747 (n_6010, n7083);
  and g12748 (\f[44] , n_6009, n_6010);
  and g12749 (n7085, n_6003, n_6004);
  not g12750 (n_6011, n7085);
  and g12751 (n7086, n_6009, n_6011);
  and g12752 (n7087, n_5955, n_5961);
  and g12753 (n7088, n_5949, n_5952);
  and g12754 (n7089, \b[33] , n951);
  and g12755 (n7090, \b[31] , n1056);
  and g12756 (n7091, \b[32] , n946);
  and g12762 (n7094, n954, n4223);
  not g12765 (n_6016, n7095);
  and g12766 (n7096, \a[14] , n_6016);
  not g12767 (n_6017, n7096);
  and g12768 (n7097, \a[14] , n_6017);
  and g12769 (n7098, n_6016, n_6017);
  not g12770 (n_6018, n7097);
  not g12771 (n_6019, n7098);
  and g12772 (n7099, n_6018, n_6019);
  and g12773 (n7100, n_5941, n_5944);
  and g12774 (n7101, n_5933, n_5936);
  and g12775 (n7102, \b[27] , n1627);
  and g12776 (n7103, \b[25] , n1763);
  and g12777 (n7104, \b[26] , n1622);
  and g12783 (n7107, n1630, n2990);
  not g12786 (n_6024, n7108);
  and g12787 (n7109, \a[20] , n_6024);
  not g12788 (n_6025, n7109);
  and g12789 (n7110, \a[20] , n_6025);
  and g12790 (n7111, n_6024, n_6025);
  not g12791 (n_6026, n7110);
  not g12792 (n_6027, n7111);
  and g12793 (n7112, n_6026, n_6027);
  and g12794 (n7113, \b[21] , n2539);
  and g12795 (n7114, \b[19] , n2685);
  and g12796 (n7115, \b[20] , n2534);
  and g12802 (n7118, n1984, n2542);
  not g12805 (n_6032, n7119);
  and g12806 (n7120, \a[26] , n_6032);
  not g12807 (n_6033, n7120);
  and g12808 (n7121, \a[26] , n_6033);
  and g12809 (n7122, n_6032, n_6033);
  not g12810 (n_6034, n7121);
  not g12811 (n_6035, n7122);
  and g12812 (n7123, n_6034, n_6035);
  and g12813 (n7124, n_5893, n_5896);
  and g12814 (n7125, n_5885, n_5888);
  and g12815 (n7126, n_5877, n_5880);
  and g12816 (n7127, \b[12] , n4287);
  and g12817 (n7128, \b[10] , n4532);
  and g12818 (n7129, \b[11] , n4282);
  and g12824 (n7132, n842, n4290);
  not g12827 (n_6040, n7133);
  and g12828 (n7134, \a[35] , n_6040);
  not g12829 (n_6041, n7134);
  and g12830 (n7135, \a[35] , n_6041);
  and g12831 (n7136, n_6040, n_6041);
  not g12832 (n_6042, n7135);
  not g12833 (n_6043, n7136);
  and g12834 (n7137, n_6042, n_6043);
  and g12835 (n7138, n_5858, n_5863);
  and g12836 (n7139, \b[6] , n5777);
  and g12837 (n7140, \b[4] , n6059);
  and g12838 (n7141, \b[5] , n5772);
  and g12844 (n7144, n459, n5780);
  not g12847 (n_6048, n7145);
  and g12848 (n7146, \a[41] , n_6048);
  not g12849 (n_6049, n7146);
  and g12850 (n7147, \a[41] , n_6049);
  and g12851 (n7148, n_6048, n_6049);
  not g12852 (n_6050, n7147);
  not g12853 (n_6051, n7148);
  and g12854 (n7149, n_6050, n_6051);
  not g12855 (n_6053, \a[45] );
  and g12856 (n7150, \a[44] , n_6053);
  and g12857 (n7151, n_5572, \a[45] );
  not g12858 (n_6054, n7150);
  not g12859 (n_6055, n7151);
  and g12860 (n7152, n_6054, n_6055);
  not g12861 (n_6056, n7152);
  and g12862 (n7153, \b[0] , n_6056);
  and g12863 (n7154, n_5840, n7153);
  not g12864 (n_6057, n7153);
  and g12865 (n7155, n6914, n_6057);
  not g12866 (n_6058, n7154);
  not g12867 (n_6059, n7155);
  and g12868 (n7156, n_6058, n_6059);
  and g12869 (n7157, \b[3] , n6595);
  and g12870 (n7158, \b[1] , n6902);
  and g12871 (n7159, \b[2] , n6590);
  and g12877 (n7162, n318, n6598);
  not g12880 (n_6064, n7163);
  and g12881 (n7164, \a[44] , n_6064);
  not g12882 (n_6065, n7164);
  and g12883 (n7165, \a[44] , n_6065);
  and g12884 (n7166, n_6064, n_6065);
  not g12885 (n_6066, n7165);
  not g12886 (n_6067, n7166);
  and g12887 (n7167, n_6066, n_6067);
  not g12888 (n_6068, n7156);
  not g12889 (n_6069, n7167);
  and g12890 (n7168, n_6068, n_6069);
  and g12891 (n7169, n7156, n7167);
  not g12892 (n_6070, n7168);
  not g12893 (n_6071, n7169);
  and g12894 (n7170, n_6070, n_6071);
  not g12895 (n_6072, n7149);
  and g12896 (n7171, n_6072, n7170);
  not g12897 (n_6073, n7171);
  and g12898 (n7172, n7170, n_6073);
  and g12899 (n7173, n_6072, n_6073);
  not g12900 (n_6074, n7172);
  not g12901 (n_6075, n7173);
  and g12902 (n7174, n_6074, n_6075);
  and g12903 (n7175, n_5850, n_5855);
  and g12904 (n7176, n7174, n7175);
  not g12905 (n_6076, n7174);
  not g12906 (n_6077, n7175);
  and g12907 (n7177, n_6076, n_6077);
  not g12908 (n_6078, n7176);
  not g12909 (n_6079, n7177);
  and g12910 (n7178, n_6078, n_6079);
  and g12911 (n7179, \b[9] , n5035);
  and g12912 (n7180, \b[7] , n5277);
  and g12913 (n7181, \b[8] , n5030);
  and g12919 (n7184, n651, n5038);
  not g12922 (n_6084, n7185);
  and g12923 (n7186, \a[38] , n_6084);
  not g12924 (n_6085, n7186);
  and g12925 (n7187, \a[38] , n_6085);
  and g12926 (n7188, n_6084, n_6085);
  not g12927 (n_6086, n7187);
  not g12928 (n_6087, n7188);
  and g12929 (n7189, n_6086, n_6087);
  not g12930 (n_6088, n7178);
  and g12931 (n7190, n_6088, n7189);
  not g12932 (n_6089, n7189);
  and g12933 (n7191, n7178, n_6089);
  not g12934 (n_6090, n7190);
  not g12935 (n_6091, n7191);
  and g12936 (n7192, n_6090, n_6091);
  not g12937 (n_6092, n7138);
  and g12938 (n7193, n_6092, n7192);
  not g12939 (n_6093, n7192);
  and g12940 (n7194, n7138, n_6093);
  not g12941 (n_6094, n7193);
  not g12942 (n_6095, n7194);
  and g12943 (n7195, n_6094, n_6095);
  not g12944 (n_6096, n7137);
  and g12945 (n7196, n_6096, n7195);
  not g12946 (n_6097, n7196);
  and g12947 (n7197, n_6096, n_6097);
  and g12948 (n7198, n7195, n_6097);
  not g12949 (n_6098, n7197);
  not g12950 (n_6099, n7198);
  and g12951 (n7199, n_6098, n_6099);
  not g12952 (n_6100, n7126);
  not g12953 (n_6101, n7199);
  and g12954 (n7200, n_6100, n_6101);
  not g12955 (n_6102, n7200);
  and g12956 (n7201, n_6100, n_6102);
  and g12957 (n7202, n_6101, n_6102);
  not g12958 (n_6103, n7201);
  not g12959 (n_6104, n7202);
  and g12960 (n7203, n_6103, n_6104);
  and g12961 (n7204, \b[15] , n3638);
  and g12962 (n7205, \b[13] , n3843);
  and g12963 (n7206, \b[14] , n3633);
  and g12969 (n7209, n1131, n3641);
  not g12972 (n_6109, n7210);
  and g12973 (n7211, \a[32] , n_6109);
  not g12974 (n_6110, n7211);
  and g12975 (n7212, \a[32] , n_6110);
  and g12976 (n7213, n_6109, n_6110);
  not g12977 (n_6111, n7212);
  not g12978 (n_6112, n7213);
  and g12979 (n7214, n_6111, n_6112);
  not g12980 (n_6113, n7203);
  not g12981 (n_6114, n7214);
  and g12982 (n7215, n_6113, n_6114);
  not g12983 (n_6115, n7215);
  and g12984 (n7216, n_6113, n_6115);
  and g12985 (n7217, n_6114, n_6115);
  not g12986 (n_6116, n7216);
  not g12987 (n_6117, n7217);
  and g12988 (n7218, n_6116, n_6117);
  not g12989 (n_6118, n7125);
  and g12990 (n7219, n_6118, n7218);
  not g12991 (n_6119, n7218);
  and g12992 (n7220, n7125, n_6119);
  not g12993 (n_6120, n7219);
  not g12994 (n_6121, n7220);
  and g12995 (n7221, n_6120, n_6121);
  and g12996 (n7222, \b[18] , n3050);
  and g12997 (n7223, \b[16] , n3243);
  and g12998 (n7224, \b[17] , n3045);
  and g13004 (n7227, n1566, n3053);
  not g13007 (n_6126, n7228);
  and g13008 (n7229, \a[29] , n_6126);
  not g13009 (n_6127, n7229);
  and g13010 (n7230, \a[29] , n_6127);
  and g13011 (n7231, n_6126, n_6127);
  not g13012 (n_6128, n7230);
  not g13013 (n_6129, n7231);
  and g13014 (n7232, n_6128, n_6129);
  not g13015 (n_6130, n7221);
  not g13016 (n_6131, n7232);
  and g13017 (n7233, n_6130, n_6131);
  and g13018 (n7234, n7221, n7232);
  not g13019 (n_6132, n7233);
  not g13020 (n_6133, n7234);
  and g13021 (n7235, n_6132, n_6133);
  not g13022 (n_6134, n7124);
  and g13023 (n7236, n_6134, n7235);
  not g13024 (n_6135, n7235);
  and g13025 (n7237, n7124, n_6135);
  not g13026 (n_6136, n7236);
  not g13027 (n_6137, n7237);
  and g13028 (n7238, n_6136, n_6137);
  not g13029 (n_6138, n7123);
  and g13030 (n7239, n_6138, n7238);
  not g13031 (n_6139, n7239);
  and g13032 (n7240, n7238, n_6139);
  and g13033 (n7241, n_6138, n_6139);
  not g13034 (n_6140, n7240);
  not g13035 (n_6141, n7241);
  and g13036 (n7242, n_6140, n_6141);
  and g13037 (n7243, n_5899, n_5905);
  and g13038 (n7244, n7242, n7243);
  not g13039 (n_6142, n7242);
  not g13040 (n_6143, n7243);
  and g13041 (n7245, n_6142, n_6143);
  not g13042 (n_6144, n7244);
  not g13043 (n_6145, n7245);
  and g13044 (n7246, n_6144, n_6145);
  and g13045 (n7247, \b[24] , n2048);
  and g13046 (n7248, \b[22] , n2198);
  and g13047 (n7249, \b[23] , n2043);
  and g13053 (n7252, n2051, n2458);
  not g13056 (n_6150, n7253);
  and g13057 (n7254, \a[23] , n_6150);
  not g13058 (n_6151, n7254);
  and g13059 (n7255, \a[23] , n_6151);
  and g13060 (n7256, n_6150, n_6151);
  not g13061 (n_6152, n7255);
  not g13062 (n_6153, n7256);
  and g13063 (n7257, n_6152, n_6153);
  not g13064 (n_6154, n7246);
  and g13065 (n7258, n_6154, n7257);
  not g13066 (n_6155, n7257);
  and g13067 (n7259, n7246, n_6155);
  not g13068 (n_6156, n7258);
  not g13069 (n_6157, n7259);
  and g13070 (n7260, n_6156, n_6157);
  not g13071 (n_6158, n6995);
  and g13072 (n7261, n_6158, n7260);
  not g13073 (n_6159, n7260);
  and g13074 (n7262, n6995, n_6159);
  not g13075 (n_6160, n7261);
  not g13076 (n_6161, n7262);
  and g13077 (n7263, n_6160, n_6161);
  not g13078 (n_6162, n7112);
  and g13079 (n7264, n_6162, n7263);
  not g13080 (n_6163, n7264);
  and g13081 (n7265, n7263, n_6163);
  and g13082 (n7266, n_6162, n_6163);
  not g13083 (n_6164, n7265);
  not g13084 (n_6165, n7266);
  and g13085 (n7267, n_6164, n_6165);
  not g13086 (n_6166, n7101);
  and g13087 (n7268, n_6166, n7267);
  not g13088 (n_6167, n7267);
  and g13089 (n7269, n7101, n_6167);
  not g13090 (n_6168, n7268);
  not g13091 (n_6169, n7269);
  and g13092 (n7270, n_6168, n_6169);
  and g13093 (n7271, \b[30] , n1302);
  and g13094 (n7272, \b[28] , n1391);
  and g13095 (n7273, \b[29] , n1297);
  and g13101 (n7276, n1305, n3577);
  not g13104 (n_6174, n7277);
  and g13105 (n7278, \a[17] , n_6174);
  not g13106 (n_6175, n7278);
  and g13107 (n7279, \a[17] , n_6175);
  and g13108 (n7280, n_6174, n_6175);
  not g13109 (n_6176, n7279);
  not g13110 (n_6177, n7280);
  and g13111 (n7281, n_6176, n_6177);
  not g13112 (n_6178, n7270);
  not g13113 (n_6179, n7281);
  and g13114 (n7282, n_6178, n_6179);
  and g13115 (n7283, n7270, n7281);
  not g13116 (n_6180, n7282);
  not g13117 (n_6181, n7283);
  and g13118 (n7284, n_6180, n_6181);
  not g13119 (n_6182, n7100);
  and g13120 (n7285, n_6182, n7284);
  not g13121 (n_6183, n7284);
  and g13122 (n7286, n7100, n_6183);
  not g13123 (n_6184, n7285);
  not g13124 (n_6185, n7286);
  and g13125 (n7287, n_6184, n_6185);
  not g13126 (n_6186, n7099);
  and g13127 (n7288, n_6186, n7287);
  not g13128 (n_6187, n7288);
  and g13129 (n7289, n7287, n_6187);
  and g13130 (n7290, n_6186, n_6187);
  not g13131 (n_6188, n7289);
  not g13132 (n_6189, n7290);
  and g13133 (n7291, n_6188, n_6189);
  not g13134 (n_6190, n7088);
  and g13135 (n7292, n_6190, n7291);
  not g13136 (n_6191, n7291);
  and g13137 (n7293, n7088, n_6191);
  not g13138 (n_6192, n7292);
  not g13139 (n_6193, n7293);
  and g13140 (n7294, n_6192, n_6193);
  and g13141 (n7295, \b[36] , n700);
  and g13142 (n7296, \b[34] , n767);
  and g13143 (n7297, \b[35] , n695);
  and g13149 (n7300, n703, n4922);
  not g13152 (n_6198, n7301);
  and g13153 (n7302, \a[11] , n_6198);
  not g13154 (n_6199, n7302);
  and g13155 (n7303, \a[11] , n_6199);
  and g13156 (n7304, n_6198, n_6199);
  not g13157 (n_6200, n7303);
  not g13158 (n_6201, n7304);
  and g13159 (n7305, n_6200, n_6201);
  not g13160 (n_6202, n7294);
  not g13161 (n_6203, n7305);
  and g13162 (n7306, n_6202, n_6203);
  and g13163 (n7307, n7294, n7305);
  not g13164 (n_6204, n7306);
  not g13165 (n_6205, n7307);
  and g13166 (n7308, n_6204, n_6205);
  not g13167 (n_6206, n7308);
  and g13168 (n7309, n7087, n_6206);
  not g13169 (n_6207, n7087);
  and g13170 (n7310, n_6207, n7308);
  not g13171 (n_6208, n7309);
  not g13172 (n_6209, n7310);
  and g13173 (n7311, n_6208, n_6209);
  and g13174 (n7312, \b[39] , n511);
  and g13175 (n7313, \b[37] , n541);
  and g13176 (n7314, \b[38] , n506);
  and g13182 (n7317, n514, n5451);
  not g13185 (n_6214, n7318);
  and g13186 (n7319, \a[8] , n_6214);
  not g13187 (n_6215, n7319);
  and g13188 (n7320, \a[8] , n_6215);
  and g13189 (n7321, n_6214, n_6215);
  not g13190 (n_6216, n7320);
  not g13191 (n_6217, n7321);
  and g13192 (n7322, n_6216, n_6217);
  not g13193 (n_6218, n7322);
  and g13194 (n7323, n7311, n_6218);
  not g13195 (n_6219, n7323);
  and g13196 (n7324, n7311, n_6219);
  and g13197 (n7325, n_6218, n_6219);
  not g13198 (n_6220, n7324);
  not g13199 (n_6221, n7325);
  and g13200 (n7326, n_6220, n_6221);
  and g13201 (n7327, n_5971, n_5976);
  and g13202 (n7328, n7326, n7327);
  not g13203 (n_6222, n7326);
  not g13204 (n_6223, n7327);
  and g13205 (n7329, n_6222, n_6223);
  not g13206 (n_6224, n7328);
  not g13207 (n_6225, n7329);
  and g13208 (n7330, n_6224, n_6225);
  and g13209 (n7331, \b[42] , n362);
  and g13210 (n7332, \b[40] , n403);
  and g13211 (n7333, \b[41] , n357);
  and g13217 (n7336, n365, n6489);
  not g13220 (n_6230, n7337);
  and g13221 (n7338, \a[5] , n_6230);
  not g13222 (n_6231, n7338);
  and g13223 (n7339, \a[5] , n_6231);
  and g13224 (n7340, n_6230, n_6231);
  not g13225 (n_6232, n7339);
  not g13226 (n_6233, n7340);
  and g13227 (n7341, n_6232, n_6233);
  not g13228 (n_6234, n7341);
  and g13229 (n7342, n7330, n_6234);
  not g13230 (n_6235, n7342);
  and g13231 (n7343, n7330, n_6235);
  and g13232 (n7344, n_6234, n_6235);
  not g13233 (n_6236, n7343);
  not g13234 (n_6237, n7344);
  and g13235 (n7345, n_6236, n_6237);
  and g13236 (n7346, n_5979, n_5984);
  and g13237 (n7347, n7345, n7346);
  not g13238 (n_6238, n7345);
  not g13239 (n_6239, n7346);
  and g13240 (n7348, n_6238, n_6239);
  not g13241 (n_6240, n7347);
  not g13242 (n_6241, n7348);
  and g13243 (n7349, n_6240, n_6241);
  and g13244 (n7350, \b[45] , n266);
  and g13245 (n7351, \b[43] , n284);
  and g13246 (n7352, \b[44] , n261);
  and g13252 (n7355, n_5993, n_5996);
  not g13253 (n_6246, \b[45] );
  and g13254 (n7356, n_5991, n_6246);
  and g13255 (n7357, \b[44] , \b[45] );
  not g13256 (n_6247, n7356);
  not g13257 (n_6248, n7357);
  and g13258 (n7358, n_6247, n_6248);
  not g13259 (n_6249, n7355);
  and g13260 (n7359, n_6249, n7358);
  not g13261 (n_6250, n7358);
  and g13262 (n7360, n7355, n_6250);
  not g13263 (n_6251, n7359);
  not g13264 (n_6252, n7360);
  and g13265 (n7361, n_6251, n_6252);
  and g13266 (n7362, n269, n7361);
  not g13269 (n_6254, n7363);
  and g13270 (n7364, \a[2] , n_6254);
  not g13271 (n_6255, n7364);
  and g13272 (n7365, \a[2] , n_6255);
  and g13273 (n7366, n_6254, n_6255);
  not g13274 (n_6256, n7365);
  not g13275 (n_6257, n7366);
  and g13276 (n7367, n_6256, n_6257);
  not g13277 (n_6258, n7349);
  and g13278 (n7368, n_6258, n7367);
  not g13279 (n_6259, n7367);
  and g13280 (n7369, n7349, n_6259);
  not g13281 (n_6260, n7368);
  not g13282 (n_6261, n7369);
  and g13283 (n7370, n_6260, n_6261);
  not g13284 (n_6262, n7086);
  and g13285 (n7371, n_6262, n7370);
  not g13286 (n_6263, n7370);
  and g13287 (n7372, n7086, n_6263);
  not g13288 (n_6264, n7371);
  not g13289 (n_6265, n7372);
  and g13290 (\f[45] , n_6264, n_6265);
  and g13291 (n7374, n_6219, n_6225);
  and g13292 (n7375, \b[34] , n951);
  and g13293 (n7376, \b[32] , n1056);
  and g13294 (n7377, \b[33] , n946);
  and g13300 (n7380, n954, n4466);
  not g13303 (n_6270, n7381);
  and g13304 (n7382, \a[14] , n_6270);
  not g13305 (n_6271, n7382);
  and g13306 (n7383, \a[14] , n_6271);
  and g13307 (n7384, n_6270, n_6271);
  not g13308 (n_6272, n7383);
  not g13309 (n_6273, n7384);
  and g13310 (n7385, n_6272, n_6273);
  and g13311 (n7386, n_6180, n_6184);
  and g13312 (n7387, n_6166, n_6167);
  not g13313 (n_6274, n7387);
  and g13314 (n7388, n_6163, n_6274);
  and g13315 (n7389, \b[28] , n1627);
  and g13316 (n7390, \b[26] , n1763);
  and g13317 (n7391, \b[27] , n1622);
  and g13323 (n7394, n1630, n3189);
  not g13326 (n_6279, n7395);
  and g13327 (n7396, \a[20] , n_6279);
  not g13328 (n_6280, n7396);
  and g13329 (n7397, \a[20] , n_6280);
  and g13330 (n7398, n_6279, n_6280);
  not g13331 (n_6281, n7397);
  not g13332 (n_6282, n7398);
  and g13333 (n7399, n_6281, n_6282);
  and g13334 (n7400, \b[16] , n3638);
  and g13335 (n7401, \b[14] , n3843);
  and g13336 (n7402, \b[15] , n3633);
  and g13342 (n7405, n1237, n3641);
  not g13345 (n_6287, n7406);
  and g13346 (n7407, \a[32] , n_6287);
  not g13347 (n_6288, n7407);
  and g13348 (n7408, \a[32] , n_6288);
  and g13349 (n7409, n_6287, n_6288);
  not g13350 (n_6289, n7408);
  not g13351 (n_6290, n7409);
  and g13352 (n7410, n_6289, n_6290);
  and g13353 (n7411, n_6097, n_6102);
  and g13354 (n7412, n_6091, n_6094);
  and g13355 (n7413, \b[7] , n5777);
  and g13356 (n7414, \b[5] , n6059);
  and g13357 (n7415, \b[6] , n5772);
  and g13363 (n7418, n484, n5780);
  not g13366 (n_6295, n7419);
  and g13367 (n7420, \a[41] , n_6295);
  not g13368 (n_6296, n7420);
  and g13369 (n7421, \a[41] , n_6296);
  and g13370 (n7422, n_6295, n_6296);
  not g13371 (n_6297, n7421);
  not g13372 (n_6298, n7422);
  and g13373 (n7423, n_6297, n_6298);
  and g13374 (n7424, n6914, n7153);
  not g13375 (n_6299, n7424);
  and g13376 (n7425, n_6070, n_6299);
  and g13377 (n7426, \b[4] , n6595);
  and g13378 (n7427, \b[2] , n6902);
  and g13379 (n7428, \b[3] , n6590);
  and g13385 (n7431, n346, n6598);
  not g13388 (n_6304, n7432);
  and g13389 (n7433, \a[44] , n_6304);
  not g13390 (n_6305, n7433);
  and g13391 (n7434, \a[44] , n_6305);
  and g13392 (n7435, n_6304, n_6305);
  not g13393 (n_6306, n7434);
  not g13394 (n_6307, n7435);
  and g13395 (n7436, n_6306, n_6307);
  and g13396 (n7437, \a[47] , n_6057);
  and g13397 (n7438, n_6053, \a[46] );
  not g13398 (n_6310, \a[46] );
  and g13399 (n7439, \a[45] , n_6310);
  not g13400 (n_6311, n7438);
  not g13401 (n_6312, n7439);
  and g13402 (n7440, n_6311, n_6312);
  not g13403 (n_6313, n7440);
  and g13404 (n7441, n7152, n_6313);
  and g13405 (n7442, \b[0] , n7441);
  and g13406 (n7443, n_6310, \a[47] );
  not g13407 (n_6314, \a[47] );
  and g13408 (n7444, \a[46] , n_6314);
  not g13409 (n_6315, n7443);
  not g13410 (n_6316, n7444);
  and g13411 (n7445, n_6315, n_6316);
  and g13412 (n7446, n_6056, n7445);
  and g13413 (n7447, \b[1] , n7446);
  not g13414 (n_6317, n7442);
  not g13415 (n_6318, n7447);
  and g13416 (n7448, n_6317, n_6318);
  not g13417 (n_6319, n7445);
  and g13418 (n7449, n_6056, n_6319);
  and g13419 (n7450, n_21, n7449);
  not g13420 (n_6320, n7450);
  and g13421 (n7451, n7448, n_6320);
  not g13422 (n_6321, n7451);
  and g13423 (n7452, \a[47] , n_6321);
  not g13424 (n_6322, n7452);
  and g13425 (n7453, \a[47] , n_6322);
  and g13426 (n7454, n_6321, n_6322);
  not g13427 (n_6323, n7453);
  not g13428 (n_6324, n7454);
  and g13429 (n7455, n_6323, n_6324);
  not g13430 (n_6325, n7455);
  and g13431 (n7456, n7437, n_6325);
  not g13432 (n_6326, n7437);
  and g13433 (n7457, n_6326, n7455);
  not g13434 (n_6327, n7456);
  not g13435 (n_6328, n7457);
  and g13436 (n7458, n_6327, n_6328);
  not g13437 (n_6329, n7458);
  and g13438 (n7459, n7436, n_6329);
  not g13439 (n_6330, n7436);
  and g13440 (n7460, n_6330, n7458);
  not g13441 (n_6331, n7459);
  not g13442 (n_6332, n7460);
  and g13443 (n7461, n_6331, n_6332);
  not g13444 (n_6333, n7425);
  and g13445 (n7462, n_6333, n7461);
  not g13446 (n_6334, n7461);
  and g13447 (n7463, n7425, n_6334);
  not g13448 (n_6335, n7462);
  not g13449 (n_6336, n7463);
  and g13450 (n7464, n_6335, n_6336);
  not g13451 (n_6337, n7423);
  and g13452 (n7465, n_6337, n7464);
  not g13453 (n_6338, n7465);
  and g13454 (n7466, n7464, n_6338);
  and g13455 (n7467, n_6337, n_6338);
  not g13456 (n_6339, n7466);
  not g13457 (n_6340, n7467);
  and g13458 (n7468, n_6339, n_6340);
  and g13459 (n7469, n_6073, n_6079);
  and g13460 (n7470, n7468, n7469);
  not g13461 (n_6341, n7468);
  not g13462 (n_6342, n7469);
  and g13463 (n7471, n_6341, n_6342);
  not g13464 (n_6343, n7470);
  not g13465 (n_6344, n7471);
  and g13466 (n7472, n_6343, n_6344);
  and g13467 (n7473, \b[10] , n5035);
  and g13468 (n7474, \b[8] , n5277);
  and g13469 (n7475, \b[9] , n5030);
  and g13475 (n7478, n738, n5038);
  not g13478 (n_6349, n7479);
  and g13479 (n7480, \a[38] , n_6349);
  not g13480 (n_6350, n7480);
  and g13481 (n7481, \a[38] , n_6350);
  and g13482 (n7482, n_6349, n_6350);
  not g13483 (n_6351, n7481);
  not g13484 (n_6352, n7482);
  and g13485 (n7483, n_6351, n_6352);
  not g13486 (n_6353, n7483);
  and g13487 (n7484, n7472, n_6353);
  not g13488 (n_6354, n7472);
  and g13489 (n7485, n_6354, n7483);
  not g13490 (n_6355, n7412);
  not g13491 (n_6356, n7485);
  and g13492 (n7486, n_6355, n_6356);
  not g13493 (n_6357, n7484);
  and g13494 (n7487, n_6357, n7486);
  not g13495 (n_6358, n7487);
  and g13496 (n7488, n_6355, n_6358);
  and g13497 (n7489, n_6357, n_6358);
  and g13498 (n7490, n_6356, n7489);
  not g13499 (n_6359, n7488);
  not g13500 (n_6360, n7490);
  and g13501 (n7491, n_6359, n_6360);
  and g13502 (n7492, \b[13] , n4287);
  and g13503 (n7493, \b[11] , n4532);
  and g13504 (n7494, \b[12] , n4282);
  and g13510 (n7497, n1008, n4290);
  not g13513 (n_6365, n7498);
  and g13514 (n7499, \a[35] , n_6365);
  not g13515 (n_6366, n7499);
  and g13516 (n7500, \a[35] , n_6366);
  and g13517 (n7501, n_6365, n_6366);
  not g13518 (n_6367, n7500);
  not g13519 (n_6368, n7501);
  and g13520 (n7502, n_6367, n_6368);
  and g13521 (n7503, n7491, n7502);
  not g13522 (n_6369, n7491);
  not g13523 (n_6370, n7502);
  and g13524 (n7504, n_6369, n_6370);
  not g13525 (n_6371, n7503);
  not g13526 (n_6372, n7504);
  and g13527 (n7505, n_6371, n_6372);
  not g13528 (n_6373, n7411);
  and g13529 (n7506, n_6373, n7505);
  not g13530 (n_6374, n7505);
  and g13531 (n7507, n7411, n_6374);
  not g13532 (n_6375, n7506);
  not g13533 (n_6376, n7507);
  and g13534 (n7508, n_6375, n_6376);
  not g13535 (n_6377, n7410);
  and g13536 (n7509, n_6377, n7508);
  not g13537 (n_6378, n7509);
  and g13538 (n7510, n7508, n_6378);
  and g13539 (n7511, n_6377, n_6378);
  not g13540 (n_6379, n7510);
  not g13541 (n_6380, n7511);
  and g13542 (n7512, n_6379, n_6380);
  and g13543 (n7513, n_6118, n_6119);
  not g13544 (n_6381, n7513);
  and g13545 (n7514, n_6115, n_6381);
  and g13546 (n7515, n7512, n7514);
  not g13547 (n_6382, n7512);
  not g13548 (n_6383, n7514);
  and g13549 (n7516, n_6382, n_6383);
  not g13550 (n_6384, n7515);
  not g13551 (n_6385, n7516);
  and g13552 (n7517, n_6384, n_6385);
  and g13553 (n7518, \b[19] , n3050);
  and g13554 (n7519, \b[17] , n3243);
  and g13555 (n7520, \b[18] , n3045);
  and g13561 (n7523, n1708, n3053);
  not g13564 (n_6390, n7524);
  and g13565 (n7525, \a[29] , n_6390);
  not g13566 (n_6391, n7525);
  and g13567 (n7526, \a[29] , n_6391);
  and g13568 (n7527, n_6390, n_6391);
  not g13569 (n_6392, n7526);
  not g13570 (n_6393, n7527);
  and g13571 (n7528, n_6392, n_6393);
  not g13572 (n_6394, n7528);
  and g13573 (n7529, n7517, n_6394);
  not g13574 (n_6395, n7529);
  and g13575 (n7530, n7517, n_6395);
  and g13576 (n7531, n_6394, n_6395);
  not g13577 (n_6396, n7530);
  not g13578 (n_6397, n7531);
  and g13579 (n7532, n_6396, n_6397);
  and g13580 (n7533, n_6132, n_6136);
  and g13581 (n7534, n7532, n7533);
  not g13582 (n_6398, n7532);
  not g13583 (n_6399, n7533);
  and g13584 (n7535, n_6398, n_6399);
  not g13585 (n_6400, n7534);
  not g13586 (n_6401, n7535);
  and g13587 (n7536, n_6400, n_6401);
  and g13588 (n7537, \b[22] , n2539);
  and g13589 (n7538, \b[20] , n2685);
  and g13590 (n7539, \b[21] , n2534);
  and g13596 (n7542, n2145, n2542);
  not g13599 (n_6406, n7543);
  and g13600 (n7544, \a[26] , n_6406);
  not g13601 (n_6407, n7544);
  and g13602 (n7545, \a[26] , n_6407);
  and g13603 (n7546, n_6406, n_6407);
  not g13604 (n_6408, n7545);
  not g13605 (n_6409, n7546);
  and g13606 (n7547, n_6408, n_6409);
  not g13607 (n_6410, n7547);
  and g13608 (n7548, n7536, n_6410);
  not g13609 (n_6411, n7548);
  and g13610 (n7549, n7536, n_6411);
  and g13611 (n7550, n_6410, n_6411);
  not g13612 (n_6412, n7549);
  not g13613 (n_6413, n7550);
  and g13614 (n7551, n_6412, n_6413);
  and g13615 (n7552, n_6139, n_6145);
  and g13616 (n7553, n7551, n7552);
  not g13617 (n_6414, n7551);
  not g13618 (n_6415, n7552);
  and g13619 (n7554, n_6414, n_6415);
  not g13620 (n_6416, n7553);
  not g13621 (n_6417, n7554);
  and g13622 (n7555, n_6416, n_6417);
  and g13623 (n7556, \b[25] , n2048);
  and g13624 (n7557, \b[23] , n2198);
  and g13625 (n7558, \b[24] , n2043);
  and g13631 (n7561, n2051, n2485);
  not g13634 (n_6422, n7562);
  and g13635 (n7563, \a[23] , n_6422);
  not g13636 (n_6423, n7563);
  and g13637 (n7564, \a[23] , n_6423);
  and g13638 (n7565, n_6422, n_6423);
  not g13639 (n_6424, n7564);
  not g13640 (n_6425, n7565);
  and g13641 (n7566, n_6424, n_6425);
  not g13642 (n_6426, n7566);
  and g13643 (n7567, n7555, n_6426);
  not g13644 (n_6427, n7567);
  and g13645 (n7568, n7555, n_6427);
  and g13646 (n7569, n_6426, n_6427);
  not g13647 (n_6428, n7568);
  not g13648 (n_6429, n7569);
  and g13649 (n7570, n_6428, n_6429);
  and g13650 (n7571, n_6157, n_6160);
  not g13651 (n_6430, n7570);
  not g13652 (n_6431, n7571);
  and g13653 (n7572, n_6430, n_6431);
  and g13654 (n7573, n7570, n7571);
  not g13655 (n_6432, n7572);
  not g13656 (n_6433, n7573);
  and g13657 (n7574, n_6432, n_6433);
  not g13658 (n_6434, n7399);
  and g13659 (n7575, n_6434, n7574);
  not g13660 (n_6435, n7575);
  and g13661 (n7576, n_6434, n_6435);
  and g13662 (n7577, n7574, n_6435);
  not g13663 (n_6436, n7576);
  not g13664 (n_6437, n7577);
  and g13665 (n7578, n_6436, n_6437);
  not g13666 (n_6438, n7388);
  not g13667 (n_6439, n7578);
  and g13668 (n7579, n_6438, n_6439);
  not g13669 (n_6440, n7579);
  and g13670 (n7580, n_6438, n_6440);
  and g13671 (n7581, n_6439, n_6440);
  not g13672 (n_6441, n7580);
  not g13673 (n_6442, n7581);
  and g13674 (n7582, n_6441, n_6442);
  and g13675 (n7583, \b[31] , n1302);
  and g13676 (n7584, \b[29] , n1391);
  and g13677 (n7585, \b[30] , n1297);
  and g13683 (n7588, n1305, n3796);
  not g13686 (n_6447, n7589);
  and g13687 (n7590, \a[17] , n_6447);
  not g13688 (n_6448, n7590);
  and g13689 (n7591, \a[17] , n_6448);
  and g13690 (n7592, n_6447, n_6448);
  not g13691 (n_6449, n7591);
  not g13692 (n_6450, n7592);
  and g13693 (n7593, n_6449, n_6450);
  and g13694 (n7594, n7582, n7593);
  not g13695 (n_6451, n7582);
  not g13696 (n_6452, n7593);
  and g13697 (n7595, n_6451, n_6452);
  not g13698 (n_6453, n7594);
  not g13699 (n_6454, n7595);
  and g13700 (n7596, n_6453, n_6454);
  not g13701 (n_6455, n7386);
  and g13702 (n7597, n_6455, n7596);
  not g13703 (n_6456, n7596);
  and g13704 (n7598, n7386, n_6456);
  not g13705 (n_6457, n7597);
  not g13706 (n_6458, n7598);
  and g13707 (n7599, n_6457, n_6458);
  not g13708 (n_6459, n7385);
  and g13709 (n7600, n_6459, n7599);
  not g13710 (n_6460, n7600);
  and g13711 (n7601, n7599, n_6460);
  and g13712 (n7602, n_6459, n_6460);
  not g13713 (n_6461, n7601);
  not g13714 (n_6462, n7602);
  and g13715 (n7603, n_6461, n_6462);
  and g13716 (n7604, n_6190, n_6191);
  not g13717 (n_6463, n7604);
  and g13718 (n7605, n_6187, n_6463);
  and g13719 (n7606, n7603, n7605);
  not g13720 (n_6464, n7603);
  not g13721 (n_6465, n7605);
  and g13722 (n7607, n_6464, n_6465);
  not g13723 (n_6466, n7606);
  not g13724 (n_6467, n7607);
  and g13725 (n7608, n_6466, n_6467);
  and g13726 (n7609, \b[37] , n700);
  and g13727 (n7610, \b[35] , n767);
  and g13728 (n7611, \b[36] , n695);
  and g13734 (n7614, n703, n5181);
  not g13737 (n_6472, n7615);
  and g13738 (n7616, \a[11] , n_6472);
  not g13739 (n_6473, n7616);
  and g13740 (n7617, \a[11] , n_6473);
  and g13741 (n7618, n_6472, n_6473);
  not g13742 (n_6474, n7617);
  not g13743 (n_6475, n7618);
  and g13744 (n7619, n_6474, n_6475);
  not g13745 (n_6476, n7619);
  and g13746 (n7620, n7608, n_6476);
  not g13747 (n_6477, n7620);
  and g13748 (n7621, n7608, n_6477);
  and g13749 (n7622, n_6476, n_6477);
  not g13750 (n_6478, n7621);
  not g13751 (n_6479, n7622);
  and g13752 (n7623, n_6478, n_6479);
  and g13753 (n7624, n_6204, n_6209);
  and g13754 (n7625, n7623, n7624);
  not g13755 (n_6480, n7623);
  not g13756 (n_6481, n7624);
  and g13757 (n7626, n_6480, n_6481);
  not g13758 (n_6482, n7625);
  not g13759 (n_6483, n7626);
  and g13760 (n7627, n_6482, n_6483);
  and g13761 (n7628, \b[40] , n511);
  and g13762 (n7629, \b[38] , n541);
  and g13763 (n7630, \b[39] , n506);
  and g13769 (n7633, n514, n5955);
  not g13772 (n_6488, n7634);
  and g13773 (n7635, \a[8] , n_6488);
  not g13774 (n_6489, n7635);
  and g13775 (n7636, \a[8] , n_6489);
  and g13776 (n7637, n_6488, n_6489);
  not g13777 (n_6490, n7636);
  not g13778 (n_6491, n7637);
  and g13779 (n7638, n_6490, n_6491);
  not g13780 (n_6492, n7638);
  and g13781 (n7639, n7627, n_6492);
  not g13782 (n_6493, n7627);
  and g13783 (n7640, n_6493, n7638);
  not g13784 (n_6494, n7374);
  not g13785 (n_6495, n7640);
  and g13786 (n7641, n_6494, n_6495);
  not g13787 (n_6496, n7639);
  and g13788 (n7642, n_6496, n7641);
  not g13789 (n_6497, n7642);
  and g13790 (n7643, n_6494, n_6497);
  and g13791 (n7644, n_6496, n_6497);
  and g13792 (n7645, n_6495, n7644);
  not g13793 (n_6498, n7643);
  not g13794 (n_6499, n7645);
  and g13795 (n7646, n_6498, n_6499);
  and g13796 (n7647, \b[43] , n362);
  and g13797 (n7648, \b[41] , n403);
  and g13798 (n7649, \b[42] , n357);
  and g13804 (n7652, n365, n6515);
  not g13807 (n_6504, n7653);
  and g13808 (n7654, \a[5] , n_6504);
  not g13809 (n_6505, n7654);
  and g13810 (n7655, \a[5] , n_6505);
  and g13811 (n7656, n_6504, n_6505);
  not g13812 (n_6506, n7655);
  not g13813 (n_6507, n7656);
  and g13814 (n7657, n_6506, n_6507);
  not g13815 (n_6508, n7646);
  not g13816 (n_6509, n7657);
  and g13817 (n7658, n_6508, n_6509);
  not g13818 (n_6510, n7658);
  and g13819 (n7659, n_6508, n_6510);
  and g13820 (n7660, n_6509, n_6510);
  not g13821 (n_6511, n7659);
  not g13822 (n_6512, n7660);
  and g13823 (n7661, n_6511, n_6512);
  and g13824 (n7662, n_6235, n_6241);
  and g13825 (n7663, n7661, n7662);
  not g13826 (n_6513, n7661);
  not g13827 (n_6514, n7662);
  and g13828 (n7664, n_6513, n_6514);
  not g13829 (n_6515, n7663);
  not g13830 (n_6516, n7664);
  and g13831 (n7665, n_6515, n_6516);
  and g13832 (n7666, \b[46] , n266);
  and g13833 (n7667, \b[44] , n284);
  and g13834 (n7668, \b[45] , n261);
  and g13840 (n7671, n_6248, n_6251);
  not g13841 (n_6521, \b[46] );
  and g13842 (n7672, n_6246, n_6521);
  and g13843 (n7673, \b[45] , \b[46] );
  not g13844 (n_6522, n7672);
  not g13845 (n_6523, n7673);
  and g13846 (n7674, n_6522, n_6523);
  not g13847 (n_6524, n7671);
  and g13848 (n7675, n_6524, n7674);
  not g13849 (n_6525, n7674);
  and g13850 (n7676, n7671, n_6525);
  not g13851 (n_6526, n7675);
  not g13852 (n_6527, n7676);
  and g13853 (n7677, n_6526, n_6527);
  and g13854 (n7678, n269, n7677);
  not g13857 (n_6529, n7679);
  and g13858 (n7680, \a[2] , n_6529);
  not g13859 (n_6530, n7680);
  and g13860 (n7681, \a[2] , n_6530);
  and g13861 (n7682, n_6529, n_6530);
  not g13862 (n_6531, n7681);
  not g13863 (n_6532, n7682);
  and g13864 (n7683, n_6531, n_6532);
  not g13865 (n_6533, n7683);
  and g13866 (n7684, n7665, n_6533);
  not g13867 (n_6534, n7684);
  and g13868 (n7685, n7665, n_6534);
  and g13869 (n7686, n_6533, n_6534);
  not g13870 (n_6535, n7685);
  not g13871 (n_6536, n7686);
  and g13872 (n7687, n_6535, n_6536);
  and g13873 (n7688, n_6261, n_6264);
  not g13874 (n_6537, n7687);
  not g13875 (n_6538, n7688);
  and g13876 (n7689, n_6537, n_6538);
  and g13877 (n7690, n7687, n7688);
  not g13878 (n_6539, n7689);
  not g13879 (n_6540, n7690);
  and g13880 (\f[46] , n_6539, n_6540);
  and g13881 (n7692, \b[47] , n266);
  and g13882 (n7693, \b[45] , n284);
  and g13883 (n7694, \b[46] , n261);
  and g13889 (n7697, n_6523, n_6526);
  not g13890 (n_6545, \b[47] );
  and g13891 (n7698, n_6521, n_6545);
  and g13892 (n7699, \b[46] , \b[47] );
  not g13893 (n_6546, n7698);
  not g13894 (n_6547, n7699);
  and g13895 (n7700, n_6546, n_6547);
  not g13896 (n_6548, n7697);
  and g13897 (n7701, n_6548, n7700);
  not g13898 (n_6549, n7700);
  and g13899 (n7702, n7697, n_6549);
  not g13900 (n_6550, n7701);
  not g13901 (n_6551, n7702);
  and g13902 (n7703, n_6550, n_6551);
  and g13903 (n7704, n269, n7703);
  not g13906 (n_6553, n7705);
  and g13907 (n7706, \a[2] , n_6553);
  not g13908 (n_6554, n7706);
  and g13909 (n7707, \a[2] , n_6554);
  and g13910 (n7708, n_6553, n_6554);
  not g13911 (n_6555, n7707);
  not g13912 (n_6556, n7708);
  and g13913 (n7709, n_6555, n_6556);
  and g13914 (n7710, n_6510, n_6516);
  and g13915 (n7711, \b[35] , n951);
  and g13916 (n7712, \b[33] , n1056);
  and g13917 (n7713, \b[34] , n946);
  and g13923 (n7716, n954, n4696);
  not g13926 (n_6561, n7717);
  and g13927 (n7718, \a[14] , n_6561);
  not g13928 (n_6562, n7718);
  and g13929 (n7719, \a[14] , n_6562);
  and g13930 (n7720, n_6561, n_6562);
  not g13931 (n_6563, n7719);
  not g13932 (n_6564, n7720);
  and g13933 (n7721, n_6563, n_6564);
  and g13934 (n7722, n_6454, n_6457);
  and g13935 (n7723, \b[32] , n1302);
  and g13936 (n7724, \b[30] , n1391);
  and g13937 (n7725, \b[31] , n1297);
  and g13943 (n7728, n1305, n4013);
  not g13946 (n_6569, n7729);
  and g13947 (n7730, \a[17] , n_6569);
  not g13948 (n_6570, n7730);
  and g13949 (n7731, \a[17] , n_6570);
  and g13950 (n7732, n_6569, n_6570);
  not g13951 (n_6571, n7731);
  not g13952 (n_6572, n7732);
  and g13953 (n7733, n_6571, n_6572);
  and g13954 (n7734, n_6435, n_6440);
  and g13955 (n7735, \b[29] , n1627);
  and g13956 (n7736, \b[27] , n1763);
  and g13957 (n7737, \b[28] , n1622);
  and g13963 (n7740, n1630, n3383);
  not g13966 (n_6577, n7741);
  and g13967 (n7742, \a[20] , n_6577);
  not g13968 (n_6578, n7742);
  and g13969 (n7743, \a[20] , n_6578);
  and g13970 (n7744, n_6577, n_6578);
  not g13971 (n_6579, n7743);
  not g13972 (n_6580, n7744);
  and g13973 (n7745, n_6579, n_6580);
  and g13974 (n7746, n_6427, n_6432);
  and g13975 (n7747, n_6411, n_6417);
  and g13976 (n7748, n_6378, n_6385);
  and g13977 (n7749, \b[17] , n3638);
  and g13978 (n7750, \b[15] , n3843);
  and g13979 (n7751, \b[16] , n3633);
  and g13985 (n7754, n1356, n3641);
  not g13988 (n_6585, n7755);
  and g13989 (n7756, \a[32] , n_6585);
  not g13990 (n_6586, n7756);
  and g13991 (n7757, \a[32] , n_6586);
  and g13992 (n7758, n_6585, n_6586);
  not g13993 (n_6587, n7757);
  not g13994 (n_6588, n7758);
  and g13995 (n7759, n_6587, n_6588);
  and g13996 (n7760, n_6372, n_6375);
  and g13997 (n7761, \b[14] , n4287);
  and g13998 (n7762, \b[12] , n4532);
  and g13999 (n7763, \b[13] , n4282);
  and g14005 (n7766, n1034, n4290);
  not g14008 (n_6593, n7767);
  and g14009 (n7768, \a[35] , n_6593);
  not g14010 (n_6594, n7768);
  and g14011 (n7769, \a[35] , n_6594);
  and g14012 (n7770, n_6593, n_6594);
  not g14013 (n_6595, n7769);
  not g14014 (n_6596, n7770);
  and g14015 (n7771, n_6595, n_6596);
  and g14016 (n7772, n_6338, n_6344);
  and g14017 (n7773, \b[8] , n5777);
  and g14018 (n7774, \b[6] , n6059);
  and g14019 (n7775, \b[7] , n5772);
  and g14025 (n7778, n585, n5780);
  not g14028 (n_6601, n7779);
  and g14029 (n7780, \a[41] , n_6601);
  not g14030 (n_6602, n7780);
  and g14031 (n7781, \a[41] , n_6602);
  and g14032 (n7782, n_6601, n_6602);
  not g14033 (n_6603, n7781);
  not g14034 (n_6604, n7782);
  and g14035 (n7783, n_6603, n_6604);
  and g14036 (n7784, n_6332, n_6335);
  and g14037 (n7785, \b[2] , n7446);
  and g14038 (n7786, n7152, n_6319);
  and g14039 (n7787, n7440, n7786);
  and g14040 (n7788, \b[0] , n7787);
  and g14041 (n7789, \b[1] , n7441);
  and g14047 (n7792, n296, n7449);
  not g14050 (n_6609, n7793);
  and g14051 (n7794, \a[47] , n_6609);
  not g14052 (n_6610, n7794);
  and g14053 (n7795, \a[47] , n_6610);
  and g14054 (n7796, n_6609, n_6610);
  not g14055 (n_6611, n7795);
  not g14056 (n_6612, n7796);
  and g14057 (n7797, n_6611, n_6612);
  and g14058 (n7798, n_6327, n7797);
  not g14059 (n_6613, n7797);
  and g14060 (n7799, n7456, n_6613);
  not g14061 (n_6614, n7798);
  not g14062 (n_6615, n7799);
  and g14063 (n7800, n_6614, n_6615);
  and g14064 (n7801, \b[5] , n6595);
  and g14065 (n7802, \b[3] , n6902);
  and g14066 (n7803, \b[4] , n6590);
  and g14072 (n7806, n394, n6598);
  not g14075 (n_6620, n7807);
  and g14076 (n7808, \a[44] , n_6620);
  not g14077 (n_6621, n7808);
  and g14078 (n7809, \a[44] , n_6621);
  and g14079 (n7810, n_6620, n_6621);
  not g14080 (n_6622, n7809);
  not g14081 (n_6623, n7810);
  and g14082 (n7811, n_6622, n_6623);
  not g14083 (n_6624, n7811);
  and g14084 (n7812, n7800, n_6624);
  not g14085 (n_6625, n7812);
  and g14086 (n7813, n7800, n_6625);
  and g14087 (n7814, n_6624, n_6625);
  not g14088 (n_6626, n7813);
  not g14089 (n_6627, n7814);
  and g14090 (n7815, n_6626, n_6627);
  not g14091 (n_6628, n7784);
  not g14092 (n_6629, n7815);
  and g14093 (n7816, n_6628, n_6629);
  and g14094 (n7817, n7784, n7815);
  not g14095 (n_6630, n7816);
  not g14096 (n_6631, n7817);
  and g14097 (n7818, n_6630, n_6631);
  not g14098 (n_6632, n7783);
  and g14099 (n7819, n_6632, n7818);
  not g14100 (n_6633, n7819);
  and g14101 (n7820, n_6632, n_6633);
  and g14102 (n7821, n7818, n_6633);
  not g14103 (n_6634, n7820);
  not g14104 (n_6635, n7821);
  and g14105 (n7822, n_6634, n_6635);
  not g14106 (n_6636, n7772);
  not g14107 (n_6637, n7822);
  and g14108 (n7823, n_6636, n_6637);
  not g14109 (n_6638, n7823);
  and g14110 (n7824, n_6636, n_6638);
  and g14111 (n7825, n_6637, n_6638);
  not g14112 (n_6639, n7824);
  not g14113 (n_6640, n7825);
  and g14114 (n7826, n_6639, n_6640);
  and g14115 (n7827, \b[11] , n5035);
  and g14116 (n7828, \b[9] , n5277);
  and g14117 (n7829, \b[10] , n5030);
  and g14123 (n7832, n818, n5038);
  not g14126 (n_6645, n7833);
  and g14127 (n7834, \a[38] , n_6645);
  not g14128 (n_6646, n7834);
  and g14129 (n7835, \a[38] , n_6646);
  and g14130 (n7836, n_6645, n_6646);
  not g14131 (n_6647, n7835);
  not g14132 (n_6648, n7836);
  and g14133 (n7837, n_6647, n_6648);
  and g14134 (n7838, n7826, n7837);
  not g14135 (n_6649, n7826);
  not g14136 (n_6650, n7837);
  and g14137 (n7839, n_6649, n_6650);
  not g14138 (n_6651, n7838);
  not g14139 (n_6652, n7839);
  and g14140 (n7840, n_6651, n_6652);
  not g14141 (n_6653, n7489);
  and g14142 (n7841, n_6653, n7840);
  not g14143 (n_6654, n7840);
  and g14144 (n7842, n7489, n_6654);
  not g14145 (n_6655, n7841);
  not g14146 (n_6656, n7842);
  and g14147 (n7843, n_6655, n_6656);
  not g14148 (n_6657, n7771);
  and g14149 (n7844, n_6657, n7843);
  not g14150 (n_6658, n7844);
  and g14151 (n7845, n7843, n_6658);
  and g14152 (n7846, n_6657, n_6658);
  not g14153 (n_6659, n7845);
  not g14154 (n_6660, n7846);
  and g14155 (n7847, n_6659, n_6660);
  not g14156 (n_6661, n7760);
  not g14157 (n_6662, n7847);
  and g14158 (n7848, n_6661, n_6662);
  and g14159 (n7849, n7760, n7847);
  not g14160 (n_6663, n7848);
  not g14161 (n_6664, n7849);
  and g14162 (n7850, n_6663, n_6664);
  not g14163 (n_6665, n7759);
  and g14164 (n7851, n_6665, n7850);
  not g14165 (n_6666, n7851);
  and g14166 (n7852, n_6665, n_6666);
  and g14167 (n7853, n7850, n_6666);
  not g14168 (n_6667, n7852);
  not g14169 (n_6668, n7853);
  and g14170 (n7854, n_6667, n_6668);
  not g14171 (n_6669, n7748);
  not g14172 (n_6670, n7854);
  and g14173 (n7855, n_6669, n_6670);
  not g14174 (n_6671, n7855);
  and g14175 (n7856, n_6669, n_6671);
  and g14176 (n7857, n_6670, n_6671);
  not g14177 (n_6672, n7856);
  not g14178 (n_6673, n7857);
  and g14179 (n7858, n_6672, n_6673);
  and g14180 (n7859, \b[20] , n3050);
  and g14181 (n7860, \b[18] , n3243);
  and g14182 (n7861, \b[19] , n3045);
  and g14188 (n7864, n1846, n3053);
  not g14191 (n_6678, n7865);
  and g14192 (n7866, \a[29] , n_6678);
  not g14193 (n_6679, n7866);
  and g14194 (n7867, \a[29] , n_6679);
  and g14195 (n7868, n_6678, n_6679);
  not g14196 (n_6680, n7867);
  not g14197 (n_6681, n7868);
  and g14198 (n7869, n_6680, n_6681);
  not g14199 (n_6682, n7858);
  not g14200 (n_6683, n7869);
  and g14201 (n7870, n_6682, n_6683);
  not g14202 (n_6684, n7870);
  and g14203 (n7871, n_6682, n_6684);
  and g14204 (n7872, n_6683, n_6684);
  not g14205 (n_6685, n7871);
  not g14206 (n_6686, n7872);
  and g14207 (n7873, n_6685, n_6686);
  and g14208 (n7874, n_6395, n_6401);
  and g14209 (n7875, n7873, n7874);
  not g14210 (n_6687, n7873);
  not g14211 (n_6688, n7874);
  and g14212 (n7876, n_6687, n_6688);
  not g14213 (n_6689, n7875);
  not g14214 (n_6690, n7876);
  and g14215 (n7877, n_6689, n_6690);
  and g14216 (n7878, \b[23] , n2539);
  and g14217 (n7879, \b[21] , n2685);
  and g14218 (n7880, \b[22] , n2534);
  and g14224 (n7883, n2300, n2542);
  not g14227 (n_6695, n7884);
  and g14228 (n7885, \a[26] , n_6695);
  not g14229 (n_6696, n7885);
  and g14230 (n7886, \a[26] , n_6696);
  and g14231 (n7887, n_6695, n_6696);
  not g14232 (n_6697, n7886);
  not g14233 (n_6698, n7887);
  and g14234 (n7888, n_6697, n_6698);
  not g14235 (n_6699, n7888);
  and g14236 (n7889, n7877, n_6699);
  not g14237 (n_6700, n7877);
  and g14238 (n7890, n_6700, n7888);
  not g14239 (n_6701, n7747);
  not g14240 (n_6702, n7890);
  and g14241 (n7891, n_6701, n_6702);
  not g14242 (n_6703, n7889);
  and g14243 (n7892, n_6703, n7891);
  not g14244 (n_6704, n7892);
  and g14245 (n7893, n_6701, n_6704);
  and g14246 (n7894, n_6703, n_6704);
  and g14247 (n7895, n_6702, n7894);
  not g14248 (n_6705, n7893);
  not g14249 (n_6706, n7895);
  and g14250 (n7896, n_6705, n_6706);
  and g14251 (n7897, \b[26] , n2048);
  and g14252 (n7898, \b[24] , n2198);
  and g14253 (n7899, \b[25] , n2043);
  and g14259 (n7902, n2051, n2813);
  not g14262 (n_6711, n7903);
  and g14263 (n7904, \a[23] , n_6711);
  not g14264 (n_6712, n7904);
  and g14265 (n7905, \a[23] , n_6712);
  and g14266 (n7906, n_6711, n_6712);
  not g14267 (n_6713, n7905);
  not g14268 (n_6714, n7906);
  and g14269 (n7907, n_6713, n_6714);
  and g14270 (n7908, n7896, n7907);
  not g14271 (n_6715, n7896);
  not g14272 (n_6716, n7907);
  and g14273 (n7909, n_6715, n_6716);
  not g14274 (n_6717, n7908);
  not g14275 (n_6718, n7909);
  and g14276 (n7910, n_6717, n_6718);
  not g14277 (n_6719, n7746);
  and g14278 (n7911, n_6719, n7910);
  not g14279 (n_6720, n7910);
  and g14280 (n7912, n7746, n_6720);
  not g14281 (n_6721, n7911);
  not g14282 (n_6722, n7912);
  and g14283 (n7913, n_6721, n_6722);
  not g14284 (n_6723, n7913);
  and g14285 (n7914, n7745, n_6723);
  not g14286 (n_6724, n7745);
  and g14287 (n7915, n_6724, n7913);
  not g14288 (n_6725, n7914);
  not g14289 (n_6726, n7915);
  and g14290 (n7916, n_6725, n_6726);
  not g14291 (n_6727, n7734);
  and g14292 (n7917, n_6727, n7916);
  not g14293 (n_6728, n7916);
  and g14294 (n7918, n7734, n_6728);
  not g14295 (n_6729, n7917);
  not g14296 (n_6730, n7918);
  and g14297 (n7919, n_6729, n_6730);
  not g14298 (n_6731, n7919);
  and g14299 (n7920, n7733, n_6731);
  not g14300 (n_6732, n7733);
  and g14301 (n7921, n_6732, n7919);
  not g14302 (n_6733, n7920);
  not g14303 (n_6734, n7921);
  and g14304 (n7922, n_6733, n_6734);
  not g14305 (n_6735, n7722);
  and g14306 (n7923, n_6735, n7922);
  not g14307 (n_6736, n7922);
  and g14308 (n7924, n7722, n_6736);
  not g14309 (n_6737, n7923);
  not g14310 (n_6738, n7924);
  and g14311 (n7925, n_6737, n_6738);
  not g14312 (n_6739, n7721);
  and g14313 (n7926, n_6739, n7925);
  not g14314 (n_6740, n7926);
  and g14315 (n7927, n7925, n_6740);
  and g14316 (n7928, n_6739, n_6740);
  not g14317 (n_6741, n7927);
  not g14318 (n_6742, n7928);
  and g14319 (n7929, n_6741, n_6742);
  and g14320 (n7930, n_6460, n_6467);
  and g14321 (n7931, n7929, n7930);
  not g14322 (n_6743, n7929);
  not g14323 (n_6744, n7930);
  and g14324 (n7932, n_6743, n_6744);
  not g14325 (n_6745, n7931);
  not g14326 (n_6746, n7932);
  and g14327 (n7933, n_6745, n_6746);
  and g14328 (n7934, \b[38] , n700);
  and g14329 (n7935, \b[36] , n767);
  and g14330 (n7936, \b[37] , n695);
  and g14336 (n7939, n703, n5205);
  not g14339 (n_6751, n7940);
  and g14340 (n7941, \a[11] , n_6751);
  not g14341 (n_6752, n7941);
  and g14342 (n7942, \a[11] , n_6752);
  and g14343 (n7943, n_6751, n_6752);
  not g14344 (n_6753, n7942);
  not g14345 (n_6754, n7943);
  and g14346 (n7944, n_6753, n_6754);
  not g14347 (n_6755, n7944);
  and g14348 (n7945, n7933, n_6755);
  not g14349 (n_6756, n7945);
  and g14350 (n7946, n7933, n_6756);
  and g14351 (n7947, n_6755, n_6756);
  not g14352 (n_6757, n7946);
  not g14353 (n_6758, n7947);
  and g14354 (n7948, n_6757, n_6758);
  and g14355 (n7949, n_6477, n_6483);
  and g14356 (n7950, n7948, n7949);
  not g14357 (n_6759, n7948);
  not g14358 (n_6760, n7949);
  and g14359 (n7951, n_6759, n_6760);
  not g14360 (n_6761, n7950);
  not g14361 (n_6762, n7951);
  and g14362 (n7952, n_6761, n_6762);
  and g14363 (n7953, \b[41] , n511);
  and g14364 (n7954, \b[39] , n541);
  and g14365 (n7955, \b[40] , n506);
  and g14371 (n7958, n514, n6219);
  not g14374 (n_6767, n7959);
  and g14375 (n7960, \a[8] , n_6767);
  not g14376 (n_6768, n7960);
  and g14377 (n7961, \a[8] , n_6768);
  and g14378 (n7962, n_6767, n_6768);
  not g14379 (n_6769, n7961);
  not g14380 (n_6770, n7962);
  and g14381 (n7963, n_6769, n_6770);
  not g14382 (n_6771, n7963);
  and g14383 (n7964, n7952, n_6771);
  not g14384 (n_6772, n7952);
  and g14385 (n7965, n_6772, n7963);
  not g14386 (n_6773, n7644);
  not g14387 (n_6774, n7965);
  and g14388 (n7966, n_6773, n_6774);
  not g14389 (n_6775, n7964);
  and g14390 (n7967, n_6775, n7966);
  not g14391 (n_6776, n7967);
  and g14392 (n7968, n_6773, n_6776);
  and g14393 (n7969, n_6775, n_6776);
  and g14394 (n7970, n_6774, n7969);
  not g14395 (n_6777, n7968);
  not g14396 (n_6778, n7970);
  and g14397 (n7971, n_6777, n_6778);
  and g14398 (n7972, \b[44] , n362);
  and g14399 (n7973, \b[42] , n403);
  and g14400 (n7974, \b[43] , n357);
  and g14406 (n7977, n365, n7072);
  not g14409 (n_6783, n7978);
  and g14410 (n7979, \a[5] , n_6783);
  not g14411 (n_6784, n7979);
  and g14412 (n7980, \a[5] , n_6784);
  and g14413 (n7981, n_6783, n_6784);
  not g14414 (n_6785, n7980);
  not g14415 (n_6786, n7981);
  and g14416 (n7982, n_6785, n_6786);
  and g14417 (n7983, n7971, n7982);
  not g14418 (n_6787, n7971);
  not g14419 (n_6788, n7982);
  and g14420 (n7984, n_6787, n_6788);
  not g14421 (n_6789, n7983);
  not g14422 (n_6790, n7984);
  and g14423 (n7985, n_6789, n_6790);
  not g14424 (n_6791, n7710);
  and g14425 (n7986, n_6791, n7985);
  not g14426 (n_6792, n7985);
  and g14427 (n7987, n7710, n_6792);
  not g14428 (n_6793, n7986);
  not g14429 (n_6794, n7987);
  and g14430 (n7988, n_6793, n_6794);
  not g14431 (n_6795, n7709);
  and g14432 (n7989, n_6795, n7988);
  not g14433 (n_6796, n7989);
  and g14434 (n7990, n7988, n_6796);
  and g14435 (n7991, n_6795, n_6796);
  not g14436 (n_6797, n7990);
  not g14437 (n_6798, n7991);
  and g14438 (n7992, n_6797, n_6798);
  and g14439 (n7993, n_6534, n_6539);
  not g14440 (n_6799, n7992);
  not g14441 (n_6800, n7993);
  and g14442 (n7994, n_6799, n_6800);
  and g14443 (n7995, n7992, n7993);
  not g14444 (n_6801, n7994);
  not g14445 (n_6802, n7995);
  and g14446 (\f[47] , n_6801, n_6802);
  and g14447 (n7997, n_6796, n_6801);
  and g14448 (n7998, \b[48] , n266);
  and g14449 (n7999, \b[46] , n284);
  and g14450 (n8000, \b[47] , n261);
  and g14456 (n8003, n_6547, n_6550);
  not g14457 (n_6807, \b[48] );
  and g14458 (n8004, n_6545, n_6807);
  and g14459 (n8005, \b[47] , \b[48] );
  not g14460 (n_6808, n8004);
  not g14461 (n_6809, n8005);
  and g14462 (n8006, n_6808, n_6809);
  not g14463 (n_6810, n8003);
  and g14464 (n8007, n_6810, n8006);
  not g14465 (n_6811, n8006);
  and g14466 (n8008, n8003, n_6811);
  not g14467 (n_6812, n8007);
  not g14468 (n_6813, n8008);
  and g14469 (n8009, n_6812, n_6813);
  and g14470 (n8010, n269, n8009);
  not g14473 (n_6815, n8011);
  and g14474 (n8012, \a[2] , n_6815);
  not g14475 (n_6816, n8012);
  and g14476 (n8013, \a[2] , n_6816);
  and g14477 (n8014, n_6815, n_6816);
  not g14478 (n_6817, n8013);
  not g14479 (n_6818, n8014);
  and g14480 (n8015, n_6817, n_6818);
  and g14481 (n8016, n_6790, n_6793);
  and g14482 (n8017, n_6740, n_6746);
  and g14483 (n8018, n_6734, n_6737);
  and g14484 (n8019, \b[33] , n1302);
  and g14485 (n8020, \b[31] , n1391);
  and g14486 (n8021, \b[32] , n1297);
  and g14492 (n8024, n1305, n4223);
  not g14495 (n_6823, n8025);
  and g14496 (n8026, \a[17] , n_6823);
  not g14497 (n_6824, n8026);
  and g14498 (n8027, \a[17] , n_6824);
  and g14499 (n8028, n_6823, n_6824);
  not g14500 (n_6825, n8027);
  not g14501 (n_6826, n8028);
  and g14502 (n8029, n_6825, n_6826);
  and g14503 (n8030, n_6726, n_6729);
  and g14504 (n8031, n_6718, n_6721);
  and g14505 (n8032, \b[27] , n2048);
  and g14506 (n8033, \b[25] , n2198);
  and g14507 (n8034, \b[26] , n2043);
  and g14513 (n8037, n2051, n2990);
  not g14516 (n_6831, n8038);
  and g14517 (n8039, \a[23] , n_6831);
  not g14518 (n_6832, n8039);
  and g14519 (n8040, \a[23] , n_6832);
  and g14520 (n8041, n_6831, n_6832);
  not g14521 (n_6833, n8040);
  not g14522 (n_6834, n8041);
  and g14523 (n8042, n_6833, n_6834);
  and g14524 (n8043, n_6658, n_6663);
  and g14525 (n8044, \b[15] , n4287);
  and g14526 (n8045, \b[13] , n4532);
  and g14527 (n8046, \b[14] , n4282);
  and g14533 (n8049, n1131, n4290);
  not g14536 (n_6839, n8050);
  and g14537 (n8051, \a[35] , n_6839);
  not g14538 (n_6840, n8051);
  and g14539 (n8052, \a[35] , n_6840);
  and g14540 (n8053, n_6839, n_6840);
  not g14541 (n_6841, n8052);
  not g14542 (n_6842, n8053);
  and g14543 (n8054, n_6841, n_6842);
  and g14544 (n8055, n_6652, n_6655);
  and g14545 (n8056, \b[12] , n5035);
  and g14546 (n8057, \b[10] , n5277);
  and g14547 (n8058, \b[11] , n5030);
  and g14553 (n8061, n842, n5038);
  not g14556 (n_6847, n8062);
  and g14557 (n8063, \a[38] , n_6847);
  not g14558 (n_6848, n8063);
  and g14559 (n8064, \a[38] , n_6848);
  and g14560 (n8065, n_6847, n_6848);
  not g14561 (n_6849, n8064);
  not g14562 (n_6850, n8065);
  and g14563 (n8066, n_6849, n_6850);
  and g14564 (n8067, n_6633, n_6638);
  and g14565 (n8068, \b[6] , n6595);
  and g14566 (n8069, \b[4] , n6902);
  and g14567 (n8070, \b[5] , n6590);
  and g14573 (n8073, n459, n6598);
  not g14576 (n_6855, n8074);
  and g14577 (n8075, \a[44] , n_6855);
  not g14578 (n_6856, n8075);
  and g14579 (n8076, \a[44] , n_6856);
  and g14580 (n8077, n_6855, n_6856);
  not g14581 (n_6857, n8076);
  not g14582 (n_6858, n8077);
  and g14583 (n8078, n_6857, n_6858);
  not g14584 (n_6860, \a[48] );
  and g14585 (n8079, \a[47] , n_6860);
  and g14586 (n8080, n_6314, \a[48] );
  not g14587 (n_6861, n8079);
  not g14588 (n_6862, n8080);
  and g14589 (n8081, n_6861, n_6862);
  not g14590 (n_6863, n8081);
  and g14591 (n8082, \b[0] , n_6863);
  and g14592 (n8083, n_6615, n8082);
  not g14593 (n_6864, n8082);
  and g14594 (n8084, n7799, n_6864);
  not g14595 (n_6865, n8083);
  not g14596 (n_6866, n8084);
  and g14597 (n8085, n_6865, n_6866);
  and g14598 (n8086, \b[3] , n7446);
  and g14599 (n8087, \b[1] , n7787);
  and g14600 (n8088, \b[2] , n7441);
  and g14606 (n8091, n318, n7449);
  not g14609 (n_6871, n8092);
  and g14610 (n8093, \a[47] , n_6871);
  not g14611 (n_6872, n8093);
  and g14612 (n8094, \a[47] , n_6872);
  and g14613 (n8095, n_6871, n_6872);
  not g14614 (n_6873, n8094);
  not g14615 (n_6874, n8095);
  and g14616 (n8096, n_6873, n_6874);
  not g14617 (n_6875, n8085);
  not g14618 (n_6876, n8096);
  and g14619 (n8097, n_6875, n_6876);
  and g14620 (n8098, n8085, n8096);
  not g14621 (n_6877, n8097);
  not g14622 (n_6878, n8098);
  and g14623 (n8099, n_6877, n_6878);
  not g14624 (n_6879, n8078);
  and g14625 (n8100, n_6879, n8099);
  not g14626 (n_6880, n8100);
  and g14627 (n8101, n8099, n_6880);
  and g14628 (n8102, n_6879, n_6880);
  not g14629 (n_6881, n8101);
  not g14630 (n_6882, n8102);
  and g14631 (n8103, n_6881, n_6882);
  and g14632 (n8104, n_6625, n_6630);
  and g14633 (n8105, n8103, n8104);
  not g14634 (n_6883, n8103);
  not g14635 (n_6884, n8104);
  and g14636 (n8106, n_6883, n_6884);
  not g14637 (n_6885, n8105);
  not g14638 (n_6886, n8106);
  and g14639 (n8107, n_6885, n_6886);
  and g14640 (n8108, \b[9] , n5777);
  and g14641 (n8109, \b[7] , n6059);
  and g14642 (n8110, \b[8] , n5772);
  and g14648 (n8113, n651, n5780);
  not g14651 (n_6891, n8114);
  and g14652 (n8115, \a[41] , n_6891);
  not g14653 (n_6892, n8115);
  and g14654 (n8116, \a[41] , n_6892);
  and g14655 (n8117, n_6891, n_6892);
  not g14656 (n_6893, n8116);
  not g14657 (n_6894, n8117);
  and g14658 (n8118, n_6893, n_6894);
  not g14659 (n_6895, n8107);
  and g14660 (n8119, n_6895, n8118);
  not g14661 (n_6896, n8118);
  and g14662 (n8120, n8107, n_6896);
  not g14663 (n_6897, n8119);
  not g14664 (n_6898, n8120);
  and g14665 (n8121, n_6897, n_6898);
  not g14666 (n_6899, n8067);
  and g14667 (n8122, n_6899, n8121);
  not g14668 (n_6900, n8121);
  and g14669 (n8123, n8067, n_6900);
  not g14670 (n_6901, n8122);
  not g14671 (n_6902, n8123);
  and g14672 (n8124, n_6901, n_6902);
  not g14673 (n_6903, n8066);
  and g14674 (n8125, n_6903, n8124);
  not g14675 (n_6904, n8125);
  and g14676 (n8126, n_6903, n_6904);
  and g14677 (n8127, n8124, n_6904);
  not g14678 (n_6905, n8126);
  not g14679 (n_6906, n8127);
  and g14680 (n8128, n_6905, n_6906);
  not g14681 (n_6907, n8055);
  not g14682 (n_6908, n8128);
  and g14683 (n8129, n_6907, n_6908);
  and g14684 (n8130, n8055, n_6906);
  and g14685 (n8131, n_6905, n8130);
  not g14686 (n_6909, n8129);
  not g14687 (n_6910, n8131);
  and g14688 (n8132, n_6909, n_6910);
  not g14689 (n_6911, n8054);
  and g14690 (n8133, n_6911, n8132);
  not g14691 (n_6912, n8132);
  and g14692 (n8134, n8054, n_6912);
  not g14693 (n_6913, n8133);
  not g14694 (n_6914, n8134);
  and g14695 (n8135, n_6913, n_6914);
  not g14696 (n_6915, n8043);
  and g14697 (n8136, n_6915, n8135);
  not g14698 (n_6916, n8135);
  and g14699 (n8137, n8043, n_6916);
  not g14700 (n_6917, n8136);
  not g14701 (n_6918, n8137);
  and g14702 (n8138, n_6917, n_6918);
  and g14703 (n8139, \b[18] , n3638);
  and g14704 (n8140, \b[16] , n3843);
  and g14705 (n8141, \b[17] , n3633);
  and g14711 (n8144, n1566, n3641);
  not g14714 (n_6923, n8145);
  and g14715 (n8146, \a[32] , n_6923);
  not g14716 (n_6924, n8146);
  and g14717 (n8147, \a[32] , n_6924);
  and g14718 (n8148, n_6923, n_6924);
  not g14719 (n_6925, n8147);
  not g14720 (n_6926, n8148);
  and g14721 (n8149, n_6925, n_6926);
  not g14722 (n_6927, n8149);
  and g14723 (n8150, n8138, n_6927);
  not g14724 (n_6928, n8150);
  and g14725 (n8151, n8138, n_6928);
  and g14726 (n8152, n_6927, n_6928);
  not g14727 (n_6929, n8151);
  not g14728 (n_6930, n8152);
  and g14729 (n8153, n_6929, n_6930);
  and g14730 (n8154, n_6666, n_6671);
  and g14731 (n8155, n8153, n8154);
  not g14732 (n_6931, n8153);
  not g14733 (n_6932, n8154);
  and g14734 (n8156, n_6931, n_6932);
  not g14735 (n_6933, n8155);
  not g14736 (n_6934, n8156);
  and g14737 (n8157, n_6933, n_6934);
  and g14738 (n8158, \b[21] , n3050);
  and g14739 (n8159, \b[19] , n3243);
  and g14740 (n8160, \b[20] , n3045);
  and g14746 (n8163, n1984, n3053);
  not g14749 (n_6939, n8164);
  and g14750 (n8165, \a[29] , n_6939);
  not g14751 (n_6940, n8165);
  and g14752 (n8166, \a[29] , n_6940);
  and g14753 (n8167, n_6939, n_6940);
  not g14754 (n_6941, n8166);
  not g14755 (n_6942, n8167);
  and g14756 (n8168, n_6941, n_6942);
  not g14757 (n_6943, n8168);
  and g14758 (n8169, n8157, n_6943);
  not g14759 (n_6944, n8169);
  and g14760 (n8170, n8157, n_6944);
  and g14761 (n8171, n_6943, n_6944);
  not g14762 (n_6945, n8170);
  not g14763 (n_6946, n8171);
  and g14764 (n8172, n_6945, n_6946);
  and g14765 (n8173, n_6684, n_6690);
  and g14766 (n8174, n8172, n8173);
  not g14767 (n_6947, n8172);
  not g14768 (n_6948, n8173);
  and g14769 (n8175, n_6947, n_6948);
  not g14770 (n_6949, n8174);
  not g14771 (n_6950, n8175);
  and g14772 (n8176, n_6949, n_6950);
  and g14773 (n8177, \b[24] , n2539);
  and g14774 (n8178, \b[22] , n2685);
  and g14775 (n8179, \b[23] , n2534);
  and g14781 (n8182, n2458, n2542);
  not g14784 (n_6955, n8183);
  and g14785 (n8184, \a[26] , n_6955);
  not g14786 (n_6956, n8184);
  and g14787 (n8185, \a[26] , n_6956);
  and g14788 (n8186, n_6955, n_6956);
  not g14789 (n_6957, n8185);
  not g14790 (n_6958, n8186);
  and g14791 (n8187, n_6957, n_6958);
  not g14792 (n_6959, n8176);
  and g14793 (n8188, n_6959, n8187);
  not g14794 (n_6960, n8187);
  and g14795 (n8189, n8176, n_6960);
  not g14796 (n_6961, n8188);
  not g14797 (n_6962, n8189);
  and g14798 (n8190, n_6961, n_6962);
  not g14799 (n_6963, n7894);
  and g14800 (n8191, n_6963, n8190);
  not g14801 (n_6964, n8190);
  and g14802 (n8192, n7894, n_6964);
  not g14803 (n_6965, n8191);
  not g14804 (n_6966, n8192);
  and g14805 (n8193, n_6965, n_6966);
  not g14806 (n_6967, n8042);
  and g14807 (n8194, n_6967, n8193);
  not g14808 (n_6968, n8194);
  and g14809 (n8195, n8193, n_6968);
  and g14810 (n8196, n_6967, n_6968);
  not g14811 (n_6969, n8195);
  not g14812 (n_6970, n8196);
  and g14813 (n8197, n_6969, n_6970);
  not g14814 (n_6971, n8031);
  and g14815 (n8198, n_6971, n8197);
  not g14816 (n_6972, n8197);
  and g14817 (n8199, n8031, n_6972);
  not g14818 (n_6973, n8198);
  not g14819 (n_6974, n8199);
  and g14820 (n8200, n_6973, n_6974);
  and g14821 (n8201, \b[30] , n1627);
  and g14822 (n8202, \b[28] , n1763);
  and g14823 (n8203, \b[29] , n1622);
  and g14829 (n8206, n1630, n3577);
  not g14832 (n_6979, n8207);
  and g14833 (n8208, \a[20] , n_6979);
  not g14834 (n_6980, n8208);
  and g14835 (n8209, \a[20] , n_6980);
  and g14836 (n8210, n_6979, n_6980);
  not g14837 (n_6981, n8209);
  not g14838 (n_6982, n8210);
  and g14839 (n8211, n_6981, n_6982);
  not g14840 (n_6983, n8200);
  not g14841 (n_6984, n8211);
  and g14842 (n8212, n_6983, n_6984);
  and g14843 (n8213, n8200, n8211);
  not g14844 (n_6985, n8212);
  not g14845 (n_6986, n8213);
  and g14846 (n8214, n_6985, n_6986);
  not g14847 (n_6987, n8030);
  and g14848 (n8215, n_6987, n8214);
  not g14849 (n_6988, n8214);
  and g14850 (n8216, n8030, n_6988);
  not g14851 (n_6989, n8215);
  not g14852 (n_6990, n8216);
  and g14853 (n8217, n_6989, n_6990);
  not g14854 (n_6991, n8029);
  and g14855 (n8218, n_6991, n8217);
  not g14856 (n_6992, n8218);
  and g14857 (n8219, n8217, n_6992);
  and g14858 (n8220, n_6991, n_6992);
  not g14859 (n_6993, n8219);
  not g14860 (n_6994, n8220);
  and g14861 (n8221, n_6993, n_6994);
  not g14862 (n_6995, n8018);
  and g14863 (n8222, n_6995, n8221);
  not g14864 (n_6996, n8221);
  and g14865 (n8223, n8018, n_6996);
  not g14866 (n_6997, n8222);
  not g14867 (n_6998, n8223);
  and g14868 (n8224, n_6997, n_6998);
  and g14869 (n8225, \b[36] , n951);
  and g14870 (n8226, \b[34] , n1056);
  and g14871 (n8227, \b[35] , n946);
  and g14877 (n8230, n954, n4922);
  not g14880 (n_7003, n8231);
  and g14881 (n8232, \a[14] , n_7003);
  not g14882 (n_7004, n8232);
  and g14883 (n8233, \a[14] , n_7004);
  and g14884 (n8234, n_7003, n_7004);
  not g14885 (n_7005, n8233);
  not g14886 (n_7006, n8234);
  and g14887 (n8235, n_7005, n_7006);
  not g14888 (n_7007, n8224);
  not g14889 (n_7008, n8235);
  and g14890 (n8236, n_7007, n_7008);
  and g14891 (n8237, n8224, n8235);
  not g14892 (n_7009, n8236);
  not g14893 (n_7010, n8237);
  and g14894 (n8238, n_7009, n_7010);
  not g14895 (n_7011, n8238);
  and g14896 (n8239, n8017, n_7011);
  not g14897 (n_7012, n8017);
  and g14898 (n8240, n_7012, n8238);
  not g14899 (n_7013, n8239);
  not g14900 (n_7014, n8240);
  and g14901 (n8241, n_7013, n_7014);
  and g14902 (n8242, \b[39] , n700);
  and g14903 (n8243, \b[37] , n767);
  and g14904 (n8244, \b[38] , n695);
  and g14910 (n8247, n703, n5451);
  not g14913 (n_7019, n8248);
  and g14914 (n8249, \a[11] , n_7019);
  not g14915 (n_7020, n8249);
  and g14916 (n8250, \a[11] , n_7020);
  and g14917 (n8251, n_7019, n_7020);
  not g14918 (n_7021, n8250);
  not g14919 (n_7022, n8251);
  and g14920 (n8252, n_7021, n_7022);
  not g14921 (n_7023, n8252);
  and g14922 (n8253, n8241, n_7023);
  not g14923 (n_7024, n8253);
  and g14924 (n8254, n8241, n_7024);
  and g14925 (n8255, n_7023, n_7024);
  not g14926 (n_7025, n8254);
  not g14927 (n_7026, n8255);
  and g14928 (n8256, n_7025, n_7026);
  and g14929 (n8257, n_6756, n_6762);
  and g14930 (n8258, n8256, n8257);
  not g14931 (n_7027, n8256);
  not g14932 (n_7028, n8257);
  and g14933 (n8259, n_7027, n_7028);
  not g14934 (n_7029, n8258);
  not g14935 (n_7030, n8259);
  and g14936 (n8260, n_7029, n_7030);
  and g14937 (n8261, \b[42] , n511);
  and g14938 (n8262, \b[40] , n541);
  and g14939 (n8263, \b[41] , n506);
  and g14945 (n8266, n514, n6489);
  not g14948 (n_7035, n8267);
  and g14949 (n8268, \a[8] , n_7035);
  not g14950 (n_7036, n8268);
  and g14951 (n8269, \a[8] , n_7036);
  and g14952 (n8270, n_7035, n_7036);
  not g14953 (n_7037, n8269);
  not g14954 (n_7038, n8270);
  and g14955 (n8271, n_7037, n_7038);
  not g14956 (n_7039, n8271);
  and g14957 (n8272, n8260, n_7039);
  not g14958 (n_7040, n8272);
  and g14959 (n8273, n8260, n_7040);
  and g14960 (n8274, n_7039, n_7040);
  not g14961 (n_7041, n8273);
  not g14962 (n_7042, n8274);
  and g14963 (n8275, n_7041, n_7042);
  not g14964 (n_7043, n7969);
  and g14965 (n8276, n_7043, n8275);
  not g14966 (n_7044, n8275);
  and g14967 (n8277, n7969, n_7044);
  not g14968 (n_7045, n8276);
  not g14969 (n_7046, n8277);
  and g14970 (n8278, n_7045, n_7046);
  and g14971 (n8279, \b[45] , n362);
  and g14972 (n8280, \b[43] , n403);
  and g14973 (n8281, \b[44] , n357);
  and g14979 (n8284, n365, n7361);
  not g14982 (n_7051, n8285);
  and g14983 (n8286, \a[5] , n_7051);
  not g14984 (n_7052, n8286);
  and g14985 (n8287, \a[5] , n_7052);
  and g14986 (n8288, n_7051, n_7052);
  not g14987 (n_7053, n8287);
  not g14988 (n_7054, n8288);
  and g14989 (n8289, n_7053, n_7054);
  not g14990 (n_7055, n8278);
  not g14991 (n_7056, n8289);
  and g14992 (n8290, n_7055, n_7056);
  and g14993 (n8291, n8278, n8289);
  not g14994 (n_7057, n8290);
  not g14995 (n_7058, n8291);
  and g14996 (n8292, n_7057, n_7058);
  not g14997 (n_7059, n8016);
  and g14998 (n8293, n_7059, n8292);
  not g14999 (n_7060, n8292);
  and g15000 (n8294, n8016, n_7060);
  not g15001 (n_7061, n8293);
  not g15002 (n_7062, n8294);
  and g15003 (n8295, n_7061, n_7062);
  not g15004 (n_7063, n8295);
  and g15005 (n8296, n8015, n_7063);
  not g15006 (n_7064, n8015);
  and g15007 (n8297, n_7064, n8295);
  not g15008 (n_7065, n8296);
  not g15009 (n_7066, n8297);
  and g15010 (n8298, n_7065, n_7066);
  not g15011 (n_7067, n7997);
  and g15012 (n8299, n_7067, n8298);
  not g15013 (n_7068, n8298);
  and g15014 (n8300, n7997, n_7068);
  not g15015 (n_7069, n8299);
  not g15016 (n_7070, n8300);
  and g15017 (\f[48] , n_7069, n_7070);
  and g15018 (n8302, n_7066, n_7069);
  and g15019 (n8303, n_6971, n_6972);
  not g15020 (n_7071, n8303);
  and g15021 (n8304, n_6968, n_7071);
  and g15022 (n8305, \b[28] , n2048);
  and g15023 (n8306, \b[26] , n2198);
  and g15024 (n8307, \b[27] , n2043);
  and g15030 (n8310, n2051, n3189);
  not g15033 (n_7076, n8311);
  and g15034 (n8312, \a[23] , n_7076);
  not g15035 (n_7077, n8312);
  and g15036 (n8313, \a[23] , n_7077);
  and g15037 (n8314, n_7076, n_7077);
  not g15038 (n_7078, n8313);
  not g15039 (n_7079, n8314);
  and g15040 (n8315, n_7078, n_7079);
  and g15041 (n8316, \b[16] , n4287);
  and g15042 (n8317, \b[14] , n4532);
  and g15043 (n8318, \b[15] , n4282);
  and g15049 (n8321, n1237, n4290);
  not g15052 (n_7084, n8322);
  and g15053 (n8323, \a[35] , n_7084);
  not g15054 (n_7085, n8323);
  and g15055 (n8324, \a[35] , n_7085);
  and g15056 (n8325, n_7084, n_7085);
  not g15057 (n_7086, n8324);
  not g15058 (n_7087, n8325);
  and g15059 (n8326, n_7086, n_7087);
  and g15060 (n8327, n_6904, n_6909);
  and g15061 (n8328, n_6898, n_6901);
  and g15062 (n8329, \b[7] , n6595);
  and g15063 (n8330, \b[5] , n6902);
  and g15064 (n8331, \b[6] , n6590);
  and g15070 (n8334, n484, n6598);
  not g15073 (n_7092, n8335);
  and g15074 (n8336, \a[44] , n_7092);
  not g15075 (n_7093, n8336);
  and g15076 (n8337, \a[44] , n_7093);
  and g15077 (n8338, n_7092, n_7093);
  not g15078 (n_7094, n8337);
  not g15079 (n_7095, n8338);
  and g15080 (n8339, n_7094, n_7095);
  and g15081 (n8340, n7799, n8082);
  not g15082 (n_7096, n8340);
  and g15083 (n8341, n_6877, n_7096);
  and g15084 (n8342, \b[4] , n7446);
  and g15085 (n8343, \b[2] , n7787);
  and g15086 (n8344, \b[3] , n7441);
  and g15092 (n8347, n346, n7449);
  not g15095 (n_7101, n8348);
  and g15096 (n8349, \a[47] , n_7101);
  not g15097 (n_7102, n8349);
  and g15098 (n8350, \a[47] , n_7102);
  and g15099 (n8351, n_7101, n_7102);
  not g15100 (n_7103, n8350);
  not g15101 (n_7104, n8351);
  and g15102 (n8352, n_7103, n_7104);
  and g15103 (n8353, \a[50] , n_6864);
  and g15104 (n8354, n_6860, \a[49] );
  not g15105 (n_7107, \a[49] );
  and g15106 (n8355, \a[48] , n_7107);
  not g15107 (n_7108, n8354);
  not g15108 (n_7109, n8355);
  and g15109 (n8356, n_7108, n_7109);
  not g15110 (n_7110, n8356);
  and g15111 (n8357, n8081, n_7110);
  and g15112 (n8358, \b[0] , n8357);
  and g15113 (n8359, n_7107, \a[50] );
  not g15114 (n_7111, \a[50] );
  and g15115 (n8360, \a[49] , n_7111);
  not g15116 (n_7112, n8359);
  not g15117 (n_7113, n8360);
  and g15118 (n8361, n_7112, n_7113);
  and g15119 (n8362, n_6863, n8361);
  and g15120 (n8363, \b[1] , n8362);
  not g15121 (n_7114, n8358);
  not g15122 (n_7115, n8363);
  and g15123 (n8364, n_7114, n_7115);
  not g15124 (n_7116, n8361);
  and g15125 (n8365, n_6863, n_7116);
  and g15126 (n8366, n_21, n8365);
  not g15127 (n_7117, n8366);
  and g15128 (n8367, n8364, n_7117);
  not g15129 (n_7118, n8367);
  and g15130 (n8368, \a[50] , n_7118);
  not g15131 (n_7119, n8368);
  and g15132 (n8369, \a[50] , n_7119);
  and g15133 (n8370, n_7118, n_7119);
  not g15134 (n_7120, n8369);
  not g15135 (n_7121, n8370);
  and g15136 (n8371, n_7120, n_7121);
  not g15137 (n_7122, n8371);
  and g15138 (n8372, n8353, n_7122);
  not g15139 (n_7123, n8353);
  and g15140 (n8373, n_7123, n8371);
  not g15141 (n_7124, n8372);
  not g15142 (n_7125, n8373);
  and g15143 (n8374, n_7124, n_7125);
  not g15144 (n_7126, n8374);
  and g15145 (n8375, n8352, n_7126);
  not g15146 (n_7127, n8352);
  and g15147 (n8376, n_7127, n8374);
  not g15148 (n_7128, n8375);
  not g15149 (n_7129, n8376);
  and g15150 (n8377, n_7128, n_7129);
  not g15151 (n_7130, n8341);
  and g15152 (n8378, n_7130, n8377);
  not g15153 (n_7131, n8377);
  and g15154 (n8379, n8341, n_7131);
  not g15155 (n_7132, n8378);
  not g15156 (n_7133, n8379);
  and g15157 (n8380, n_7132, n_7133);
  not g15158 (n_7134, n8339);
  and g15159 (n8381, n_7134, n8380);
  not g15160 (n_7135, n8381);
  and g15161 (n8382, n8380, n_7135);
  and g15162 (n8383, n_7134, n_7135);
  not g15163 (n_7136, n8382);
  not g15164 (n_7137, n8383);
  and g15165 (n8384, n_7136, n_7137);
  and g15166 (n8385, n_6880, n_6886);
  and g15167 (n8386, n8384, n8385);
  not g15168 (n_7138, n8384);
  not g15169 (n_7139, n8385);
  and g15170 (n8387, n_7138, n_7139);
  not g15171 (n_7140, n8386);
  not g15172 (n_7141, n8387);
  and g15173 (n8388, n_7140, n_7141);
  and g15174 (n8389, \b[10] , n5777);
  and g15175 (n8390, \b[8] , n6059);
  and g15176 (n8391, \b[9] , n5772);
  and g15182 (n8394, n738, n5780);
  not g15185 (n_7146, n8395);
  and g15186 (n8396, \a[41] , n_7146);
  not g15187 (n_7147, n8396);
  and g15188 (n8397, \a[41] , n_7147);
  and g15189 (n8398, n_7146, n_7147);
  not g15190 (n_7148, n8397);
  not g15191 (n_7149, n8398);
  and g15192 (n8399, n_7148, n_7149);
  not g15193 (n_7150, n8399);
  and g15194 (n8400, n8388, n_7150);
  not g15195 (n_7151, n8388);
  and g15196 (n8401, n_7151, n8399);
  not g15197 (n_7152, n8328);
  not g15198 (n_7153, n8401);
  and g15199 (n8402, n_7152, n_7153);
  not g15200 (n_7154, n8400);
  and g15201 (n8403, n_7154, n8402);
  not g15202 (n_7155, n8403);
  and g15203 (n8404, n_7152, n_7155);
  and g15204 (n8405, n_7154, n_7155);
  and g15205 (n8406, n_7153, n8405);
  not g15206 (n_7156, n8404);
  not g15207 (n_7157, n8406);
  and g15208 (n8407, n_7156, n_7157);
  and g15209 (n8408, \b[13] , n5035);
  and g15210 (n8409, \b[11] , n5277);
  and g15211 (n8410, \b[12] , n5030);
  and g15217 (n8413, n1008, n5038);
  not g15220 (n_7162, n8414);
  and g15221 (n8415, \a[38] , n_7162);
  not g15222 (n_7163, n8415);
  and g15223 (n8416, \a[38] , n_7163);
  and g15224 (n8417, n_7162, n_7163);
  not g15225 (n_7164, n8416);
  not g15226 (n_7165, n8417);
  and g15227 (n8418, n_7164, n_7165);
  and g15228 (n8419, n8407, n8418);
  not g15229 (n_7166, n8407);
  not g15230 (n_7167, n8418);
  and g15231 (n8420, n_7166, n_7167);
  not g15232 (n_7168, n8419);
  not g15233 (n_7169, n8420);
  and g15234 (n8421, n_7168, n_7169);
  not g15235 (n_7170, n8327);
  and g15236 (n8422, n_7170, n8421);
  not g15237 (n_7171, n8421);
  and g15238 (n8423, n8327, n_7171);
  not g15239 (n_7172, n8422);
  not g15240 (n_7173, n8423);
  and g15241 (n8424, n_7172, n_7173);
  not g15242 (n_7174, n8326);
  and g15243 (n8425, n_7174, n8424);
  not g15244 (n_7175, n8425);
  and g15245 (n8426, n8424, n_7175);
  and g15246 (n8427, n_7174, n_7175);
  not g15247 (n_7176, n8426);
  not g15248 (n_7177, n8427);
  and g15249 (n8428, n_7176, n_7177);
  and g15250 (n8429, n_6913, n_6917);
  and g15251 (n8430, n8428, n8429);
  not g15252 (n_7178, n8428);
  not g15253 (n_7179, n8429);
  and g15254 (n8431, n_7178, n_7179);
  not g15255 (n_7180, n8430);
  not g15256 (n_7181, n8431);
  and g15257 (n8432, n_7180, n_7181);
  and g15258 (n8433, \b[19] , n3638);
  and g15259 (n8434, \b[17] , n3843);
  and g15260 (n8435, \b[18] , n3633);
  and g15266 (n8438, n1708, n3641);
  not g15269 (n_7186, n8439);
  and g15270 (n8440, \a[32] , n_7186);
  not g15271 (n_7187, n8440);
  and g15272 (n8441, \a[32] , n_7187);
  and g15273 (n8442, n_7186, n_7187);
  not g15274 (n_7188, n8441);
  not g15275 (n_7189, n8442);
  and g15276 (n8443, n_7188, n_7189);
  not g15277 (n_7190, n8443);
  and g15278 (n8444, n8432, n_7190);
  not g15279 (n_7191, n8444);
  and g15280 (n8445, n8432, n_7191);
  and g15281 (n8446, n_7190, n_7191);
  not g15282 (n_7192, n8445);
  not g15283 (n_7193, n8446);
  and g15284 (n8447, n_7192, n_7193);
  and g15285 (n8448, n_6928, n_6934);
  and g15286 (n8449, n8447, n8448);
  not g15287 (n_7194, n8447);
  not g15288 (n_7195, n8448);
  and g15289 (n8450, n_7194, n_7195);
  not g15290 (n_7196, n8449);
  not g15291 (n_7197, n8450);
  and g15292 (n8451, n_7196, n_7197);
  and g15293 (n8452, \b[22] , n3050);
  and g15294 (n8453, \b[20] , n3243);
  and g15295 (n8454, \b[21] , n3045);
  and g15301 (n8457, n2145, n3053);
  not g15304 (n_7202, n8458);
  and g15305 (n8459, \a[29] , n_7202);
  not g15306 (n_7203, n8459);
  and g15307 (n8460, \a[29] , n_7203);
  and g15308 (n8461, n_7202, n_7203);
  not g15309 (n_7204, n8460);
  not g15310 (n_7205, n8461);
  and g15311 (n8462, n_7204, n_7205);
  not g15312 (n_7206, n8462);
  and g15313 (n8463, n8451, n_7206);
  not g15314 (n_7207, n8463);
  and g15315 (n8464, n8451, n_7207);
  and g15316 (n8465, n_7206, n_7207);
  not g15317 (n_7208, n8464);
  not g15318 (n_7209, n8465);
  and g15319 (n8466, n_7208, n_7209);
  and g15320 (n8467, n_6944, n_6950);
  and g15321 (n8468, n8466, n8467);
  not g15322 (n_7210, n8466);
  not g15323 (n_7211, n8467);
  and g15324 (n8469, n_7210, n_7211);
  not g15325 (n_7212, n8468);
  not g15326 (n_7213, n8469);
  and g15327 (n8470, n_7212, n_7213);
  and g15328 (n8471, \b[25] , n2539);
  and g15329 (n8472, \b[23] , n2685);
  and g15330 (n8473, \b[24] , n2534);
  and g15336 (n8476, n2485, n2542);
  not g15339 (n_7218, n8477);
  and g15340 (n8478, \a[26] , n_7218);
  not g15341 (n_7219, n8478);
  and g15342 (n8479, \a[26] , n_7219);
  and g15343 (n8480, n_7218, n_7219);
  not g15344 (n_7220, n8479);
  not g15345 (n_7221, n8480);
  and g15346 (n8481, n_7220, n_7221);
  not g15347 (n_7222, n8481);
  and g15348 (n8482, n8470, n_7222);
  not g15349 (n_7223, n8482);
  and g15350 (n8483, n8470, n_7223);
  and g15351 (n8484, n_7222, n_7223);
  not g15352 (n_7224, n8483);
  not g15353 (n_7225, n8484);
  and g15354 (n8485, n_7224, n_7225);
  and g15355 (n8486, n_6962, n_6965);
  not g15356 (n_7226, n8485);
  not g15357 (n_7227, n8486);
  and g15358 (n8487, n_7226, n_7227);
  and g15359 (n8488, n8485, n8486);
  not g15360 (n_7228, n8487);
  not g15361 (n_7229, n8488);
  and g15362 (n8489, n_7228, n_7229);
  not g15363 (n_7230, n8315);
  and g15364 (n8490, n_7230, n8489);
  not g15365 (n_7231, n8490);
  and g15366 (n8491, n_7230, n_7231);
  and g15367 (n8492, n8489, n_7231);
  not g15368 (n_7232, n8491);
  not g15369 (n_7233, n8492);
  and g15370 (n8493, n_7232, n_7233);
  not g15371 (n_7234, n8304);
  not g15372 (n_7235, n8493);
  and g15373 (n8494, n_7234, n_7235);
  not g15374 (n_7236, n8494);
  and g15375 (n8495, n_7234, n_7236);
  and g15376 (n8496, n_7235, n_7236);
  not g15377 (n_7237, n8495);
  not g15378 (n_7238, n8496);
  and g15379 (n8497, n_7237, n_7238);
  and g15380 (n8498, \b[31] , n1627);
  and g15381 (n8499, \b[29] , n1763);
  and g15382 (n8500, \b[30] , n1622);
  and g15388 (n8503, n1630, n3796);
  not g15391 (n_7243, n8504);
  and g15392 (n8505, \a[20] , n_7243);
  not g15393 (n_7244, n8505);
  and g15394 (n8506, \a[20] , n_7244);
  and g15395 (n8507, n_7243, n_7244);
  not g15396 (n_7245, n8506);
  not g15397 (n_7246, n8507);
  and g15398 (n8508, n_7245, n_7246);
  not g15399 (n_7247, n8497);
  not g15400 (n_7248, n8508);
  and g15401 (n8509, n_7247, n_7248);
  not g15402 (n_7249, n8509);
  and g15403 (n8510, n_7247, n_7249);
  and g15404 (n8511, n_7248, n_7249);
  not g15405 (n_7250, n8510);
  not g15406 (n_7251, n8511);
  and g15407 (n8512, n_7250, n_7251);
  and g15408 (n8513, n_6985, n_6989);
  and g15409 (n8514, n8512, n8513);
  not g15410 (n_7252, n8512);
  not g15411 (n_7253, n8513);
  and g15412 (n8515, n_7252, n_7253);
  not g15413 (n_7254, n8514);
  not g15414 (n_7255, n8515);
  and g15415 (n8516, n_7254, n_7255);
  and g15416 (n8517, \b[34] , n1302);
  and g15417 (n8518, \b[32] , n1391);
  and g15418 (n8519, \b[33] , n1297);
  and g15424 (n8522, n1305, n4466);
  not g15427 (n_7260, n8523);
  and g15428 (n8524, \a[17] , n_7260);
  not g15429 (n_7261, n8524);
  and g15430 (n8525, \a[17] , n_7261);
  and g15431 (n8526, n_7260, n_7261);
  not g15432 (n_7262, n8525);
  not g15433 (n_7263, n8526);
  and g15434 (n8527, n_7262, n_7263);
  not g15435 (n_7264, n8527);
  and g15436 (n8528, n8516, n_7264);
  not g15437 (n_7265, n8528);
  and g15438 (n8529, n8516, n_7265);
  and g15439 (n8530, n_7264, n_7265);
  not g15440 (n_7266, n8529);
  not g15441 (n_7267, n8530);
  and g15442 (n8531, n_7266, n_7267);
  and g15443 (n8532, n_6995, n_6996);
  not g15444 (n_7268, n8532);
  and g15445 (n8533, n_6992, n_7268);
  and g15446 (n8534, n8531, n8533);
  not g15447 (n_7269, n8531);
  not g15448 (n_7270, n8533);
  and g15449 (n8535, n_7269, n_7270);
  not g15450 (n_7271, n8534);
  not g15451 (n_7272, n8535);
  and g15452 (n8536, n_7271, n_7272);
  and g15453 (n8537, \b[37] , n951);
  and g15454 (n8538, \b[35] , n1056);
  and g15455 (n8539, \b[36] , n946);
  and g15461 (n8542, n954, n5181);
  not g15464 (n_7277, n8543);
  and g15465 (n8544, \a[14] , n_7277);
  not g15466 (n_7278, n8544);
  and g15467 (n8545, \a[14] , n_7278);
  and g15468 (n8546, n_7277, n_7278);
  not g15469 (n_7279, n8545);
  not g15470 (n_7280, n8546);
  and g15471 (n8547, n_7279, n_7280);
  not g15472 (n_7281, n8547);
  and g15473 (n8548, n8536, n_7281);
  not g15474 (n_7282, n8548);
  and g15475 (n8549, n8536, n_7282);
  and g15476 (n8550, n_7281, n_7282);
  not g15477 (n_7283, n8549);
  not g15478 (n_7284, n8550);
  and g15479 (n8551, n_7283, n_7284);
  and g15480 (n8552, n_7009, n_7014);
  and g15481 (n8553, n8551, n8552);
  not g15482 (n_7285, n8551);
  not g15483 (n_7286, n8552);
  and g15484 (n8554, n_7285, n_7286);
  not g15485 (n_7287, n8553);
  not g15486 (n_7288, n8554);
  and g15487 (n8555, n_7287, n_7288);
  and g15488 (n8556, \b[40] , n700);
  and g15489 (n8557, \b[38] , n767);
  and g15490 (n8558, \b[39] , n695);
  and g15496 (n8561, n703, n5955);
  not g15499 (n_7293, n8562);
  and g15500 (n8563, \a[11] , n_7293);
  not g15501 (n_7294, n8563);
  and g15502 (n8564, \a[11] , n_7294);
  and g15503 (n8565, n_7293, n_7294);
  not g15504 (n_7295, n8564);
  not g15505 (n_7296, n8565);
  and g15506 (n8566, n_7295, n_7296);
  not g15507 (n_7297, n8566);
  and g15508 (n8567, n8555, n_7297);
  not g15509 (n_7298, n8567);
  and g15510 (n8568, n8555, n_7298);
  and g15511 (n8569, n_7297, n_7298);
  not g15512 (n_7299, n8568);
  not g15513 (n_7300, n8569);
  and g15514 (n8570, n_7299, n_7300);
  and g15515 (n8571, n_7024, n_7030);
  and g15516 (n8572, n8570, n8571);
  not g15517 (n_7301, n8570);
  not g15518 (n_7302, n8571);
  and g15519 (n8573, n_7301, n_7302);
  not g15520 (n_7303, n8572);
  not g15521 (n_7304, n8573);
  and g15522 (n8574, n_7303, n_7304);
  and g15523 (n8575, \b[43] , n511);
  and g15524 (n8576, \b[41] , n541);
  and g15525 (n8577, \b[42] , n506);
  and g15531 (n8580, n514, n6515);
  not g15534 (n_7309, n8581);
  and g15535 (n8582, \a[8] , n_7309);
  not g15536 (n_7310, n8582);
  and g15537 (n8583, \a[8] , n_7310);
  and g15538 (n8584, n_7309, n_7310);
  not g15539 (n_7311, n8583);
  not g15540 (n_7312, n8584);
  and g15541 (n8585, n_7311, n_7312);
  not g15542 (n_7313, n8585);
  and g15543 (n8586, n8574, n_7313);
  not g15544 (n_7314, n8586);
  and g15545 (n8587, n8574, n_7314);
  and g15546 (n8588, n_7313, n_7314);
  not g15547 (n_7315, n8587);
  not g15548 (n_7316, n8588);
  and g15549 (n8589, n_7315, n_7316);
  and g15550 (n8590, n_7043, n_7044);
  not g15551 (n_7317, n8590);
  and g15552 (n8591, n_7040, n_7317);
  and g15553 (n8592, n8589, n8591);
  not g15554 (n_7318, n8589);
  not g15555 (n_7319, n8591);
  and g15556 (n8593, n_7318, n_7319);
  not g15557 (n_7320, n8592);
  not g15558 (n_7321, n8593);
  and g15559 (n8594, n_7320, n_7321);
  and g15560 (n8595, \b[46] , n362);
  and g15561 (n8596, \b[44] , n403);
  and g15562 (n8597, \b[45] , n357);
  and g15568 (n8600, n365, n7677);
  not g15571 (n_7326, n8601);
  and g15572 (n8602, \a[5] , n_7326);
  not g15573 (n_7327, n8602);
  and g15574 (n8603, \a[5] , n_7327);
  and g15575 (n8604, n_7326, n_7327);
  not g15576 (n_7328, n8603);
  not g15577 (n_7329, n8604);
  and g15578 (n8605, n_7328, n_7329);
  not g15579 (n_7330, n8605);
  and g15580 (n8606, n8594, n_7330);
  not g15581 (n_7331, n8606);
  and g15582 (n8607, n8594, n_7331);
  and g15583 (n8608, n_7330, n_7331);
  not g15584 (n_7332, n8607);
  not g15585 (n_7333, n8608);
  and g15586 (n8609, n_7332, n_7333);
  and g15587 (n8610, n_7057, n_7061);
  and g15588 (n8611, n8609, n8610);
  not g15589 (n_7334, n8609);
  not g15590 (n_7335, n8610);
  and g15591 (n8612, n_7334, n_7335);
  not g15592 (n_7336, n8611);
  not g15593 (n_7337, n8612);
  and g15594 (n8613, n_7336, n_7337);
  and g15595 (n8614, \b[49] , n266);
  and g15596 (n8615, \b[47] , n284);
  and g15597 (n8616, \b[48] , n261);
  and g15603 (n8619, n_6809, n_6812);
  not g15604 (n_7342, \b[49] );
  and g15605 (n8620, n_6807, n_7342);
  and g15606 (n8621, \b[48] , \b[49] );
  not g15607 (n_7343, n8620);
  not g15608 (n_7344, n8621);
  and g15609 (n8622, n_7343, n_7344);
  not g15610 (n_7345, n8619);
  and g15611 (n8623, n_7345, n8622);
  not g15612 (n_7346, n8622);
  and g15613 (n8624, n8619, n_7346);
  not g15614 (n_7347, n8623);
  not g15615 (n_7348, n8624);
  and g15616 (n8625, n_7347, n_7348);
  and g15617 (n8626, n269, n8625);
  not g15620 (n_7350, n8627);
  and g15621 (n8628, \a[2] , n_7350);
  not g15622 (n_7351, n8628);
  and g15623 (n8629, \a[2] , n_7351);
  and g15624 (n8630, n_7350, n_7351);
  not g15625 (n_7352, n8629);
  not g15626 (n_7353, n8630);
  and g15627 (n8631, n_7352, n_7353);
  not g15628 (n_7354, n8613);
  and g15629 (n8632, n_7354, n8631);
  not g15630 (n_7355, n8631);
  and g15631 (n8633, n8613, n_7355);
  not g15632 (n_7356, n8632);
  not g15633 (n_7357, n8633);
  and g15634 (n8634, n_7356, n_7357);
  not g15635 (n_7358, n8302);
  and g15636 (n8635, n_7358, n8634);
  not g15637 (n_7359, n8634);
  and g15638 (n8636, n8302, n_7359);
  not g15639 (n_7360, n8635);
  not g15640 (n_7361, n8636);
  and g15641 (\f[49] , n_7360, n_7361);
  and g15642 (n8638, n_7314, n_7321);
  and g15643 (n8639, \b[35] , n1302);
  and g15644 (n8640, \b[33] , n1391);
  and g15645 (n8641, \b[34] , n1297);
  and g15651 (n8644, n1305, n4696);
  not g15654 (n_7366, n8645);
  and g15655 (n8646, \a[17] , n_7366);
  not g15656 (n_7367, n8646);
  and g15657 (n8647, \a[17] , n_7367);
  and g15658 (n8648, n_7366, n_7367);
  not g15659 (n_7368, n8647);
  not g15660 (n_7369, n8648);
  and g15661 (n8649, n_7368, n_7369);
  and g15662 (n8650, n_7249, n_7255);
  and g15663 (n8651, \b[32] , n1627);
  and g15664 (n8652, \b[30] , n1763);
  and g15665 (n8653, \b[31] , n1622);
  and g15671 (n8656, n1630, n4013);
  not g15674 (n_7374, n8657);
  and g15675 (n8658, \a[20] , n_7374);
  not g15676 (n_7375, n8658);
  and g15677 (n8659, \a[20] , n_7375);
  and g15678 (n8660, n_7374, n_7375);
  not g15679 (n_7376, n8659);
  not g15680 (n_7377, n8660);
  and g15681 (n8661, n_7376, n_7377);
  and g15682 (n8662, n_7231, n_7236);
  and g15683 (n8663, \b[29] , n2048);
  and g15684 (n8664, \b[27] , n2198);
  and g15685 (n8665, \b[28] , n2043);
  and g15691 (n8668, n2051, n3383);
  not g15694 (n_7382, n8669);
  and g15695 (n8670, \a[23] , n_7382);
  not g15696 (n_7383, n8670);
  and g15697 (n8671, \a[23] , n_7383);
  and g15698 (n8672, n_7382, n_7383);
  not g15699 (n_7384, n8671);
  not g15700 (n_7385, n8672);
  and g15701 (n8673, n_7384, n_7385);
  and g15702 (n8674, n_7223, n_7228);
  and g15703 (n8675, n_7207, n_7213);
  and g15704 (n8676, n_7175, n_7181);
  and g15705 (n8677, \b[17] , n4287);
  and g15706 (n8678, \b[15] , n4532);
  and g15707 (n8679, \b[16] , n4282);
  and g15713 (n8682, n1356, n4290);
  not g15716 (n_7390, n8683);
  and g15717 (n8684, \a[35] , n_7390);
  not g15718 (n_7391, n8684);
  and g15719 (n8685, \a[35] , n_7391);
  and g15720 (n8686, n_7390, n_7391);
  not g15721 (n_7392, n8685);
  not g15722 (n_7393, n8686);
  and g15723 (n8687, n_7392, n_7393);
  and g15724 (n8688, n_7169, n_7172);
  and g15725 (n8689, \b[14] , n5035);
  and g15726 (n8690, \b[12] , n5277);
  and g15727 (n8691, \b[13] , n5030);
  and g15733 (n8694, n1034, n5038);
  not g15736 (n_7398, n8695);
  and g15737 (n8696, \a[38] , n_7398);
  not g15738 (n_7399, n8696);
  and g15739 (n8697, \a[38] , n_7399);
  and g15740 (n8698, n_7398, n_7399);
  not g15741 (n_7400, n8697);
  not g15742 (n_7401, n8698);
  and g15743 (n8699, n_7400, n_7401);
  and g15744 (n8700, n_7135, n_7141);
  and g15745 (n8701, \b[8] , n6595);
  and g15746 (n8702, \b[6] , n6902);
  and g15747 (n8703, \b[7] , n6590);
  and g15753 (n8706, n585, n6598);
  not g15756 (n_7406, n8707);
  and g15757 (n8708, \a[44] , n_7406);
  not g15758 (n_7407, n8708);
  and g15759 (n8709, \a[44] , n_7407);
  and g15760 (n8710, n_7406, n_7407);
  not g15761 (n_7408, n8709);
  not g15762 (n_7409, n8710);
  and g15763 (n8711, n_7408, n_7409);
  and g15764 (n8712, n_7129, n_7132);
  and g15765 (n8713, \b[2] , n8362);
  and g15766 (n8714, n8081, n_7116);
  and g15767 (n8715, n8356, n8714);
  and g15768 (n8716, \b[0] , n8715);
  and g15769 (n8717, \b[1] , n8357);
  and g15775 (n8720, n296, n8365);
  not g15778 (n_7414, n8721);
  and g15779 (n8722, \a[50] , n_7414);
  not g15780 (n_7415, n8722);
  and g15781 (n8723, \a[50] , n_7415);
  and g15782 (n8724, n_7414, n_7415);
  not g15783 (n_7416, n8723);
  not g15784 (n_7417, n8724);
  and g15785 (n8725, n_7416, n_7417);
  and g15786 (n8726, n_7124, n8725);
  not g15787 (n_7418, n8725);
  and g15788 (n8727, n8372, n_7418);
  not g15789 (n_7419, n8726);
  not g15790 (n_7420, n8727);
  and g15791 (n8728, n_7419, n_7420);
  and g15792 (n8729, \b[5] , n7446);
  and g15793 (n8730, \b[3] , n7787);
  and g15794 (n8731, \b[4] , n7441);
  and g15800 (n8734, n394, n7449);
  not g15803 (n_7425, n8735);
  and g15804 (n8736, \a[47] , n_7425);
  not g15805 (n_7426, n8736);
  and g15806 (n8737, \a[47] , n_7426);
  and g15807 (n8738, n_7425, n_7426);
  not g15808 (n_7427, n8737);
  not g15809 (n_7428, n8738);
  and g15810 (n8739, n_7427, n_7428);
  not g15811 (n_7429, n8739);
  and g15812 (n8740, n8728, n_7429);
  not g15813 (n_7430, n8740);
  and g15814 (n8741, n8728, n_7430);
  and g15815 (n8742, n_7429, n_7430);
  not g15816 (n_7431, n8741);
  not g15817 (n_7432, n8742);
  and g15818 (n8743, n_7431, n_7432);
  not g15819 (n_7433, n8712);
  not g15820 (n_7434, n8743);
  and g15821 (n8744, n_7433, n_7434);
  and g15822 (n8745, n8712, n8743);
  not g15823 (n_7435, n8744);
  not g15824 (n_7436, n8745);
  and g15825 (n8746, n_7435, n_7436);
  not g15826 (n_7437, n8711);
  and g15827 (n8747, n_7437, n8746);
  not g15828 (n_7438, n8747);
  and g15829 (n8748, n_7437, n_7438);
  and g15830 (n8749, n8746, n_7438);
  not g15831 (n_7439, n8748);
  not g15832 (n_7440, n8749);
  and g15833 (n8750, n_7439, n_7440);
  not g15834 (n_7441, n8700);
  not g15835 (n_7442, n8750);
  and g15836 (n8751, n_7441, n_7442);
  not g15837 (n_7443, n8751);
  and g15838 (n8752, n_7441, n_7443);
  and g15839 (n8753, n_7442, n_7443);
  not g15840 (n_7444, n8752);
  not g15841 (n_7445, n8753);
  and g15842 (n8754, n_7444, n_7445);
  and g15843 (n8755, \b[11] , n5777);
  and g15844 (n8756, \b[9] , n6059);
  and g15845 (n8757, \b[10] , n5772);
  and g15851 (n8760, n818, n5780);
  not g15854 (n_7450, n8761);
  and g15855 (n8762, \a[41] , n_7450);
  not g15856 (n_7451, n8762);
  and g15857 (n8763, \a[41] , n_7451);
  and g15858 (n8764, n_7450, n_7451);
  not g15859 (n_7452, n8763);
  not g15860 (n_7453, n8764);
  and g15861 (n8765, n_7452, n_7453);
  and g15862 (n8766, n8754, n8765);
  not g15863 (n_7454, n8754);
  not g15864 (n_7455, n8765);
  and g15865 (n8767, n_7454, n_7455);
  not g15866 (n_7456, n8766);
  not g15867 (n_7457, n8767);
  and g15868 (n8768, n_7456, n_7457);
  not g15869 (n_7458, n8405);
  and g15870 (n8769, n_7458, n8768);
  not g15871 (n_7459, n8768);
  and g15872 (n8770, n8405, n_7459);
  not g15873 (n_7460, n8769);
  not g15874 (n_7461, n8770);
  and g15875 (n8771, n_7460, n_7461);
  not g15876 (n_7462, n8699);
  and g15877 (n8772, n_7462, n8771);
  not g15878 (n_7463, n8772);
  and g15879 (n8773, n8771, n_7463);
  and g15880 (n8774, n_7462, n_7463);
  not g15881 (n_7464, n8773);
  not g15882 (n_7465, n8774);
  and g15883 (n8775, n_7464, n_7465);
  not g15884 (n_7466, n8688);
  not g15885 (n_7467, n8775);
  and g15886 (n8776, n_7466, n_7467);
  and g15887 (n8777, n8688, n8775);
  not g15888 (n_7468, n8776);
  not g15889 (n_7469, n8777);
  and g15890 (n8778, n_7468, n_7469);
  not g15891 (n_7470, n8687);
  and g15892 (n8779, n_7470, n8778);
  not g15893 (n_7471, n8779);
  and g15894 (n8780, n_7470, n_7471);
  and g15895 (n8781, n8778, n_7471);
  not g15896 (n_7472, n8780);
  not g15897 (n_7473, n8781);
  and g15898 (n8782, n_7472, n_7473);
  not g15899 (n_7474, n8676);
  not g15900 (n_7475, n8782);
  and g15901 (n8783, n_7474, n_7475);
  not g15902 (n_7476, n8783);
  and g15903 (n8784, n_7474, n_7476);
  and g15904 (n8785, n_7475, n_7476);
  not g15905 (n_7477, n8784);
  not g15906 (n_7478, n8785);
  and g15907 (n8786, n_7477, n_7478);
  and g15908 (n8787, \b[20] , n3638);
  and g15909 (n8788, \b[18] , n3843);
  and g15910 (n8789, \b[19] , n3633);
  and g15916 (n8792, n1846, n3641);
  not g15919 (n_7483, n8793);
  and g15920 (n8794, \a[32] , n_7483);
  not g15921 (n_7484, n8794);
  and g15922 (n8795, \a[32] , n_7484);
  and g15923 (n8796, n_7483, n_7484);
  not g15924 (n_7485, n8795);
  not g15925 (n_7486, n8796);
  and g15926 (n8797, n_7485, n_7486);
  not g15927 (n_7487, n8786);
  not g15928 (n_7488, n8797);
  and g15929 (n8798, n_7487, n_7488);
  not g15930 (n_7489, n8798);
  and g15931 (n8799, n_7487, n_7489);
  and g15932 (n8800, n_7488, n_7489);
  not g15933 (n_7490, n8799);
  not g15934 (n_7491, n8800);
  and g15935 (n8801, n_7490, n_7491);
  and g15936 (n8802, n_7191, n_7197);
  and g15937 (n8803, n8801, n8802);
  not g15938 (n_7492, n8801);
  not g15939 (n_7493, n8802);
  and g15940 (n8804, n_7492, n_7493);
  not g15941 (n_7494, n8803);
  not g15942 (n_7495, n8804);
  and g15943 (n8805, n_7494, n_7495);
  and g15944 (n8806, \b[23] , n3050);
  and g15945 (n8807, \b[21] , n3243);
  and g15946 (n8808, \b[22] , n3045);
  and g15952 (n8811, n2300, n3053);
  not g15955 (n_7500, n8812);
  and g15956 (n8813, \a[29] , n_7500);
  not g15957 (n_7501, n8813);
  and g15958 (n8814, \a[29] , n_7501);
  and g15959 (n8815, n_7500, n_7501);
  not g15960 (n_7502, n8814);
  not g15961 (n_7503, n8815);
  and g15962 (n8816, n_7502, n_7503);
  not g15963 (n_7504, n8816);
  and g15964 (n8817, n8805, n_7504);
  not g15965 (n_7505, n8805);
  and g15966 (n8818, n_7505, n8816);
  not g15967 (n_7506, n8675);
  not g15968 (n_7507, n8818);
  and g15969 (n8819, n_7506, n_7507);
  not g15970 (n_7508, n8817);
  and g15971 (n8820, n_7508, n8819);
  not g15972 (n_7509, n8820);
  and g15973 (n8821, n_7506, n_7509);
  and g15974 (n8822, n_7508, n_7509);
  and g15975 (n8823, n_7507, n8822);
  not g15976 (n_7510, n8821);
  not g15977 (n_7511, n8823);
  and g15978 (n8824, n_7510, n_7511);
  and g15979 (n8825, \b[26] , n2539);
  and g15980 (n8826, \b[24] , n2685);
  and g15981 (n8827, \b[25] , n2534);
  and g15987 (n8830, n2542, n2813);
  not g15990 (n_7516, n8831);
  and g15991 (n8832, \a[26] , n_7516);
  not g15992 (n_7517, n8832);
  and g15993 (n8833, \a[26] , n_7517);
  and g15994 (n8834, n_7516, n_7517);
  not g15995 (n_7518, n8833);
  not g15996 (n_7519, n8834);
  and g15997 (n8835, n_7518, n_7519);
  and g15998 (n8836, n8824, n8835);
  not g15999 (n_7520, n8824);
  not g16000 (n_7521, n8835);
  and g16001 (n8837, n_7520, n_7521);
  not g16002 (n_7522, n8836);
  not g16003 (n_7523, n8837);
  and g16004 (n8838, n_7522, n_7523);
  not g16005 (n_7524, n8674);
  and g16006 (n8839, n_7524, n8838);
  not g16007 (n_7525, n8838);
  and g16008 (n8840, n8674, n_7525);
  not g16009 (n_7526, n8839);
  not g16010 (n_7527, n8840);
  and g16011 (n8841, n_7526, n_7527);
  not g16012 (n_7528, n8841);
  and g16013 (n8842, n8673, n_7528);
  not g16014 (n_7529, n8673);
  and g16015 (n8843, n_7529, n8841);
  not g16016 (n_7530, n8842);
  not g16017 (n_7531, n8843);
  and g16018 (n8844, n_7530, n_7531);
  not g16019 (n_7532, n8662);
  and g16020 (n8845, n_7532, n8844);
  not g16021 (n_7533, n8844);
  and g16022 (n8846, n8662, n_7533);
  not g16023 (n_7534, n8845);
  not g16024 (n_7535, n8846);
  and g16025 (n8847, n_7534, n_7535);
  not g16026 (n_7536, n8847);
  and g16027 (n8848, n8661, n_7536);
  not g16028 (n_7537, n8661);
  and g16029 (n8849, n_7537, n8847);
  not g16030 (n_7538, n8848);
  not g16031 (n_7539, n8849);
  and g16032 (n8850, n_7538, n_7539);
  not g16033 (n_7540, n8650);
  and g16034 (n8851, n_7540, n8850);
  not g16035 (n_7541, n8850);
  and g16036 (n8852, n8650, n_7541);
  not g16037 (n_7542, n8851);
  not g16038 (n_7543, n8852);
  and g16039 (n8853, n_7542, n_7543);
  not g16040 (n_7544, n8649);
  and g16041 (n8854, n_7544, n8853);
  not g16042 (n_7545, n8854);
  and g16043 (n8855, n8853, n_7545);
  and g16044 (n8856, n_7544, n_7545);
  not g16045 (n_7546, n8855);
  not g16046 (n_7547, n8856);
  and g16047 (n8857, n_7546, n_7547);
  and g16048 (n8858, n_7265, n_7272);
  and g16049 (n8859, n8857, n8858);
  not g16050 (n_7548, n8857);
  not g16051 (n_7549, n8858);
  and g16052 (n8860, n_7548, n_7549);
  not g16053 (n_7550, n8859);
  not g16054 (n_7551, n8860);
  and g16055 (n8861, n_7550, n_7551);
  and g16056 (n8862, \b[38] , n951);
  and g16057 (n8863, \b[36] , n1056);
  and g16058 (n8864, \b[37] , n946);
  and g16064 (n8867, n954, n5205);
  not g16067 (n_7556, n8868);
  and g16068 (n8869, \a[14] , n_7556);
  not g16069 (n_7557, n8869);
  and g16070 (n8870, \a[14] , n_7557);
  and g16071 (n8871, n_7556, n_7557);
  not g16072 (n_7558, n8870);
  not g16073 (n_7559, n8871);
  and g16074 (n8872, n_7558, n_7559);
  not g16075 (n_7560, n8872);
  and g16076 (n8873, n8861, n_7560);
  not g16077 (n_7561, n8873);
  and g16078 (n8874, n8861, n_7561);
  and g16079 (n8875, n_7560, n_7561);
  not g16080 (n_7562, n8874);
  not g16081 (n_7563, n8875);
  and g16082 (n8876, n_7562, n_7563);
  and g16083 (n8877, n_7282, n_7288);
  and g16084 (n8878, n8876, n8877);
  not g16085 (n_7564, n8876);
  not g16086 (n_7565, n8877);
  and g16087 (n8879, n_7564, n_7565);
  not g16088 (n_7566, n8878);
  not g16089 (n_7567, n8879);
  and g16090 (n8880, n_7566, n_7567);
  and g16091 (n8881, \b[41] , n700);
  and g16092 (n8882, \b[39] , n767);
  and g16093 (n8883, \b[40] , n695);
  and g16099 (n8886, n703, n6219);
  not g16102 (n_7572, n8887);
  and g16103 (n8888, \a[11] , n_7572);
  not g16104 (n_7573, n8888);
  and g16105 (n8889, \a[11] , n_7573);
  and g16106 (n8890, n_7572, n_7573);
  not g16107 (n_7574, n8889);
  not g16108 (n_7575, n8890);
  and g16109 (n8891, n_7574, n_7575);
  not g16110 (n_7576, n8891);
  and g16111 (n8892, n8880, n_7576);
  not g16112 (n_7577, n8892);
  and g16113 (n8893, n8880, n_7577);
  and g16114 (n8894, n_7576, n_7577);
  not g16115 (n_7578, n8893);
  not g16116 (n_7579, n8894);
  and g16117 (n8895, n_7578, n_7579);
  and g16118 (n8896, n_7298, n_7304);
  and g16119 (n8897, n8895, n8896);
  not g16120 (n_7580, n8895);
  not g16121 (n_7581, n8896);
  and g16122 (n8898, n_7580, n_7581);
  not g16123 (n_7582, n8897);
  not g16124 (n_7583, n8898);
  and g16125 (n8899, n_7582, n_7583);
  and g16126 (n8900, \b[44] , n511);
  and g16127 (n8901, \b[42] , n541);
  and g16128 (n8902, \b[43] , n506);
  and g16134 (n8905, n514, n7072);
  not g16137 (n_7588, n8906);
  and g16138 (n8907, \a[8] , n_7588);
  not g16139 (n_7589, n8907);
  and g16140 (n8908, \a[8] , n_7589);
  and g16141 (n8909, n_7588, n_7589);
  not g16142 (n_7590, n8908);
  not g16143 (n_7591, n8909);
  and g16144 (n8910, n_7590, n_7591);
  not g16145 (n_7592, n8910);
  and g16146 (n8911, n8899, n_7592);
  not g16147 (n_7593, n8899);
  and g16148 (n8912, n_7593, n8910);
  not g16149 (n_7594, n8638);
  not g16150 (n_7595, n8912);
  and g16151 (n8913, n_7594, n_7595);
  not g16152 (n_7596, n8911);
  and g16153 (n8914, n_7596, n8913);
  not g16154 (n_7597, n8914);
  and g16155 (n8915, n_7594, n_7597);
  and g16156 (n8916, n_7596, n_7597);
  and g16157 (n8917, n_7595, n8916);
  not g16158 (n_7598, n8915);
  not g16159 (n_7599, n8917);
  and g16160 (n8918, n_7598, n_7599);
  and g16161 (n8919, \b[47] , n362);
  and g16162 (n8920, \b[45] , n403);
  and g16163 (n8921, \b[46] , n357);
  and g16169 (n8924, n365, n7703);
  not g16172 (n_7604, n8925);
  and g16173 (n8926, \a[5] , n_7604);
  not g16174 (n_7605, n8926);
  and g16175 (n8927, \a[5] , n_7605);
  and g16176 (n8928, n_7604, n_7605);
  not g16177 (n_7606, n8927);
  not g16178 (n_7607, n8928);
  and g16179 (n8929, n_7606, n_7607);
  not g16180 (n_7608, n8918);
  not g16181 (n_7609, n8929);
  and g16182 (n8930, n_7608, n_7609);
  not g16183 (n_7610, n8930);
  and g16184 (n8931, n_7608, n_7610);
  and g16185 (n8932, n_7609, n_7610);
  not g16186 (n_7611, n8931);
  not g16187 (n_7612, n8932);
  and g16188 (n8933, n_7611, n_7612);
  and g16189 (n8934, n_7331, n_7337);
  and g16190 (n8935, n8933, n8934);
  not g16191 (n_7613, n8933);
  not g16192 (n_7614, n8934);
  and g16193 (n8936, n_7613, n_7614);
  not g16194 (n_7615, n8935);
  not g16195 (n_7616, n8936);
  and g16196 (n8937, n_7615, n_7616);
  and g16197 (n8938, \b[50] , n266);
  and g16198 (n8939, \b[48] , n284);
  and g16199 (n8940, \b[49] , n261);
  and g16205 (n8943, n_7344, n_7347);
  not g16206 (n_7621, \b[50] );
  and g16207 (n8944, n_7342, n_7621);
  and g16208 (n8945, \b[49] , \b[50] );
  not g16209 (n_7622, n8944);
  not g16210 (n_7623, n8945);
  and g16211 (n8946, n_7622, n_7623);
  not g16212 (n_7624, n8943);
  and g16213 (n8947, n_7624, n8946);
  not g16214 (n_7625, n8946);
  and g16215 (n8948, n8943, n_7625);
  not g16216 (n_7626, n8947);
  not g16217 (n_7627, n8948);
  and g16218 (n8949, n_7626, n_7627);
  and g16219 (n8950, n269, n8949);
  not g16222 (n_7629, n8951);
  and g16223 (n8952, \a[2] , n_7629);
  not g16224 (n_7630, n8952);
  and g16225 (n8953, \a[2] , n_7630);
  and g16226 (n8954, n_7629, n_7630);
  not g16227 (n_7631, n8953);
  not g16228 (n_7632, n8954);
  and g16229 (n8955, n_7631, n_7632);
  not g16230 (n_7633, n8955);
  and g16231 (n8956, n8937, n_7633);
  not g16232 (n_7634, n8956);
  and g16233 (n8957, n8937, n_7634);
  and g16234 (n8958, n_7633, n_7634);
  not g16235 (n_7635, n8957);
  not g16236 (n_7636, n8958);
  and g16237 (n8959, n_7635, n_7636);
  and g16238 (n8960, n_7357, n_7360);
  not g16239 (n_7637, n8959);
  not g16240 (n_7638, n8960);
  and g16241 (n8961, n_7637, n_7638);
  and g16242 (n8962, n8959, n8960);
  not g16243 (n_7639, n8961);
  not g16244 (n_7640, n8962);
  and g16245 (\f[50] , n_7639, n_7640);
  and g16246 (n8964, n_7634, n_7639);
  and g16247 (n8965, \b[51] , n266);
  and g16248 (n8966, \b[49] , n284);
  and g16249 (n8967, \b[50] , n261);
  and g16255 (n8970, n_7623, n_7626);
  not g16256 (n_7645, \b[51] );
  and g16257 (n8971, n_7621, n_7645);
  and g16258 (n8972, \b[50] , \b[51] );
  not g16259 (n_7646, n8971);
  not g16260 (n_7647, n8972);
  and g16261 (n8973, n_7646, n_7647);
  not g16262 (n_7648, n8970);
  and g16263 (n8974, n_7648, n8973);
  not g16264 (n_7649, n8973);
  and g16265 (n8975, n8970, n_7649);
  not g16266 (n_7650, n8974);
  not g16267 (n_7651, n8975);
  and g16268 (n8976, n_7650, n_7651);
  and g16269 (n8977, n269, n8976);
  not g16272 (n_7653, n8978);
  and g16273 (n8979, \a[2] , n_7653);
  not g16274 (n_7654, n8979);
  and g16275 (n8980, \a[2] , n_7654);
  and g16276 (n8981, n_7653, n_7654);
  not g16277 (n_7655, n8980);
  not g16278 (n_7656, n8981);
  and g16279 (n8982, n_7655, n_7656);
  and g16280 (n8983, n_7610, n_7616);
  and g16281 (n8984, \b[45] , n511);
  and g16282 (n8985, \b[43] , n541);
  and g16283 (n8986, \b[44] , n506);
  and g16289 (n8989, n514, n7361);
  not g16292 (n_7661, n8990);
  and g16293 (n8991, \a[8] , n_7661);
  not g16294 (n_7662, n8991);
  and g16295 (n8992, \a[8] , n_7662);
  and g16296 (n8993, n_7661, n_7662);
  not g16297 (n_7663, n8992);
  not g16298 (n_7664, n8993);
  and g16299 (n8994, n_7663, n_7664);
  and g16300 (n8995, n_7545, n_7551);
  and g16301 (n8996, n_7539, n_7542);
  and g16302 (n8997, \b[33] , n1627);
  and g16303 (n8998, \b[31] , n1763);
  and g16304 (n8999, \b[32] , n1622);
  and g16310 (n9002, n1630, n4223);
  not g16313 (n_7669, n9003);
  and g16314 (n9004, \a[20] , n_7669);
  not g16315 (n_7670, n9004);
  and g16316 (n9005, \a[20] , n_7670);
  and g16317 (n9006, n_7669, n_7670);
  not g16318 (n_7671, n9005);
  not g16319 (n_7672, n9006);
  and g16320 (n9007, n_7671, n_7672);
  and g16321 (n9008, n_7531, n_7534);
  and g16322 (n9009, n_7523, n_7526);
  and g16323 (n9010, \b[27] , n2539);
  and g16324 (n9011, \b[25] , n2685);
  and g16325 (n9012, \b[26] , n2534);
  and g16331 (n9015, n2542, n2990);
  not g16334 (n_7677, n9016);
  and g16335 (n9017, \a[26] , n_7677);
  not g16336 (n_7678, n9017);
  and g16337 (n9018, \a[26] , n_7678);
  and g16338 (n9019, n_7677, n_7678);
  not g16339 (n_7679, n9018);
  not g16340 (n_7680, n9019);
  and g16341 (n9020, n_7679, n_7680);
  and g16342 (n9021, n_7471, n_7476);
  and g16343 (n9022, \b[18] , n4287);
  and g16344 (n9023, \b[16] , n4532);
  and g16345 (n9024, \b[17] , n4282);
  and g16351 (n9027, n1566, n4290);
  not g16354 (n_7685, n9028);
  and g16355 (n9029, \a[35] , n_7685);
  not g16356 (n_7686, n9029);
  and g16357 (n9030, \a[35] , n_7686);
  and g16358 (n9031, n_7685, n_7686);
  not g16359 (n_7687, n9030);
  not g16360 (n_7688, n9031);
  and g16361 (n9032, n_7687, n_7688);
  and g16362 (n9033, n_7463, n_7468);
  and g16363 (n9034, \b[15] , n5035);
  and g16364 (n9035, \b[13] , n5277);
  and g16365 (n9036, \b[14] , n5030);
  and g16371 (n9039, n1131, n5038);
  not g16374 (n_7693, n9040);
  and g16375 (n9041, \a[38] , n_7693);
  not g16376 (n_7694, n9041);
  and g16377 (n9042, \a[38] , n_7694);
  and g16378 (n9043, n_7693, n_7694);
  not g16379 (n_7695, n9042);
  not g16380 (n_7696, n9043);
  and g16381 (n9044, n_7695, n_7696);
  and g16382 (n9045, n_7457, n_7460);
  and g16383 (n9046, \b[12] , n5777);
  and g16384 (n9047, \b[10] , n6059);
  and g16385 (n9048, \b[11] , n5772);
  and g16391 (n9051, n842, n5780);
  not g16394 (n_7701, n9052);
  and g16395 (n9053, \a[41] , n_7701);
  not g16396 (n_7702, n9053);
  and g16397 (n9054, \a[41] , n_7702);
  and g16398 (n9055, n_7701, n_7702);
  not g16399 (n_7703, n9054);
  not g16400 (n_7704, n9055);
  and g16401 (n9056, n_7703, n_7704);
  and g16402 (n9057, n_7438, n_7443);
  and g16403 (n9058, \b[6] , n7446);
  and g16404 (n9059, \b[4] , n7787);
  and g16405 (n9060, \b[5] , n7441);
  and g16411 (n9063, n459, n7449);
  not g16414 (n_7709, n9064);
  and g16415 (n9065, \a[47] , n_7709);
  not g16416 (n_7710, n9065);
  and g16417 (n9066, \a[47] , n_7710);
  and g16418 (n9067, n_7709, n_7710);
  not g16419 (n_7711, n9066);
  not g16420 (n_7712, n9067);
  and g16421 (n9068, n_7711, n_7712);
  not g16422 (n_7714, \a[51] );
  and g16423 (n9069, \a[50] , n_7714);
  and g16424 (n9070, n_7111, \a[51] );
  not g16425 (n_7715, n9069);
  not g16426 (n_7716, n9070);
  and g16427 (n9071, n_7715, n_7716);
  not g16428 (n_7717, n9071);
  and g16429 (n9072, \b[0] , n_7717);
  and g16430 (n9073, n_7420, n9072);
  not g16431 (n_7718, n9072);
  and g16432 (n9074, n8727, n_7718);
  not g16433 (n_7719, n9073);
  not g16434 (n_7720, n9074);
  and g16435 (n9075, n_7719, n_7720);
  and g16436 (n9076, \b[3] , n8362);
  and g16437 (n9077, \b[1] , n8715);
  and g16438 (n9078, \b[2] , n8357);
  and g16444 (n9081, n318, n8365);
  not g16447 (n_7725, n9082);
  and g16448 (n9083, \a[50] , n_7725);
  not g16449 (n_7726, n9083);
  and g16450 (n9084, \a[50] , n_7726);
  and g16451 (n9085, n_7725, n_7726);
  not g16452 (n_7727, n9084);
  not g16453 (n_7728, n9085);
  and g16454 (n9086, n_7727, n_7728);
  not g16455 (n_7729, n9075);
  not g16456 (n_7730, n9086);
  and g16457 (n9087, n_7729, n_7730);
  and g16458 (n9088, n9075, n9086);
  not g16459 (n_7731, n9087);
  not g16460 (n_7732, n9088);
  and g16461 (n9089, n_7731, n_7732);
  not g16462 (n_7733, n9068);
  and g16463 (n9090, n_7733, n9089);
  not g16464 (n_7734, n9090);
  and g16465 (n9091, n9089, n_7734);
  and g16466 (n9092, n_7733, n_7734);
  not g16467 (n_7735, n9091);
  not g16468 (n_7736, n9092);
  and g16469 (n9093, n_7735, n_7736);
  and g16470 (n9094, n_7430, n_7435);
  and g16471 (n9095, n9093, n9094);
  not g16472 (n_7737, n9093);
  not g16473 (n_7738, n9094);
  and g16474 (n9096, n_7737, n_7738);
  not g16475 (n_7739, n9095);
  not g16476 (n_7740, n9096);
  and g16477 (n9097, n_7739, n_7740);
  and g16478 (n9098, \b[9] , n6595);
  and g16479 (n9099, \b[7] , n6902);
  and g16480 (n9100, \b[8] , n6590);
  and g16486 (n9103, n651, n6598);
  not g16489 (n_7745, n9104);
  and g16490 (n9105, \a[44] , n_7745);
  not g16491 (n_7746, n9105);
  and g16492 (n9106, \a[44] , n_7746);
  and g16493 (n9107, n_7745, n_7746);
  not g16494 (n_7747, n9106);
  not g16495 (n_7748, n9107);
  and g16496 (n9108, n_7747, n_7748);
  not g16497 (n_7749, n9097);
  and g16498 (n9109, n_7749, n9108);
  not g16499 (n_7750, n9108);
  and g16500 (n9110, n9097, n_7750);
  not g16501 (n_7751, n9109);
  not g16502 (n_7752, n9110);
  and g16503 (n9111, n_7751, n_7752);
  not g16504 (n_7753, n9057);
  and g16505 (n9112, n_7753, n9111);
  not g16506 (n_7754, n9111);
  and g16507 (n9113, n9057, n_7754);
  not g16508 (n_7755, n9112);
  not g16509 (n_7756, n9113);
  and g16510 (n9114, n_7755, n_7756);
  not g16511 (n_7757, n9056);
  and g16512 (n9115, n_7757, n9114);
  not g16513 (n_7758, n9115);
  and g16514 (n9116, n_7757, n_7758);
  and g16515 (n9117, n9114, n_7758);
  not g16516 (n_7759, n9116);
  not g16517 (n_7760, n9117);
  and g16518 (n9118, n_7759, n_7760);
  not g16519 (n_7761, n9045);
  not g16520 (n_7762, n9118);
  and g16521 (n9119, n_7761, n_7762);
  and g16522 (n9120, n9045, n_7760);
  and g16523 (n9121, n_7759, n9120);
  not g16524 (n_7763, n9119);
  not g16525 (n_7764, n9121);
  and g16526 (n9122, n_7763, n_7764);
  not g16527 (n_7765, n9044);
  and g16528 (n9123, n_7765, n9122);
  not g16529 (n_7766, n9122);
  and g16530 (n9124, n9044, n_7766);
  not g16531 (n_7767, n9123);
  not g16532 (n_7768, n9124);
  and g16533 (n9125, n_7767, n_7768);
  not g16534 (n_7769, n9033);
  and g16535 (n9126, n_7769, n9125);
  not g16536 (n_7770, n9125);
  and g16537 (n9127, n9033, n_7770);
  not g16538 (n_7771, n9126);
  not g16539 (n_7772, n9127);
  and g16540 (n9128, n_7771, n_7772);
  not g16541 (n_7773, n9032);
  and g16542 (n9129, n_7773, n9128);
  not g16543 (n_7774, n9128);
  and g16544 (n9130, n9032, n_7774);
  not g16545 (n_7775, n9129);
  not g16546 (n_7776, n9130);
  and g16547 (n9131, n_7775, n_7776);
  not g16548 (n_7777, n9021);
  and g16549 (n9132, n_7777, n9131);
  not g16550 (n_7778, n9131);
  and g16551 (n9133, n9021, n_7778);
  not g16552 (n_7779, n9132);
  not g16553 (n_7780, n9133);
  and g16554 (n9134, n_7779, n_7780);
  and g16555 (n9135, \b[21] , n3638);
  and g16556 (n9136, \b[19] , n3843);
  and g16557 (n9137, \b[20] , n3633);
  and g16563 (n9140, n1984, n3641);
  not g16566 (n_7785, n9141);
  and g16567 (n9142, \a[32] , n_7785);
  not g16568 (n_7786, n9142);
  and g16569 (n9143, \a[32] , n_7786);
  and g16570 (n9144, n_7785, n_7786);
  not g16571 (n_7787, n9143);
  not g16572 (n_7788, n9144);
  and g16573 (n9145, n_7787, n_7788);
  not g16574 (n_7789, n9145);
  and g16575 (n9146, n9134, n_7789);
  not g16576 (n_7790, n9146);
  and g16577 (n9147, n9134, n_7790);
  and g16578 (n9148, n_7789, n_7790);
  not g16579 (n_7791, n9147);
  not g16580 (n_7792, n9148);
  and g16581 (n9149, n_7791, n_7792);
  and g16582 (n9150, n_7489, n_7495);
  and g16583 (n9151, n9149, n9150);
  not g16584 (n_7793, n9149);
  not g16585 (n_7794, n9150);
  and g16586 (n9152, n_7793, n_7794);
  not g16587 (n_7795, n9151);
  not g16588 (n_7796, n9152);
  and g16589 (n9153, n_7795, n_7796);
  and g16590 (n9154, \b[24] , n3050);
  and g16591 (n9155, \b[22] , n3243);
  and g16592 (n9156, \b[23] , n3045);
  and g16598 (n9159, n2458, n3053);
  not g16601 (n_7801, n9160);
  and g16602 (n9161, \a[29] , n_7801);
  not g16603 (n_7802, n9161);
  and g16604 (n9162, \a[29] , n_7802);
  and g16605 (n9163, n_7801, n_7802);
  not g16606 (n_7803, n9162);
  not g16607 (n_7804, n9163);
  and g16608 (n9164, n_7803, n_7804);
  not g16609 (n_7805, n9153);
  and g16610 (n9165, n_7805, n9164);
  not g16611 (n_7806, n9164);
  and g16612 (n9166, n9153, n_7806);
  not g16613 (n_7807, n9165);
  not g16614 (n_7808, n9166);
  and g16615 (n9167, n_7807, n_7808);
  not g16616 (n_7809, n8822);
  and g16617 (n9168, n_7809, n9167);
  not g16618 (n_7810, n9167);
  and g16619 (n9169, n8822, n_7810);
  not g16620 (n_7811, n9168);
  not g16621 (n_7812, n9169);
  and g16622 (n9170, n_7811, n_7812);
  not g16623 (n_7813, n9020);
  and g16624 (n9171, n_7813, n9170);
  not g16625 (n_7814, n9171);
  and g16626 (n9172, n9170, n_7814);
  and g16627 (n9173, n_7813, n_7814);
  not g16628 (n_7815, n9172);
  not g16629 (n_7816, n9173);
  and g16630 (n9174, n_7815, n_7816);
  not g16631 (n_7817, n9009);
  and g16632 (n9175, n_7817, n9174);
  not g16633 (n_7818, n9174);
  and g16634 (n9176, n9009, n_7818);
  not g16635 (n_7819, n9175);
  not g16636 (n_7820, n9176);
  and g16637 (n9177, n_7819, n_7820);
  and g16638 (n9178, \b[30] , n2048);
  and g16639 (n9179, \b[28] , n2198);
  and g16640 (n9180, \b[29] , n2043);
  and g16646 (n9183, n2051, n3577);
  not g16649 (n_7825, n9184);
  and g16650 (n9185, \a[23] , n_7825);
  not g16651 (n_7826, n9185);
  and g16652 (n9186, \a[23] , n_7826);
  and g16653 (n9187, n_7825, n_7826);
  not g16654 (n_7827, n9186);
  not g16655 (n_7828, n9187);
  and g16656 (n9188, n_7827, n_7828);
  not g16657 (n_7829, n9177);
  not g16658 (n_7830, n9188);
  and g16659 (n9189, n_7829, n_7830);
  and g16660 (n9190, n9177, n9188);
  not g16661 (n_7831, n9189);
  not g16662 (n_7832, n9190);
  and g16663 (n9191, n_7831, n_7832);
  not g16664 (n_7833, n9008);
  and g16665 (n9192, n_7833, n9191);
  not g16666 (n_7834, n9191);
  and g16667 (n9193, n9008, n_7834);
  not g16668 (n_7835, n9192);
  not g16669 (n_7836, n9193);
  and g16670 (n9194, n_7835, n_7836);
  not g16671 (n_7837, n9007);
  and g16672 (n9195, n_7837, n9194);
  not g16673 (n_7838, n9195);
  and g16674 (n9196, n9194, n_7838);
  and g16675 (n9197, n_7837, n_7838);
  not g16676 (n_7839, n9196);
  not g16677 (n_7840, n9197);
  and g16678 (n9198, n_7839, n_7840);
  not g16679 (n_7841, n8996);
  and g16680 (n9199, n_7841, n9198);
  not g16681 (n_7842, n9198);
  and g16682 (n9200, n8996, n_7842);
  not g16683 (n_7843, n9199);
  not g16684 (n_7844, n9200);
  and g16685 (n9201, n_7843, n_7844);
  and g16686 (n9202, \b[36] , n1302);
  and g16687 (n9203, \b[34] , n1391);
  and g16688 (n9204, \b[35] , n1297);
  and g16694 (n9207, n1305, n4922);
  not g16697 (n_7849, n9208);
  and g16698 (n9209, \a[17] , n_7849);
  not g16699 (n_7850, n9209);
  and g16700 (n9210, \a[17] , n_7850);
  and g16701 (n9211, n_7849, n_7850);
  not g16702 (n_7851, n9210);
  not g16703 (n_7852, n9211);
  and g16704 (n9212, n_7851, n_7852);
  not g16705 (n_7853, n9201);
  not g16706 (n_7854, n9212);
  and g16707 (n9213, n_7853, n_7854);
  and g16708 (n9214, n9201, n9212);
  not g16709 (n_7855, n9213);
  not g16710 (n_7856, n9214);
  and g16711 (n9215, n_7855, n_7856);
  not g16712 (n_7857, n9215);
  and g16713 (n9216, n8995, n_7857);
  not g16714 (n_7858, n8995);
  and g16715 (n9217, n_7858, n9215);
  not g16716 (n_7859, n9216);
  not g16717 (n_7860, n9217);
  and g16718 (n9218, n_7859, n_7860);
  and g16719 (n9219, \b[39] , n951);
  and g16720 (n9220, \b[37] , n1056);
  and g16721 (n9221, \b[38] , n946);
  and g16727 (n9224, n954, n5451);
  not g16730 (n_7865, n9225);
  and g16731 (n9226, \a[14] , n_7865);
  not g16732 (n_7866, n9226);
  and g16733 (n9227, \a[14] , n_7866);
  and g16734 (n9228, n_7865, n_7866);
  not g16735 (n_7867, n9227);
  not g16736 (n_7868, n9228);
  and g16737 (n9229, n_7867, n_7868);
  not g16738 (n_7869, n9229);
  and g16739 (n9230, n9218, n_7869);
  not g16740 (n_7870, n9230);
  and g16741 (n9231, n9218, n_7870);
  and g16742 (n9232, n_7869, n_7870);
  not g16743 (n_7871, n9231);
  not g16744 (n_7872, n9232);
  and g16745 (n9233, n_7871, n_7872);
  and g16746 (n9234, n_7561, n_7567);
  and g16747 (n9235, n9233, n9234);
  not g16748 (n_7873, n9233);
  not g16749 (n_7874, n9234);
  and g16750 (n9236, n_7873, n_7874);
  not g16751 (n_7875, n9235);
  not g16752 (n_7876, n9236);
  and g16753 (n9237, n_7875, n_7876);
  and g16754 (n9238, \b[42] , n700);
  and g16755 (n9239, \b[40] , n767);
  and g16756 (n9240, \b[41] , n695);
  and g16762 (n9243, n703, n6489);
  not g16765 (n_7881, n9244);
  and g16766 (n9245, \a[11] , n_7881);
  not g16767 (n_7882, n9245);
  and g16768 (n9246, \a[11] , n_7882);
  and g16769 (n9247, n_7881, n_7882);
  not g16770 (n_7883, n9246);
  not g16771 (n_7884, n9247);
  and g16772 (n9248, n_7883, n_7884);
  not g16773 (n_7885, n9237);
  and g16774 (n9249, n_7885, n9248);
  not g16775 (n_7886, n9248);
  and g16776 (n9250, n9237, n_7886);
  not g16777 (n_7887, n9249);
  not g16778 (n_7888, n9250);
  and g16779 (n9251, n_7887, n_7888);
  and g16780 (n9252, n_7577, n_7583);
  not g16781 (n_7889, n9252);
  and g16782 (n9253, n9251, n_7889);
  not g16783 (n_7890, n9251);
  and g16784 (n9254, n_7890, n9252);
  not g16785 (n_7891, n9253);
  not g16786 (n_7892, n9254);
  and g16787 (n9255, n_7891, n_7892);
  not g16788 (n_7893, n8994);
  and g16789 (n9256, n_7893, n9255);
  not g16790 (n_7894, n9256);
  and g16791 (n9257, n9255, n_7894);
  and g16792 (n9258, n_7893, n_7894);
  not g16793 (n_7895, n9257);
  not g16794 (n_7896, n9258);
  and g16795 (n9259, n_7895, n_7896);
  not g16796 (n_7897, n8916);
  and g16797 (n9260, n_7897, n9259);
  not g16798 (n_7898, n9259);
  and g16799 (n9261, n8916, n_7898);
  not g16800 (n_7899, n9260);
  not g16801 (n_7900, n9261);
  and g16802 (n9262, n_7899, n_7900);
  and g16803 (n9263, \b[48] , n362);
  and g16804 (n9264, \b[46] , n403);
  and g16805 (n9265, \b[47] , n357);
  and g16811 (n9268, n365, n8009);
  not g16814 (n_7905, n9269);
  and g16815 (n9270, \a[5] , n_7905);
  not g16816 (n_7906, n9270);
  and g16817 (n9271, \a[5] , n_7906);
  and g16818 (n9272, n_7905, n_7906);
  not g16819 (n_7907, n9271);
  not g16820 (n_7908, n9272);
  and g16821 (n9273, n_7907, n_7908);
  and g16822 (n9274, n9262, n9273);
  not g16823 (n_7909, n9262);
  not g16824 (n_7910, n9273);
  and g16825 (n9275, n_7909, n_7910);
  not g16826 (n_7911, n9274);
  not g16827 (n_7912, n9275);
  and g16828 (n9276, n_7911, n_7912);
  not g16829 (n_7913, n8983);
  and g16830 (n9277, n_7913, n9276);
  not g16831 (n_7914, n9276);
  and g16832 (n9278, n8983, n_7914);
  not g16833 (n_7915, n9277);
  not g16834 (n_7916, n9278);
  and g16835 (n9279, n_7915, n_7916);
  not g16836 (n_7917, n8982);
  and g16837 (n9280, n_7917, n9279);
  not g16838 (n_7918, n9279);
  and g16839 (n9281, n8982, n_7918);
  not g16840 (n_7919, n9280);
  not g16841 (n_7920, n9281);
  and g16842 (n9282, n_7919, n_7920);
  not g16843 (n_7921, n8964);
  and g16844 (n9283, n_7921, n9282);
  not g16845 (n_7922, n9282);
  and g16846 (n9284, n8964, n_7922);
  not g16847 (n_7923, n9283);
  not g16848 (n_7924, n9284);
  and g16849 (\f[51] , n_7923, n_7924);
  and g16850 (n9286, n_7919, n_7923);
  and g16851 (n9287, n_7912, n_7915);
  and g16852 (n9288, n_7888, n_7891);
  and g16853 (n9289, n_7817, n_7818);
  not g16854 (n_7925, n9289);
  and g16855 (n9290, n_7814, n_7925);
  and g16856 (n9291, n_7808, n_7811);
  and g16857 (n9292, n_7775, n_7779);
  and g16858 (n9293, \b[16] , n5035);
  and g16859 (n9294, \b[14] , n5277);
  and g16860 (n9295, \b[15] , n5030);
  and g16866 (n9298, n1237, n5038);
  not g16869 (n_7930, n9299);
  and g16870 (n9300, \a[38] , n_7930);
  not g16871 (n_7931, n9300);
  and g16872 (n9301, \a[38] , n_7931);
  and g16873 (n9302, n_7930, n_7931);
  not g16874 (n_7932, n9301);
  not g16875 (n_7933, n9302);
  and g16876 (n9303, n_7932, n_7933);
  and g16877 (n9304, n_7758, n_7763);
  and g16878 (n9305, n_7752, n_7755);
  and g16879 (n9306, \b[7] , n7446);
  and g16880 (n9307, \b[5] , n7787);
  and g16881 (n9308, \b[6] , n7441);
  and g16887 (n9311, n484, n7449);
  not g16890 (n_7938, n9312);
  and g16891 (n9313, \a[47] , n_7938);
  not g16892 (n_7939, n9313);
  and g16893 (n9314, \a[47] , n_7939);
  and g16894 (n9315, n_7938, n_7939);
  not g16895 (n_7940, n9314);
  not g16896 (n_7941, n9315);
  and g16897 (n9316, n_7940, n_7941);
  and g16898 (n9317, n8727, n9072);
  not g16899 (n_7942, n9317);
  and g16900 (n9318, n_7731, n_7942);
  and g16901 (n9319, \b[4] , n8362);
  and g16902 (n9320, \b[2] , n8715);
  and g16903 (n9321, \b[3] , n8357);
  and g16909 (n9324, n346, n8365);
  not g16912 (n_7947, n9325);
  and g16913 (n9326, \a[50] , n_7947);
  not g16914 (n_7948, n9326);
  and g16915 (n9327, \a[50] , n_7948);
  and g16916 (n9328, n_7947, n_7948);
  not g16917 (n_7949, n9327);
  not g16918 (n_7950, n9328);
  and g16919 (n9329, n_7949, n_7950);
  and g16920 (n9330, \a[53] , n_7718);
  and g16921 (n9331, n_7714, \a[52] );
  not g16922 (n_7953, \a[52] );
  and g16923 (n9332, \a[51] , n_7953);
  not g16924 (n_7954, n9331);
  not g16925 (n_7955, n9332);
  and g16926 (n9333, n_7954, n_7955);
  not g16927 (n_7956, n9333);
  and g16928 (n9334, n9071, n_7956);
  and g16929 (n9335, \b[0] , n9334);
  and g16930 (n9336, n_7953, \a[53] );
  not g16931 (n_7957, \a[53] );
  and g16932 (n9337, \a[52] , n_7957);
  not g16933 (n_7958, n9336);
  not g16934 (n_7959, n9337);
  and g16935 (n9338, n_7958, n_7959);
  and g16936 (n9339, n_7717, n9338);
  and g16937 (n9340, \b[1] , n9339);
  not g16938 (n_7960, n9335);
  not g16939 (n_7961, n9340);
  and g16940 (n9341, n_7960, n_7961);
  not g16941 (n_7962, n9338);
  and g16942 (n9342, n_7717, n_7962);
  and g16943 (n9343, n_21, n9342);
  not g16944 (n_7963, n9343);
  and g16945 (n9344, n9341, n_7963);
  not g16946 (n_7964, n9344);
  and g16947 (n9345, \a[53] , n_7964);
  not g16948 (n_7965, n9345);
  and g16949 (n9346, \a[53] , n_7965);
  and g16950 (n9347, n_7964, n_7965);
  not g16951 (n_7966, n9346);
  not g16952 (n_7967, n9347);
  and g16953 (n9348, n_7966, n_7967);
  not g16954 (n_7968, n9348);
  and g16955 (n9349, n9330, n_7968);
  not g16956 (n_7969, n9330);
  and g16957 (n9350, n_7969, n9348);
  not g16958 (n_7970, n9349);
  not g16959 (n_7971, n9350);
  and g16960 (n9351, n_7970, n_7971);
  not g16961 (n_7972, n9351);
  and g16962 (n9352, n9329, n_7972);
  not g16963 (n_7973, n9329);
  and g16964 (n9353, n_7973, n9351);
  not g16965 (n_7974, n9352);
  not g16966 (n_7975, n9353);
  and g16967 (n9354, n_7974, n_7975);
  not g16968 (n_7976, n9318);
  and g16969 (n9355, n_7976, n9354);
  not g16970 (n_7977, n9354);
  and g16971 (n9356, n9318, n_7977);
  not g16972 (n_7978, n9355);
  not g16973 (n_7979, n9356);
  and g16974 (n9357, n_7978, n_7979);
  not g16975 (n_7980, n9316);
  and g16976 (n9358, n_7980, n9357);
  not g16977 (n_7981, n9358);
  and g16978 (n9359, n9357, n_7981);
  and g16979 (n9360, n_7980, n_7981);
  not g16980 (n_7982, n9359);
  not g16981 (n_7983, n9360);
  and g16982 (n9361, n_7982, n_7983);
  and g16983 (n9362, n_7734, n_7740);
  and g16984 (n9363, n9361, n9362);
  not g16985 (n_7984, n9361);
  not g16986 (n_7985, n9362);
  and g16987 (n9364, n_7984, n_7985);
  not g16988 (n_7986, n9363);
  not g16989 (n_7987, n9364);
  and g16990 (n9365, n_7986, n_7987);
  and g16991 (n9366, \b[10] , n6595);
  and g16992 (n9367, \b[8] , n6902);
  and g16993 (n9368, \b[9] , n6590);
  and g16999 (n9371, n738, n6598);
  not g17002 (n_7992, n9372);
  and g17003 (n9373, \a[44] , n_7992);
  not g17004 (n_7993, n9373);
  and g17005 (n9374, \a[44] , n_7993);
  and g17006 (n9375, n_7992, n_7993);
  not g17007 (n_7994, n9374);
  not g17008 (n_7995, n9375);
  and g17009 (n9376, n_7994, n_7995);
  not g17010 (n_7996, n9376);
  and g17011 (n9377, n9365, n_7996);
  not g17012 (n_7997, n9365);
  and g17013 (n9378, n_7997, n9376);
  not g17014 (n_7998, n9305);
  not g17015 (n_7999, n9378);
  and g17016 (n9379, n_7998, n_7999);
  not g17017 (n_8000, n9377);
  and g17018 (n9380, n_8000, n9379);
  not g17019 (n_8001, n9380);
  and g17020 (n9381, n_7998, n_8001);
  and g17021 (n9382, n_8000, n_8001);
  and g17022 (n9383, n_7999, n9382);
  not g17023 (n_8002, n9381);
  not g17024 (n_8003, n9383);
  and g17025 (n9384, n_8002, n_8003);
  and g17026 (n9385, \b[13] , n5777);
  and g17027 (n9386, \b[11] , n6059);
  and g17028 (n9387, \b[12] , n5772);
  and g17034 (n9390, n1008, n5780);
  not g17037 (n_8008, n9391);
  and g17038 (n9392, \a[41] , n_8008);
  not g17039 (n_8009, n9392);
  and g17040 (n9393, \a[41] , n_8009);
  and g17041 (n9394, n_8008, n_8009);
  not g17042 (n_8010, n9393);
  not g17043 (n_8011, n9394);
  and g17044 (n9395, n_8010, n_8011);
  and g17045 (n9396, n9384, n9395);
  not g17046 (n_8012, n9384);
  not g17047 (n_8013, n9395);
  and g17048 (n9397, n_8012, n_8013);
  not g17049 (n_8014, n9396);
  not g17050 (n_8015, n9397);
  and g17051 (n9398, n_8014, n_8015);
  not g17052 (n_8016, n9304);
  and g17053 (n9399, n_8016, n9398);
  not g17054 (n_8017, n9398);
  and g17055 (n9400, n9304, n_8017);
  not g17056 (n_8018, n9399);
  not g17057 (n_8019, n9400);
  and g17058 (n9401, n_8018, n_8019);
  not g17059 (n_8020, n9303);
  and g17060 (n9402, n_8020, n9401);
  not g17061 (n_8021, n9402);
  and g17062 (n9403, n9401, n_8021);
  and g17063 (n9404, n_8020, n_8021);
  not g17064 (n_8022, n9403);
  not g17065 (n_8023, n9404);
  and g17066 (n9405, n_8022, n_8023);
  and g17067 (n9406, n_7767, n_7771);
  and g17068 (n9407, n9405, n9406);
  not g17069 (n_8024, n9405);
  not g17070 (n_8025, n9406);
  and g17071 (n9408, n_8024, n_8025);
  not g17072 (n_8026, n9407);
  not g17073 (n_8027, n9408);
  and g17074 (n9409, n_8026, n_8027);
  and g17075 (n9410, \b[19] , n4287);
  and g17076 (n9411, \b[17] , n4532);
  and g17077 (n9412, \b[18] , n4282);
  and g17083 (n9415, n1708, n4290);
  not g17086 (n_8032, n9416);
  and g17087 (n9417, \a[35] , n_8032);
  not g17088 (n_8033, n9417);
  and g17089 (n9418, \a[35] , n_8033);
  and g17090 (n9419, n_8032, n_8033);
  not g17091 (n_8034, n9418);
  not g17092 (n_8035, n9419);
  and g17093 (n9420, n_8034, n_8035);
  not g17094 (n_8036, n9420);
  and g17095 (n9421, n9409, n_8036);
  not g17096 (n_8037, n9409);
  and g17097 (n9422, n_8037, n9420);
  not g17098 (n_8038, n9292);
  not g17099 (n_8039, n9422);
  and g17100 (n9423, n_8038, n_8039);
  not g17101 (n_8040, n9421);
  and g17102 (n9424, n_8040, n9423);
  not g17103 (n_8041, n9424);
  and g17104 (n9425, n_8038, n_8041);
  and g17105 (n9426, n_8040, n_8041);
  and g17106 (n9427, n_8039, n9426);
  not g17107 (n_8042, n9425);
  not g17108 (n_8043, n9427);
  and g17109 (n9428, n_8042, n_8043);
  and g17110 (n9429, \b[22] , n3638);
  and g17111 (n9430, \b[20] , n3843);
  and g17112 (n9431, \b[21] , n3633);
  and g17118 (n9434, n2145, n3641);
  not g17121 (n_8048, n9435);
  and g17122 (n9436, \a[32] , n_8048);
  not g17123 (n_8049, n9436);
  and g17124 (n9437, \a[32] , n_8049);
  and g17125 (n9438, n_8048, n_8049);
  not g17126 (n_8050, n9437);
  not g17127 (n_8051, n9438);
  and g17128 (n9439, n_8050, n_8051);
  not g17129 (n_8052, n9428);
  not g17130 (n_8053, n9439);
  and g17131 (n9440, n_8052, n_8053);
  not g17132 (n_8054, n9440);
  and g17133 (n9441, n_8052, n_8054);
  and g17134 (n9442, n_8053, n_8054);
  not g17135 (n_8055, n9441);
  not g17136 (n_8056, n9442);
  and g17137 (n9443, n_8055, n_8056);
  and g17138 (n9444, n_7790, n_7796);
  and g17139 (n9445, n9443, n9444);
  not g17140 (n_8057, n9443);
  not g17141 (n_8058, n9444);
  and g17142 (n9446, n_8057, n_8058);
  not g17143 (n_8059, n9445);
  not g17144 (n_8060, n9446);
  and g17145 (n9447, n_8059, n_8060);
  and g17146 (n9448, \b[25] , n3050);
  and g17147 (n9449, \b[23] , n3243);
  and g17148 (n9450, \b[24] , n3045);
  and g17154 (n9453, n2485, n3053);
  not g17157 (n_8065, n9454);
  and g17158 (n9455, \a[29] , n_8065);
  not g17159 (n_8066, n9455);
  and g17160 (n9456, \a[29] , n_8066);
  and g17161 (n9457, n_8065, n_8066);
  not g17162 (n_8067, n9456);
  not g17163 (n_8068, n9457);
  and g17164 (n9458, n_8067, n_8068);
  not g17165 (n_8069, n9458);
  and g17166 (n9459, n9447, n_8069);
  not g17167 (n_8070, n9459);
  and g17168 (n9460, n9447, n_8070);
  and g17169 (n9461, n_8069, n_8070);
  not g17170 (n_8071, n9460);
  not g17171 (n_8072, n9461);
  and g17172 (n9462, n_8071, n_8072);
  not g17173 (n_8073, n9291);
  and g17174 (n9463, n_8073, n9462);
  not g17175 (n_8074, n9462);
  and g17176 (n9464, n9291, n_8074);
  not g17177 (n_8075, n9463);
  not g17178 (n_8076, n9464);
  and g17179 (n9465, n_8075, n_8076);
  and g17180 (n9466, \b[28] , n2539);
  and g17181 (n9467, \b[26] , n2685);
  and g17182 (n9468, \b[27] , n2534);
  and g17188 (n9471, n2542, n3189);
  not g17191 (n_8081, n9472);
  and g17192 (n9473, \a[26] , n_8081);
  not g17193 (n_8082, n9473);
  and g17194 (n9474, \a[26] , n_8082);
  and g17195 (n9475, n_8081, n_8082);
  not g17196 (n_8083, n9474);
  not g17197 (n_8084, n9475);
  and g17198 (n9476, n_8083, n_8084);
  not g17199 (n_8085, n9465);
  not g17200 (n_8086, n9476);
  and g17201 (n9477, n_8085, n_8086);
  and g17202 (n9478, n9465, n9476);
  not g17203 (n_8087, n9477);
  not g17204 (n_8088, n9478);
  and g17205 (n9479, n_8087, n_8088);
  not g17206 (n_8089, n9479);
  and g17207 (n9480, n9290, n_8089);
  not g17208 (n_8090, n9290);
  and g17209 (n9481, n_8090, n9479);
  not g17210 (n_8091, n9480);
  not g17211 (n_8092, n9481);
  and g17212 (n9482, n_8091, n_8092);
  and g17213 (n9483, \b[31] , n2048);
  and g17214 (n9484, \b[29] , n2198);
  and g17215 (n9485, \b[30] , n2043);
  and g17221 (n9488, n2051, n3796);
  not g17224 (n_8097, n9489);
  and g17225 (n9490, \a[23] , n_8097);
  not g17226 (n_8098, n9490);
  and g17227 (n9491, \a[23] , n_8098);
  and g17228 (n9492, n_8097, n_8098);
  not g17229 (n_8099, n9491);
  not g17230 (n_8100, n9492);
  and g17231 (n9493, n_8099, n_8100);
  not g17232 (n_8101, n9493);
  and g17233 (n9494, n9482, n_8101);
  not g17234 (n_8102, n9494);
  and g17235 (n9495, n9482, n_8102);
  and g17236 (n9496, n_8101, n_8102);
  not g17237 (n_8103, n9495);
  not g17238 (n_8104, n9496);
  and g17239 (n9497, n_8103, n_8104);
  and g17240 (n9498, n_7831, n_7835);
  and g17241 (n9499, n9497, n9498);
  not g17242 (n_8105, n9497);
  not g17243 (n_8106, n9498);
  and g17244 (n9500, n_8105, n_8106);
  not g17245 (n_8107, n9499);
  not g17246 (n_8108, n9500);
  and g17247 (n9501, n_8107, n_8108);
  and g17248 (n9502, \b[34] , n1627);
  and g17249 (n9503, \b[32] , n1763);
  and g17250 (n9504, \b[33] , n1622);
  and g17256 (n9507, n1630, n4466);
  not g17259 (n_8113, n9508);
  and g17260 (n9509, \a[20] , n_8113);
  not g17261 (n_8114, n9509);
  and g17262 (n9510, \a[20] , n_8114);
  and g17263 (n9511, n_8113, n_8114);
  not g17264 (n_8115, n9510);
  not g17265 (n_8116, n9511);
  and g17266 (n9512, n_8115, n_8116);
  not g17267 (n_8117, n9512);
  and g17268 (n9513, n9501, n_8117);
  not g17269 (n_8118, n9513);
  and g17270 (n9514, n9501, n_8118);
  and g17271 (n9515, n_8117, n_8118);
  not g17272 (n_8119, n9514);
  not g17273 (n_8120, n9515);
  and g17274 (n9516, n_8119, n_8120);
  and g17275 (n9517, n_7841, n_7842);
  not g17276 (n_8121, n9517);
  and g17277 (n9518, n_7838, n_8121);
  and g17278 (n9519, n9516, n9518);
  not g17279 (n_8122, n9516);
  not g17280 (n_8123, n9518);
  and g17281 (n9520, n_8122, n_8123);
  not g17282 (n_8124, n9519);
  not g17283 (n_8125, n9520);
  and g17284 (n9521, n_8124, n_8125);
  and g17285 (n9522, \b[37] , n1302);
  and g17286 (n9523, \b[35] , n1391);
  and g17287 (n9524, \b[36] , n1297);
  and g17293 (n9527, n1305, n5181);
  not g17296 (n_8130, n9528);
  and g17297 (n9529, \a[17] , n_8130);
  not g17298 (n_8131, n9529);
  and g17299 (n9530, \a[17] , n_8131);
  and g17300 (n9531, n_8130, n_8131);
  not g17301 (n_8132, n9530);
  not g17302 (n_8133, n9531);
  and g17303 (n9532, n_8132, n_8133);
  not g17304 (n_8134, n9532);
  and g17305 (n9533, n9521, n_8134);
  not g17306 (n_8135, n9533);
  and g17307 (n9534, n9521, n_8135);
  and g17308 (n9535, n_8134, n_8135);
  not g17309 (n_8136, n9534);
  not g17310 (n_8137, n9535);
  and g17311 (n9536, n_8136, n_8137);
  and g17312 (n9537, n_7855, n_7860);
  and g17313 (n9538, n9536, n9537);
  not g17314 (n_8138, n9536);
  not g17315 (n_8139, n9537);
  and g17316 (n9539, n_8138, n_8139);
  not g17317 (n_8140, n9538);
  not g17318 (n_8141, n9539);
  and g17319 (n9540, n_8140, n_8141);
  and g17320 (n9541, \b[40] , n951);
  and g17321 (n9542, \b[38] , n1056);
  and g17322 (n9543, \b[39] , n946);
  and g17328 (n9546, n954, n5955);
  not g17331 (n_8146, n9547);
  and g17332 (n9548, \a[14] , n_8146);
  not g17333 (n_8147, n9548);
  and g17334 (n9549, \a[14] , n_8147);
  and g17335 (n9550, n_8146, n_8147);
  not g17336 (n_8148, n9549);
  not g17337 (n_8149, n9550);
  and g17338 (n9551, n_8148, n_8149);
  not g17339 (n_8150, n9551);
  and g17340 (n9552, n9540, n_8150);
  not g17341 (n_8151, n9552);
  and g17342 (n9553, n9540, n_8151);
  and g17343 (n9554, n_8150, n_8151);
  not g17344 (n_8152, n9553);
  not g17345 (n_8153, n9554);
  and g17346 (n9555, n_8152, n_8153);
  and g17347 (n9556, n_7870, n_7876);
  and g17348 (n9557, n9555, n9556);
  not g17349 (n_8154, n9555);
  not g17350 (n_8155, n9556);
  and g17351 (n9558, n_8154, n_8155);
  not g17352 (n_8156, n9557);
  not g17353 (n_8157, n9558);
  and g17354 (n9559, n_8156, n_8157);
  and g17355 (n9560, \b[43] , n700);
  and g17356 (n9561, \b[41] , n767);
  and g17357 (n9562, \b[42] , n695);
  and g17363 (n9565, n703, n6515);
  not g17366 (n_8162, n9566);
  and g17367 (n9567, \a[11] , n_8162);
  not g17368 (n_8163, n9567);
  and g17369 (n9568, \a[11] , n_8163);
  and g17370 (n9569, n_8162, n_8163);
  not g17371 (n_8164, n9568);
  not g17372 (n_8165, n9569);
  and g17373 (n9570, n_8164, n_8165);
  not g17374 (n_8166, n9570);
  and g17375 (n9571, n9559, n_8166);
  not g17376 (n_8167, n9559);
  and g17377 (n9572, n_8167, n9570);
  not g17378 (n_8168, n9288);
  not g17379 (n_8169, n9572);
  and g17380 (n9573, n_8168, n_8169);
  not g17381 (n_8170, n9571);
  and g17382 (n9574, n_8170, n9573);
  not g17383 (n_8171, n9574);
  and g17384 (n9575, n_8168, n_8171);
  and g17385 (n9576, n_8170, n_8171);
  and g17386 (n9577, n_8169, n9576);
  not g17387 (n_8172, n9575);
  not g17388 (n_8173, n9577);
  and g17389 (n9578, n_8172, n_8173);
  and g17390 (n9579, \b[46] , n511);
  and g17391 (n9580, \b[44] , n541);
  and g17392 (n9581, \b[45] , n506);
  and g17398 (n9584, n514, n7677);
  not g17401 (n_8178, n9585);
  and g17402 (n9586, \a[8] , n_8178);
  not g17403 (n_8179, n9586);
  and g17404 (n9587, \a[8] , n_8179);
  and g17405 (n9588, n_8178, n_8179);
  not g17406 (n_8180, n9587);
  not g17407 (n_8181, n9588);
  and g17408 (n9589, n_8180, n_8181);
  not g17409 (n_8182, n9578);
  not g17410 (n_8183, n9589);
  and g17411 (n9590, n_8182, n_8183);
  not g17412 (n_8184, n9590);
  and g17413 (n9591, n_8182, n_8184);
  and g17414 (n9592, n_8183, n_8184);
  not g17415 (n_8185, n9591);
  not g17416 (n_8186, n9592);
  and g17417 (n9593, n_8185, n_8186);
  and g17418 (n9594, n_7897, n_7898);
  not g17419 (n_8187, n9594);
  and g17420 (n9595, n_7894, n_8187);
  and g17421 (n9596, n9593, n9595);
  not g17422 (n_8188, n9593);
  not g17423 (n_8189, n9595);
  and g17424 (n9597, n_8188, n_8189);
  not g17425 (n_8190, n9596);
  not g17426 (n_8191, n9597);
  and g17427 (n9598, n_8190, n_8191);
  and g17428 (n9599, \b[49] , n362);
  and g17429 (n9600, \b[47] , n403);
  and g17430 (n9601, \b[48] , n357);
  and g17436 (n9604, n365, n8625);
  not g17439 (n_8196, n9605);
  and g17440 (n9606, \a[5] , n_8196);
  not g17441 (n_8197, n9606);
  and g17442 (n9607, \a[5] , n_8197);
  and g17443 (n9608, n_8196, n_8197);
  not g17444 (n_8198, n9607);
  not g17445 (n_8199, n9608);
  and g17446 (n9609, n_8198, n_8199);
  not g17447 (n_8200, n9609);
  and g17448 (n9610, n9598, n_8200);
  not g17449 (n_8201, n9610);
  and g17450 (n9611, n9598, n_8201);
  and g17451 (n9612, n_8200, n_8201);
  not g17452 (n_8202, n9611);
  not g17453 (n_8203, n9612);
  and g17454 (n9613, n_8202, n_8203);
  not g17455 (n_8204, n9287);
  and g17456 (n9614, n_8204, n9613);
  not g17457 (n_8205, n9613);
  and g17458 (n9615, n9287, n_8205);
  not g17459 (n_8206, n9614);
  not g17460 (n_8207, n9615);
  and g17461 (n9616, n_8206, n_8207);
  and g17462 (n9617, \b[52] , n266);
  and g17463 (n9618, \b[50] , n284);
  and g17464 (n9619, \b[51] , n261);
  and g17470 (n9622, n_7647, n_7650);
  not g17471 (n_8212, \b[52] );
  and g17472 (n9623, n_7645, n_8212);
  and g17473 (n9624, \b[51] , \b[52] );
  not g17474 (n_8213, n9623);
  not g17475 (n_8214, n9624);
  and g17476 (n9625, n_8213, n_8214);
  not g17477 (n_8215, n9622);
  and g17478 (n9626, n_8215, n9625);
  not g17479 (n_8216, n9625);
  and g17480 (n9627, n9622, n_8216);
  not g17481 (n_8217, n9626);
  not g17482 (n_8218, n9627);
  and g17483 (n9628, n_8217, n_8218);
  and g17484 (n9629, n269, n9628);
  not g17487 (n_8220, n9630);
  and g17488 (n9631, \a[2] , n_8220);
  not g17489 (n_8221, n9631);
  and g17490 (n9632, \a[2] , n_8221);
  and g17491 (n9633, n_8220, n_8221);
  not g17492 (n_8222, n9632);
  not g17493 (n_8223, n9633);
  and g17494 (n9634, n_8222, n_8223);
  not g17495 (n_8224, n9616);
  not g17496 (n_8225, n9634);
  and g17497 (n9635, n_8224, n_8225);
  and g17498 (n9636, n9616, n9634);
  not g17499 (n_8226, n9635);
  not g17500 (n_8227, n9636);
  and g17501 (n9637, n_8226, n_8227);
  not g17502 (n_8228, n9286);
  and g17503 (n9638, n_8228, n9637);
  not g17504 (n_8229, n9637);
  and g17505 (n9639, n9286, n_8229);
  not g17506 (n_8230, n9638);
  not g17507 (n_8231, n9639);
  and g17508 (\f[52] , n_8230, n_8231);
  and g17509 (n9641, n_8226, n_8230);
  and g17510 (n9642, n_8204, n_8205);
  not g17511 (n_8232, n9642);
  and g17512 (n9643, n_8201, n_8232);
  and g17513 (n9644, \b[35] , n1627);
  and g17514 (n9645, \b[33] , n1763);
  and g17515 (n9646, \b[34] , n1622);
  and g17521 (n9649, n1630, n4696);
  not g17524 (n_8237, n9650);
  and g17525 (n9651, \a[20] , n_8237);
  not g17526 (n_8238, n9651);
  and g17527 (n9652, \a[20] , n_8238);
  and g17528 (n9653, n_8237, n_8238);
  not g17529 (n_8239, n9652);
  not g17530 (n_8240, n9653);
  and g17531 (n9654, n_8239, n_8240);
  and g17532 (n9655, n_8102, n_8108);
  and g17533 (n9656, \b[32] , n2048);
  and g17534 (n9657, \b[30] , n2198);
  and g17535 (n9658, \b[31] , n2043);
  and g17541 (n9661, n2051, n4013);
  not g17544 (n_8245, n9662);
  and g17545 (n9663, \a[23] , n_8245);
  not g17546 (n_8246, n9663);
  and g17547 (n9664, \a[23] , n_8246);
  and g17548 (n9665, n_8245, n_8246);
  not g17549 (n_8247, n9664);
  not g17550 (n_8248, n9665);
  and g17551 (n9666, n_8247, n_8248);
  and g17552 (n9667, n_8087, n_8092);
  and g17553 (n9668, \b[29] , n2539);
  and g17554 (n9669, \b[27] , n2685);
  and g17555 (n9670, \b[28] , n2534);
  and g17561 (n9673, n2542, n3383);
  not g17564 (n_8253, n9674);
  and g17565 (n9675, \a[26] , n_8253);
  not g17566 (n_8254, n9675);
  and g17567 (n9676, \a[26] , n_8254);
  and g17568 (n9677, n_8253, n_8254);
  not g17569 (n_8255, n9676);
  not g17570 (n_8256, n9677);
  and g17571 (n9678, n_8255, n_8256);
  and g17572 (n9679, n_8073, n_8074);
  not g17573 (n_8257, n9679);
  and g17574 (n9680, n_8070, n_8257);
  and g17575 (n9681, n_8054, n_8060);
  and g17576 (n9682, \b[23] , n3638);
  and g17577 (n9683, \b[21] , n3843);
  and g17578 (n9684, \b[22] , n3633);
  and g17584 (n9687, n2300, n3641);
  not g17587 (n_8262, n9688);
  and g17588 (n9689, \a[32] , n_8262);
  not g17589 (n_8263, n9689);
  and g17590 (n9690, \a[32] , n_8263);
  and g17591 (n9691, n_8262, n_8263);
  not g17592 (n_8264, n9690);
  not g17593 (n_8265, n9691);
  and g17594 (n9692, n_8264, n_8265);
  and g17595 (n9693, n_8021, n_8027);
  and g17596 (n9694, \b[17] , n5035);
  and g17597 (n9695, \b[15] , n5277);
  and g17598 (n9696, \b[16] , n5030);
  and g17604 (n9699, n1356, n5038);
  not g17607 (n_8270, n9700);
  and g17608 (n9701, \a[38] , n_8270);
  not g17609 (n_8271, n9701);
  and g17610 (n9702, \a[38] , n_8271);
  and g17611 (n9703, n_8270, n_8271);
  not g17612 (n_8272, n9702);
  not g17613 (n_8273, n9703);
  and g17614 (n9704, n_8272, n_8273);
  and g17615 (n9705, n_8015, n_8018);
  and g17616 (n9706, \b[14] , n5777);
  and g17617 (n9707, \b[12] , n6059);
  and g17618 (n9708, \b[13] , n5772);
  and g17624 (n9711, n1034, n5780);
  not g17627 (n_8278, n9712);
  and g17628 (n9713, \a[41] , n_8278);
  not g17629 (n_8279, n9713);
  and g17630 (n9714, \a[41] , n_8279);
  and g17631 (n9715, n_8278, n_8279);
  not g17632 (n_8280, n9714);
  not g17633 (n_8281, n9715);
  and g17634 (n9716, n_8280, n_8281);
  and g17635 (n9717, \b[11] , n6595);
  and g17636 (n9718, \b[9] , n6902);
  and g17637 (n9719, \b[10] , n6590);
  and g17643 (n9722, n818, n6598);
  not g17646 (n_8286, n9723);
  and g17647 (n9724, \a[44] , n_8286);
  not g17648 (n_8287, n9724);
  and g17649 (n9725, \a[44] , n_8287);
  and g17650 (n9726, n_8286, n_8287);
  not g17651 (n_8288, n9725);
  not g17652 (n_8289, n9726);
  and g17653 (n9727, n_8288, n_8289);
  and g17654 (n9728, n_7981, n_7987);
  and g17655 (n9729, n_7975, n_7978);
  and g17656 (n9730, \b[2] , n9339);
  and g17657 (n9731, n9071, n_7962);
  and g17658 (n9732, n9333, n9731);
  and g17659 (n9733, \b[0] , n9732);
  and g17660 (n9734, \b[1] , n9334);
  and g17666 (n9737, n296, n9342);
  not g17669 (n_8294, n9738);
  and g17670 (n9739, \a[53] , n_8294);
  not g17671 (n_8295, n9739);
  and g17672 (n9740, \a[53] , n_8295);
  and g17673 (n9741, n_8294, n_8295);
  not g17674 (n_8296, n9740);
  not g17675 (n_8297, n9741);
  and g17676 (n9742, n_8296, n_8297);
  and g17677 (n9743, n_7970, n9742);
  not g17678 (n_8298, n9742);
  and g17679 (n9744, n9349, n_8298);
  not g17680 (n_8299, n9743);
  not g17681 (n_8300, n9744);
  and g17682 (n9745, n_8299, n_8300);
  and g17683 (n9746, \b[5] , n8362);
  and g17684 (n9747, \b[3] , n8715);
  and g17685 (n9748, \b[4] , n8357);
  and g17691 (n9751, n394, n8365);
  not g17694 (n_8305, n9752);
  and g17695 (n9753, \a[50] , n_8305);
  not g17696 (n_8306, n9753);
  and g17697 (n9754, \a[50] , n_8306);
  and g17698 (n9755, n_8305, n_8306);
  not g17699 (n_8307, n9754);
  not g17700 (n_8308, n9755);
  and g17701 (n9756, n_8307, n_8308);
  not g17702 (n_8309, n9756);
  and g17703 (n9757, n9745, n_8309);
  not g17704 (n_8310, n9745);
  and g17705 (n9758, n_8310, n9756);
  not g17706 (n_8311, n9729);
  not g17707 (n_8312, n9758);
  and g17708 (n9759, n_8311, n_8312);
  not g17709 (n_8313, n9757);
  and g17710 (n9760, n_8313, n9759);
  not g17711 (n_8314, n9760);
  and g17712 (n9761, n_8311, n_8314);
  and g17713 (n9762, n_8313, n_8314);
  and g17714 (n9763, n_8312, n9762);
  not g17715 (n_8315, n9761);
  not g17716 (n_8316, n9763);
  and g17717 (n9764, n_8315, n_8316);
  and g17718 (n9765, \b[8] , n7446);
  and g17719 (n9766, \b[6] , n7787);
  and g17720 (n9767, \b[7] , n7441);
  and g17726 (n9770, n585, n7449);
  not g17729 (n_8321, n9771);
  and g17730 (n9772, \a[47] , n_8321);
  not g17731 (n_8322, n9772);
  and g17732 (n9773, \a[47] , n_8322);
  and g17733 (n9774, n_8321, n_8322);
  not g17734 (n_8323, n9773);
  not g17735 (n_8324, n9774);
  and g17736 (n9775, n_8323, n_8324);
  and g17737 (n9776, n9764, n9775);
  not g17738 (n_8325, n9764);
  not g17739 (n_8326, n9775);
  and g17740 (n9777, n_8325, n_8326);
  not g17741 (n_8327, n9776);
  not g17742 (n_8328, n9777);
  and g17743 (n9778, n_8327, n_8328);
  not g17744 (n_8329, n9728);
  and g17745 (n9779, n_8329, n9778);
  not g17746 (n_8330, n9778);
  and g17747 (n9780, n9728, n_8330);
  not g17748 (n_8331, n9779);
  not g17749 (n_8332, n9780);
  and g17750 (n9781, n_8331, n_8332);
  not g17751 (n_8333, n9781);
  and g17752 (n9782, n9727, n_8333);
  not g17753 (n_8334, n9727);
  and g17754 (n9783, n_8334, n9781);
  not g17755 (n_8335, n9782);
  not g17756 (n_8336, n9783);
  and g17757 (n9784, n_8335, n_8336);
  not g17758 (n_8337, n9382);
  and g17759 (n9785, n_8337, n9784);
  not g17760 (n_8338, n9784);
  and g17761 (n9786, n9382, n_8338);
  not g17762 (n_8339, n9785);
  not g17763 (n_8340, n9786);
  and g17764 (n9787, n_8339, n_8340);
  not g17765 (n_8341, n9716);
  and g17766 (n9788, n_8341, n9787);
  not g17767 (n_8342, n9788);
  and g17768 (n9789, n9787, n_8342);
  and g17769 (n9790, n_8341, n_8342);
  not g17770 (n_8343, n9789);
  not g17771 (n_8344, n9790);
  and g17772 (n9791, n_8343, n_8344);
  not g17773 (n_8345, n9705);
  not g17774 (n_8346, n9791);
  and g17775 (n9792, n_8345, n_8346);
  and g17776 (n9793, n9705, n9791);
  not g17777 (n_8347, n9792);
  not g17778 (n_8348, n9793);
  and g17779 (n9794, n_8347, n_8348);
  not g17780 (n_8349, n9704);
  and g17781 (n9795, n_8349, n9794);
  not g17782 (n_8350, n9795);
  and g17783 (n9796, n_8349, n_8350);
  and g17784 (n9797, n9794, n_8350);
  not g17785 (n_8351, n9796);
  not g17786 (n_8352, n9797);
  and g17787 (n9798, n_8351, n_8352);
  not g17788 (n_8353, n9693);
  not g17789 (n_8354, n9798);
  and g17790 (n9799, n_8353, n_8354);
  not g17791 (n_8355, n9799);
  and g17792 (n9800, n_8353, n_8355);
  and g17793 (n9801, n_8354, n_8355);
  not g17794 (n_8356, n9800);
  not g17795 (n_8357, n9801);
  and g17796 (n9802, n_8356, n_8357);
  and g17797 (n9803, \b[20] , n4287);
  and g17798 (n9804, \b[18] , n4532);
  and g17799 (n9805, \b[19] , n4282);
  and g17805 (n9808, n1846, n4290);
  not g17808 (n_8362, n9809);
  and g17809 (n9810, \a[35] , n_8362);
  not g17810 (n_8363, n9810);
  and g17811 (n9811, \a[35] , n_8363);
  and g17812 (n9812, n_8362, n_8363);
  not g17813 (n_8364, n9811);
  not g17814 (n_8365, n9812);
  and g17815 (n9813, n_8364, n_8365);
  not g17816 (n_8366, n9802);
  not g17817 (n_8367, n9813);
  and g17818 (n9814, n_8366, n_8367);
  not g17819 (n_8368, n9814);
  and g17820 (n9815, n_8366, n_8368);
  and g17821 (n9816, n_8367, n_8368);
  not g17822 (n_8369, n9815);
  not g17823 (n_8370, n9816);
  and g17824 (n9817, n_8369, n_8370);
  not g17825 (n_8371, n9426);
  not g17826 (n_8372, n9817);
  and g17827 (n9818, n_8371, n_8372);
  and g17828 (n9819, n9426, n9817);
  not g17829 (n_8373, n9818);
  not g17830 (n_8374, n9819);
  and g17831 (n9820, n_8373, n_8374);
  not g17832 (n_8375, n9692);
  and g17833 (n9821, n_8375, n9820);
  not g17834 (n_8376, n9821);
  and g17835 (n9822, n_8375, n_8376);
  and g17836 (n9823, n9820, n_8376);
  not g17837 (n_8377, n9822);
  not g17838 (n_8378, n9823);
  and g17839 (n9824, n_8377, n_8378);
  not g17840 (n_8379, n9681);
  not g17841 (n_8380, n9824);
  and g17842 (n9825, n_8379, n_8380);
  not g17843 (n_8381, n9825);
  and g17844 (n9826, n_8379, n_8381);
  and g17845 (n9827, n_8380, n_8381);
  not g17846 (n_8382, n9826);
  not g17847 (n_8383, n9827);
  and g17848 (n9828, n_8382, n_8383);
  and g17849 (n9829, \b[26] , n3050);
  and g17850 (n9830, \b[24] , n3243);
  and g17851 (n9831, \b[25] , n3045);
  and g17857 (n9834, n2813, n3053);
  not g17860 (n_8388, n9835);
  and g17861 (n9836, \a[29] , n_8388);
  not g17862 (n_8389, n9836);
  and g17863 (n9837, \a[29] , n_8389);
  and g17864 (n9838, n_8388, n_8389);
  not g17865 (n_8390, n9837);
  not g17866 (n_8391, n9838);
  and g17867 (n9839, n_8390, n_8391);
  and g17868 (n9840, n9828, n9839);
  not g17869 (n_8392, n9828);
  not g17870 (n_8393, n9839);
  and g17871 (n9841, n_8392, n_8393);
  not g17872 (n_8394, n9840);
  not g17873 (n_8395, n9841);
  and g17874 (n9842, n_8394, n_8395);
  not g17875 (n_8396, n9680);
  and g17876 (n9843, n_8396, n9842);
  not g17877 (n_8397, n9842);
  and g17878 (n9844, n9680, n_8397);
  not g17879 (n_8398, n9843);
  not g17880 (n_8399, n9844);
  and g17881 (n9845, n_8398, n_8399);
  not g17882 (n_8400, n9845);
  and g17883 (n9846, n9678, n_8400);
  not g17884 (n_8401, n9678);
  and g17885 (n9847, n_8401, n9845);
  not g17886 (n_8402, n9846);
  not g17887 (n_8403, n9847);
  and g17888 (n9848, n_8402, n_8403);
  not g17889 (n_8404, n9667);
  and g17890 (n9849, n_8404, n9848);
  not g17891 (n_8405, n9848);
  and g17892 (n9850, n9667, n_8405);
  not g17893 (n_8406, n9849);
  not g17894 (n_8407, n9850);
  and g17895 (n9851, n_8406, n_8407);
  not g17896 (n_8408, n9851);
  and g17897 (n9852, n9666, n_8408);
  not g17898 (n_8409, n9666);
  and g17899 (n9853, n_8409, n9851);
  not g17900 (n_8410, n9852);
  not g17901 (n_8411, n9853);
  and g17902 (n9854, n_8410, n_8411);
  not g17903 (n_8412, n9655);
  and g17904 (n9855, n_8412, n9854);
  not g17905 (n_8413, n9854);
  and g17906 (n9856, n9655, n_8413);
  not g17907 (n_8414, n9855);
  not g17908 (n_8415, n9856);
  and g17909 (n9857, n_8414, n_8415);
  not g17910 (n_8416, n9654);
  and g17911 (n9858, n_8416, n9857);
  not g17912 (n_8417, n9858);
  and g17913 (n9859, n9857, n_8417);
  and g17914 (n9860, n_8416, n_8417);
  not g17915 (n_8418, n9859);
  not g17916 (n_8419, n9860);
  and g17917 (n9861, n_8418, n_8419);
  and g17918 (n9862, n_8118, n_8125);
  and g17919 (n9863, n9861, n9862);
  not g17920 (n_8420, n9861);
  not g17921 (n_8421, n9862);
  and g17922 (n9864, n_8420, n_8421);
  not g17923 (n_8422, n9863);
  not g17924 (n_8423, n9864);
  and g17925 (n9865, n_8422, n_8423);
  and g17926 (n9866, \b[38] , n1302);
  and g17927 (n9867, \b[36] , n1391);
  and g17928 (n9868, \b[37] , n1297);
  and g17934 (n9871, n1305, n5205);
  not g17937 (n_8428, n9872);
  and g17938 (n9873, \a[17] , n_8428);
  not g17939 (n_8429, n9873);
  and g17940 (n9874, \a[17] , n_8429);
  and g17941 (n9875, n_8428, n_8429);
  not g17942 (n_8430, n9874);
  not g17943 (n_8431, n9875);
  and g17944 (n9876, n_8430, n_8431);
  not g17945 (n_8432, n9876);
  and g17946 (n9877, n9865, n_8432);
  not g17947 (n_8433, n9877);
  and g17948 (n9878, n9865, n_8433);
  and g17949 (n9879, n_8432, n_8433);
  not g17950 (n_8434, n9878);
  not g17951 (n_8435, n9879);
  and g17952 (n9880, n_8434, n_8435);
  and g17953 (n9881, n_8135, n_8141);
  and g17954 (n9882, n9880, n9881);
  not g17955 (n_8436, n9880);
  not g17956 (n_8437, n9881);
  and g17957 (n9883, n_8436, n_8437);
  not g17958 (n_8438, n9882);
  not g17959 (n_8439, n9883);
  and g17960 (n9884, n_8438, n_8439);
  and g17961 (n9885, \b[41] , n951);
  and g17962 (n9886, \b[39] , n1056);
  and g17963 (n9887, \b[40] , n946);
  and g17969 (n9890, n954, n6219);
  not g17972 (n_8444, n9891);
  and g17973 (n9892, \a[14] , n_8444);
  not g17974 (n_8445, n9892);
  and g17975 (n9893, \a[14] , n_8445);
  and g17976 (n9894, n_8444, n_8445);
  not g17977 (n_8446, n9893);
  not g17978 (n_8447, n9894);
  and g17979 (n9895, n_8446, n_8447);
  not g17980 (n_8448, n9895);
  and g17981 (n9896, n9884, n_8448);
  not g17982 (n_8449, n9896);
  and g17983 (n9897, n9884, n_8449);
  and g17984 (n9898, n_8448, n_8449);
  not g17985 (n_8450, n9897);
  not g17986 (n_8451, n9898);
  and g17987 (n9899, n_8450, n_8451);
  and g17988 (n9900, n_8151, n_8157);
  and g17989 (n9901, n9899, n9900);
  not g17990 (n_8452, n9899);
  not g17991 (n_8453, n9900);
  and g17992 (n9902, n_8452, n_8453);
  not g17993 (n_8454, n9901);
  not g17994 (n_8455, n9902);
  and g17995 (n9903, n_8454, n_8455);
  and g17996 (n9904, \b[44] , n700);
  and g17997 (n9905, \b[42] , n767);
  and g17998 (n9906, \b[43] , n695);
  and g18004 (n9909, n703, n7072);
  not g18007 (n_8460, n9910);
  and g18008 (n9911, \a[11] , n_8460);
  not g18009 (n_8461, n9911);
  and g18010 (n9912, \a[11] , n_8461);
  and g18011 (n9913, n_8460, n_8461);
  not g18012 (n_8462, n9912);
  not g18013 (n_8463, n9913);
  and g18014 (n9914, n_8462, n_8463);
  not g18015 (n_8464, n9914);
  and g18016 (n9915, n9903, n_8464);
  not g18017 (n_8465, n9903);
  and g18018 (n9916, n_8465, n9914);
  not g18019 (n_8466, n9576);
  not g18020 (n_8467, n9916);
  and g18021 (n9917, n_8466, n_8467);
  not g18022 (n_8468, n9915);
  and g18023 (n9918, n_8468, n9917);
  not g18024 (n_8469, n9918);
  and g18025 (n9919, n_8466, n_8469);
  and g18026 (n9920, n_8468, n_8469);
  and g18027 (n9921, n_8467, n9920);
  not g18028 (n_8470, n9919);
  not g18029 (n_8471, n9921);
  and g18030 (n9922, n_8470, n_8471);
  and g18031 (n9923, \b[47] , n511);
  and g18032 (n9924, \b[45] , n541);
  and g18033 (n9925, \b[46] , n506);
  and g18039 (n9928, n514, n7703);
  not g18042 (n_8476, n9929);
  and g18043 (n9930, \a[8] , n_8476);
  not g18044 (n_8477, n9930);
  and g18045 (n9931, \a[8] , n_8477);
  and g18046 (n9932, n_8476, n_8477);
  not g18047 (n_8478, n9931);
  not g18048 (n_8479, n9932);
  and g18049 (n9933, n_8478, n_8479);
  not g18050 (n_8480, n9922);
  not g18051 (n_8481, n9933);
  and g18052 (n9934, n_8480, n_8481);
  not g18053 (n_8482, n9934);
  and g18054 (n9935, n_8480, n_8482);
  and g18055 (n9936, n_8481, n_8482);
  not g18056 (n_8483, n9935);
  not g18057 (n_8484, n9936);
  and g18058 (n9937, n_8483, n_8484);
  and g18059 (n9938, n_8184, n_8191);
  and g18060 (n9939, n9937, n9938);
  not g18061 (n_8485, n9937);
  not g18062 (n_8486, n9938);
  and g18063 (n9940, n_8485, n_8486);
  not g18064 (n_8487, n9939);
  not g18065 (n_8488, n9940);
  and g18066 (n9941, n_8487, n_8488);
  and g18067 (n9942, \b[50] , n362);
  and g18068 (n9943, \b[48] , n403);
  and g18069 (n9944, \b[49] , n357);
  and g18075 (n9947, n365, n8949);
  not g18078 (n_8493, n9948);
  and g18079 (n9949, \a[5] , n_8493);
  not g18080 (n_8494, n9949);
  and g18081 (n9950, \a[5] , n_8494);
  and g18082 (n9951, n_8493, n_8494);
  not g18083 (n_8495, n9950);
  not g18084 (n_8496, n9951);
  and g18085 (n9952, n_8495, n_8496);
  not g18086 (n_8497, n9952);
  and g18087 (n9953, n9941, n_8497);
  not g18088 (n_8498, n9941);
  and g18089 (n9954, n_8498, n9952);
  not g18090 (n_8499, n9643);
  not g18091 (n_8500, n9954);
  and g18092 (n9955, n_8499, n_8500);
  not g18093 (n_8501, n9953);
  and g18094 (n9956, n_8501, n9955);
  not g18095 (n_8502, n9956);
  and g18096 (n9957, n_8499, n_8502);
  and g18097 (n9958, n_8501, n_8502);
  and g18098 (n9959, n_8500, n9958);
  not g18099 (n_8503, n9957);
  not g18100 (n_8504, n9959);
  and g18101 (n9960, n_8503, n_8504);
  and g18102 (n9961, \b[53] , n266);
  and g18103 (n9962, \b[51] , n284);
  and g18104 (n9963, \b[52] , n261);
  and g18110 (n9966, n_8214, n_8217);
  not g18111 (n_8509, \b[53] );
  and g18112 (n9967, n_8212, n_8509);
  and g18113 (n9968, \b[52] , \b[53] );
  not g18114 (n_8510, n9967);
  not g18115 (n_8511, n9968);
  and g18116 (n9969, n_8510, n_8511);
  not g18117 (n_8512, n9966);
  and g18118 (n9970, n_8512, n9969);
  not g18119 (n_8513, n9969);
  and g18120 (n9971, n9966, n_8513);
  not g18121 (n_8514, n9970);
  not g18122 (n_8515, n9971);
  and g18123 (n9972, n_8514, n_8515);
  and g18124 (n9973, n269, n9972);
  not g18127 (n_8517, n9974);
  and g18128 (n9975, \a[2] , n_8517);
  not g18129 (n_8518, n9975);
  and g18130 (n9976, \a[2] , n_8518);
  and g18131 (n9977, n_8517, n_8518);
  not g18132 (n_8519, n9976);
  not g18133 (n_8520, n9977);
  and g18134 (n9978, n_8519, n_8520);
  not g18135 (n_8521, n9960);
  and g18136 (n9979, n_8521, n9978);
  not g18137 (n_8522, n9978);
  and g18138 (n9980, n9960, n_8522);
  not g18139 (n_8523, n9979);
  not g18140 (n_8524, n9980);
  and g18141 (n9981, n_8523, n_8524);
  not g18142 (n_8525, n9641);
  not g18143 (n_8526, n9981);
  and g18144 (n9982, n_8525, n_8526);
  and g18145 (n9983, n9641, n9981);
  not g18146 (n_8527, n9982);
  not g18147 (n_8528, n9983);
  and g18148 (\f[53] , n_8527, n_8528);
  and g18149 (n9985, n_8521, n_8522);
  not g18150 (n_8529, n9985);
  and g18151 (n9986, n_8527, n_8529);
  and g18152 (n9987, \b[54] , n266);
  and g18153 (n9988, \b[52] , n284);
  and g18154 (n9989, \b[53] , n261);
  and g18160 (n9992, n_8511, n_8514);
  not g18161 (n_8534, \b[54] );
  and g18162 (n9993, n_8509, n_8534);
  and g18163 (n9994, \b[53] , \b[54] );
  not g18164 (n_8535, n9993);
  not g18165 (n_8536, n9994);
  and g18166 (n9995, n_8535, n_8536);
  not g18167 (n_8537, n9992);
  and g18168 (n9996, n_8537, n9995);
  not g18169 (n_8538, n9995);
  and g18170 (n9997, n9992, n_8538);
  not g18171 (n_8539, n9996);
  not g18172 (n_8540, n9997);
  and g18173 (n9998, n_8539, n_8540);
  and g18174 (n9999, n269, n9998);
  not g18177 (n_8542, n10000);
  and g18178 (n10001, \a[2] , n_8542);
  not g18179 (n_8543, n10001);
  and g18180 (n10002, \a[2] , n_8543);
  and g18181 (n10003, n_8542, n_8543);
  not g18182 (n_8544, n10002);
  not g18183 (n_8545, n10003);
  and g18184 (n10004, n_8544, n_8545);
  and g18185 (n10005, \b[45] , n700);
  and g18186 (n10006, \b[43] , n767);
  and g18187 (n10007, \b[44] , n695);
  and g18193 (n10010, n703, n7361);
  not g18196 (n_8550, n10011);
  and g18197 (n10012, \a[11] , n_8550);
  not g18198 (n_8551, n10012);
  and g18199 (n10013, \a[11] , n_8551);
  and g18200 (n10014, n_8550, n_8551);
  not g18201 (n_8552, n10013);
  not g18202 (n_8553, n10014);
  and g18203 (n10015, n_8552, n_8553);
  and g18204 (n10016, n_8449, n_8455);
  and g18205 (n10017, n_8417, n_8423);
  and g18206 (n10018, n_8411, n_8414);
  and g18207 (n10019, n_8403, n_8406);
  and g18208 (n10020, \b[30] , n2539);
  and g18209 (n10021, \b[28] , n2685);
  and g18210 (n10022, \b[29] , n2534);
  and g18216 (n10025, n2542, n3577);
  not g18219 (n_8558, n10026);
  and g18220 (n10027, \a[26] , n_8558);
  not g18221 (n_8559, n10027);
  and g18222 (n10028, \a[26] , n_8559);
  and g18223 (n10029, n_8558, n_8559);
  not g18224 (n_8560, n10028);
  not g18225 (n_8561, n10029);
  and g18226 (n10030, n_8560, n_8561);
  and g18227 (n10031, n_8395, n_8398);
  and g18228 (n10032, \b[27] , n3050);
  and g18229 (n10033, \b[25] , n3243);
  and g18230 (n10034, \b[26] , n3045);
  and g18236 (n10037, n2990, n3053);
  not g18239 (n_8566, n10038);
  and g18240 (n10039, \a[29] , n_8566);
  not g18241 (n_8567, n10039);
  and g18242 (n10040, \a[29] , n_8567);
  and g18243 (n10041, n_8566, n_8567);
  not g18244 (n_8568, n10040);
  not g18245 (n_8569, n10041);
  and g18246 (n10042, n_8568, n_8569);
  and g18247 (n10043, n_8376, n_8381);
  and g18248 (n10044, \b[24] , n3638);
  and g18249 (n10045, \b[22] , n3843);
  and g18250 (n10046, \b[23] , n3633);
  and g18256 (n10049, n2458, n3641);
  not g18259 (n_8574, n10050);
  and g18260 (n10051, \a[32] , n_8574);
  not g18261 (n_8575, n10051);
  and g18262 (n10052, \a[32] , n_8575);
  and g18263 (n10053, n_8574, n_8575);
  not g18264 (n_8576, n10052);
  not g18265 (n_8577, n10053);
  and g18266 (n10054, n_8576, n_8577);
  and g18267 (n10055, n_8368, n_8373);
  and g18268 (n10056, \b[21] , n4287);
  and g18269 (n10057, \b[19] , n4532);
  and g18270 (n10058, \b[20] , n4282);
  and g18276 (n10061, n1984, n4290);
  not g18279 (n_8582, n10062);
  and g18280 (n10063, \a[35] , n_8582);
  not g18281 (n_8583, n10063);
  and g18282 (n10064, \a[35] , n_8583);
  and g18283 (n10065, n_8582, n_8583);
  not g18284 (n_8584, n10064);
  not g18285 (n_8585, n10065);
  and g18286 (n10066, n_8584, n_8585);
  and g18287 (n10067, n_8350, n_8355);
  and g18288 (n10068, \b[18] , n5035);
  and g18289 (n10069, \b[16] , n5277);
  and g18290 (n10070, \b[17] , n5030);
  and g18296 (n10073, n1566, n5038);
  not g18299 (n_8590, n10074);
  and g18300 (n10075, \a[38] , n_8590);
  not g18301 (n_8591, n10075);
  and g18302 (n10076, \a[38] , n_8591);
  and g18303 (n10077, n_8590, n_8591);
  not g18304 (n_8592, n10076);
  not g18305 (n_8593, n10077);
  and g18306 (n10078, n_8592, n_8593);
  and g18307 (n10079, n_8342, n_8347);
  and g18308 (n10080, \b[15] , n5777);
  and g18309 (n10081, \b[13] , n6059);
  and g18310 (n10082, \b[14] , n5772);
  and g18316 (n10085, n1131, n5780);
  not g18319 (n_8598, n10086);
  and g18320 (n10087, \a[41] , n_8598);
  not g18321 (n_8599, n10087);
  and g18322 (n10088, \a[41] , n_8599);
  and g18323 (n10089, n_8598, n_8599);
  not g18324 (n_8600, n10088);
  not g18325 (n_8601, n10089);
  and g18326 (n10090, n_8600, n_8601);
  and g18327 (n10091, n_8336, n_8339);
  and g18328 (n10092, \b[12] , n6595);
  and g18329 (n10093, \b[10] , n6902);
  and g18330 (n10094, \b[11] , n6590);
  and g18336 (n10097, n842, n6598);
  not g18339 (n_8606, n10098);
  and g18340 (n10099, \a[44] , n_8606);
  not g18341 (n_8607, n10099);
  and g18342 (n10100, \a[44] , n_8607);
  and g18343 (n10101, n_8606, n_8607);
  not g18344 (n_8608, n10100);
  not g18345 (n_8609, n10101);
  and g18346 (n10102, n_8608, n_8609);
  and g18347 (n10103, n_8328, n_8331);
  and g18348 (n10104, \b[9] , n7446);
  and g18349 (n10105, \b[7] , n7787);
  and g18350 (n10106, \b[8] , n7441);
  and g18356 (n10109, n651, n7449);
  not g18359 (n_8614, n10110);
  and g18360 (n10111, \a[47] , n_8614);
  not g18361 (n_8615, n10111);
  and g18362 (n10112, \a[47] , n_8615);
  and g18363 (n10113, n_8614, n_8615);
  not g18364 (n_8616, n10112);
  not g18365 (n_8617, n10113);
  and g18366 (n10114, n_8616, n_8617);
  and g18367 (n10115, \b[6] , n8362);
  and g18368 (n10116, \b[4] , n8715);
  and g18369 (n10117, \b[5] , n8357);
  and g18375 (n10120, n459, n8365);
  not g18378 (n_8622, n10121);
  and g18379 (n10122, \a[50] , n_8622);
  not g18380 (n_8623, n10122);
  and g18381 (n10123, \a[50] , n_8623);
  and g18382 (n10124, n_8622, n_8623);
  not g18383 (n_8624, n10123);
  not g18384 (n_8625, n10124);
  and g18385 (n10125, n_8624, n_8625);
  not g18386 (n_8627, \a[54] );
  and g18387 (n10126, \a[53] , n_8627);
  and g18388 (n10127, n_7957, \a[54] );
  not g18389 (n_8628, n10126);
  not g18390 (n_8629, n10127);
  and g18391 (n10128, n_8628, n_8629);
  not g18392 (n_8630, n10128);
  and g18393 (n10129, \b[0] , n_8630);
  and g18394 (n10130, n_8300, n10129);
  not g18395 (n_8631, n10129);
  and g18396 (n10131, n9744, n_8631);
  not g18397 (n_8632, n10130);
  not g18398 (n_8633, n10131);
  and g18399 (n10132, n_8632, n_8633);
  and g18400 (n10133, \b[3] , n9339);
  and g18401 (n10134, \b[1] , n9732);
  and g18402 (n10135, \b[2] , n9334);
  and g18408 (n10138, n318, n9342);
  not g18411 (n_8638, n10139);
  and g18412 (n10140, \a[53] , n_8638);
  not g18413 (n_8639, n10140);
  and g18414 (n10141, \a[53] , n_8639);
  and g18415 (n10142, n_8638, n_8639);
  not g18416 (n_8640, n10141);
  not g18417 (n_8641, n10142);
  and g18418 (n10143, n_8640, n_8641);
  not g18419 (n_8642, n10132);
  not g18420 (n_8643, n10143);
  and g18421 (n10144, n_8642, n_8643);
  and g18422 (n10145, n10132, n10143);
  not g18423 (n_8644, n10144);
  not g18424 (n_8645, n10145);
  and g18425 (n10146, n_8644, n_8645);
  not g18426 (n_8646, n10125);
  and g18427 (n10147, n_8646, n10146);
  not g18428 (n_8647, n10147);
  and g18429 (n10148, n10146, n_8647);
  and g18430 (n10149, n_8646, n_8647);
  not g18431 (n_8648, n10148);
  not g18432 (n_8649, n10149);
  and g18433 (n10150, n_8648, n_8649);
  not g18434 (n_8650, n9762);
  not g18435 (n_8651, n10150);
  and g18436 (n10151, n_8650, n_8651);
  and g18437 (n10152, n9762, n10150);
  not g18438 (n_8652, n10151);
  not g18439 (n_8653, n10152);
  and g18440 (n10153, n_8652, n_8653);
  not g18441 (n_8654, n10114);
  and g18442 (n10154, n_8654, n10153);
  not g18443 (n_8655, n10154);
  and g18444 (n10155, n_8654, n_8655);
  and g18445 (n10156, n10153, n_8655);
  not g18446 (n_8656, n10155);
  not g18447 (n_8657, n10156);
  and g18448 (n10157, n_8656, n_8657);
  not g18449 (n_8658, n10103);
  not g18450 (n_8659, n10157);
  and g18451 (n10158, n_8658, n_8659);
  and g18452 (n10159, n10103, n_8657);
  and g18453 (n10160, n_8656, n10159);
  not g18454 (n_8660, n10158);
  not g18455 (n_8661, n10160);
  and g18456 (n10161, n_8660, n_8661);
  not g18457 (n_8662, n10102);
  and g18458 (n10162, n_8662, n10161);
  not g18459 (n_8663, n10162);
  and g18460 (n10163, n_8662, n_8663);
  and g18461 (n10164, n10161, n_8663);
  not g18462 (n_8664, n10163);
  not g18463 (n_8665, n10164);
  and g18464 (n10165, n_8664, n_8665);
  not g18465 (n_8666, n10091);
  not g18466 (n_8667, n10165);
  and g18467 (n10166, n_8666, n_8667);
  and g18468 (n10167, n10091, n_8665);
  and g18469 (n10168, n_8664, n10167);
  not g18470 (n_8668, n10166);
  not g18471 (n_8669, n10168);
  and g18472 (n10169, n_8668, n_8669);
  not g18473 (n_8670, n10090);
  and g18474 (n10170, n_8670, n10169);
  not g18475 (n_8671, n10169);
  and g18476 (n10171, n10090, n_8671);
  not g18477 (n_8672, n10170);
  not g18478 (n_8673, n10171);
  and g18479 (n10172, n_8672, n_8673);
  not g18480 (n_8674, n10079);
  and g18481 (n10173, n_8674, n10172);
  not g18482 (n_8675, n10172);
  and g18483 (n10174, n10079, n_8675);
  not g18484 (n_8676, n10173);
  not g18485 (n_8677, n10174);
  and g18486 (n10175, n_8676, n_8677);
  not g18487 (n_8678, n10078);
  and g18488 (n10176, n_8678, n10175);
  not g18489 (n_8679, n10176);
  and g18490 (n10177, n_8678, n_8679);
  and g18491 (n10178, n10175, n_8679);
  not g18492 (n_8680, n10177);
  not g18493 (n_8681, n10178);
  and g18494 (n10179, n_8680, n_8681);
  not g18495 (n_8682, n10067);
  not g18496 (n_8683, n10179);
  and g18497 (n10180, n_8682, n_8683);
  and g18498 (n10181, n10067, n_8681);
  and g18499 (n10182, n_8680, n10181);
  not g18500 (n_8684, n10180);
  not g18501 (n_8685, n10182);
  and g18502 (n10183, n_8684, n_8685);
  not g18503 (n_8686, n10066);
  and g18504 (n10184, n_8686, n10183);
  not g18505 (n_8687, n10183);
  and g18506 (n10185, n10066, n_8687);
  not g18507 (n_8688, n10184);
  not g18508 (n_8689, n10185);
  and g18509 (n10186, n_8688, n_8689);
  not g18510 (n_8690, n10055);
  and g18511 (n10187, n_8690, n10186);
  not g18512 (n_8691, n10186);
  and g18513 (n10188, n10055, n_8691);
  not g18514 (n_8692, n10187);
  not g18515 (n_8693, n10188);
  and g18516 (n10189, n_8692, n_8693);
  not g18517 (n_8694, n10054);
  and g18518 (n10190, n_8694, n10189);
  not g18519 (n_8695, n10189);
  and g18520 (n10191, n10054, n_8695);
  not g18521 (n_8696, n10190);
  not g18522 (n_8697, n10191);
  and g18523 (n10192, n_8696, n_8697);
  not g18524 (n_8698, n10043);
  and g18525 (n10193, n_8698, n10192);
  not g18526 (n_8699, n10192);
  and g18527 (n10194, n10043, n_8699);
  not g18528 (n_8700, n10193);
  not g18529 (n_8701, n10194);
  and g18530 (n10195, n_8700, n_8701);
  not g18531 (n_8702, n10042);
  and g18532 (n10196, n_8702, n10195);
  not g18533 (n_8703, n10195);
  and g18534 (n10197, n10042, n_8703);
  not g18535 (n_8704, n10196);
  not g18536 (n_8705, n10197);
  and g18537 (n10198, n_8704, n_8705);
  not g18538 (n_8706, n10031);
  and g18539 (n10199, n_8706, n10198);
  not g18540 (n_8707, n10198);
  and g18541 (n10200, n10031, n_8707);
  not g18542 (n_8708, n10199);
  not g18543 (n_8709, n10200);
  and g18544 (n10201, n_8708, n_8709);
  not g18545 (n_8710, n10030);
  and g18546 (n10202, n_8710, n10201);
  not g18547 (n_8711, n10201);
  and g18548 (n10203, n10030, n_8711);
  not g18549 (n_8712, n10202);
  not g18550 (n_8713, n10203);
  and g18551 (n10204, n_8712, n_8713);
  not g18552 (n_8714, n10019);
  and g18553 (n10205, n_8714, n10204);
  not g18554 (n_8715, n10204);
  and g18555 (n10206, n10019, n_8715);
  not g18556 (n_8716, n10205);
  not g18557 (n_8717, n10206);
  and g18558 (n10207, n_8716, n_8717);
  and g18559 (n10208, \b[33] , n2048);
  and g18560 (n10209, \b[31] , n2198);
  and g18561 (n10210, \b[32] , n2043);
  and g18567 (n10213, n2051, n4223);
  not g18570 (n_8722, n10214);
  and g18571 (n10215, \a[23] , n_8722);
  not g18572 (n_8723, n10215);
  and g18573 (n10216, \a[23] , n_8723);
  and g18574 (n10217, n_8722, n_8723);
  not g18575 (n_8724, n10216);
  not g18576 (n_8725, n10217);
  and g18577 (n10218, n_8724, n_8725);
  not g18578 (n_8726, n10218);
  and g18579 (n10219, n10207, n_8726);
  not g18580 (n_8727, n10219);
  and g18581 (n10220, n10207, n_8727);
  and g18582 (n10221, n_8726, n_8727);
  not g18583 (n_8728, n10220);
  not g18584 (n_8729, n10221);
  and g18585 (n10222, n_8728, n_8729);
  not g18586 (n_8730, n10018);
  and g18587 (n10223, n_8730, n10222);
  not g18588 (n_8731, n10222);
  and g18589 (n10224, n10018, n_8731);
  not g18590 (n_8732, n10223);
  not g18591 (n_8733, n10224);
  and g18592 (n10225, n_8732, n_8733);
  and g18593 (n10226, \b[36] , n1627);
  and g18594 (n10227, \b[34] , n1763);
  and g18595 (n10228, \b[35] , n1622);
  and g18601 (n10231, n1630, n4922);
  not g18604 (n_8738, n10232);
  and g18605 (n10233, \a[20] , n_8738);
  not g18606 (n_8739, n10233);
  and g18607 (n10234, \a[20] , n_8739);
  and g18608 (n10235, n_8738, n_8739);
  not g18609 (n_8740, n10234);
  not g18610 (n_8741, n10235);
  and g18611 (n10236, n_8740, n_8741);
  not g18612 (n_8742, n10225);
  not g18613 (n_8743, n10236);
  and g18614 (n10237, n_8742, n_8743);
  and g18615 (n10238, n10225, n10236);
  not g18616 (n_8744, n10237);
  not g18617 (n_8745, n10238);
  and g18618 (n10239, n_8744, n_8745);
  not g18619 (n_8746, n10239);
  and g18620 (n10240, n10017, n_8746);
  not g18621 (n_8747, n10017);
  and g18622 (n10241, n_8747, n10239);
  not g18623 (n_8748, n10240);
  not g18624 (n_8749, n10241);
  and g18625 (n10242, n_8748, n_8749);
  and g18626 (n10243, \b[39] , n1302);
  and g18627 (n10244, \b[37] , n1391);
  and g18628 (n10245, \b[38] , n1297);
  and g18634 (n10248, n1305, n5451);
  not g18637 (n_8754, n10249);
  and g18638 (n10250, \a[17] , n_8754);
  not g18639 (n_8755, n10250);
  and g18640 (n10251, \a[17] , n_8755);
  and g18641 (n10252, n_8754, n_8755);
  not g18642 (n_8756, n10251);
  not g18643 (n_8757, n10252);
  and g18644 (n10253, n_8756, n_8757);
  not g18645 (n_8758, n10253);
  and g18646 (n10254, n10242, n_8758);
  not g18647 (n_8759, n10254);
  and g18648 (n10255, n10242, n_8759);
  and g18649 (n10256, n_8758, n_8759);
  not g18650 (n_8760, n10255);
  not g18651 (n_8761, n10256);
  and g18652 (n10257, n_8760, n_8761);
  and g18653 (n10258, n_8433, n_8439);
  and g18654 (n10259, n10257, n10258);
  not g18655 (n_8762, n10257);
  not g18656 (n_8763, n10258);
  and g18657 (n10260, n_8762, n_8763);
  not g18658 (n_8764, n10259);
  not g18659 (n_8765, n10260);
  and g18660 (n10261, n_8764, n_8765);
  and g18661 (n10262, \b[42] , n951);
  and g18662 (n10263, \b[40] , n1056);
  and g18663 (n10264, \b[41] , n946);
  and g18669 (n10267, n954, n6489);
  not g18672 (n_8770, n10268);
  and g18673 (n10269, \a[14] , n_8770);
  not g18674 (n_8771, n10269);
  and g18675 (n10270, \a[14] , n_8771);
  and g18676 (n10271, n_8770, n_8771);
  not g18677 (n_8772, n10270);
  not g18678 (n_8773, n10271);
  and g18679 (n10272, n_8772, n_8773);
  not g18680 (n_8774, n10261);
  and g18681 (n10273, n_8774, n10272);
  not g18682 (n_8775, n10272);
  and g18683 (n10274, n10261, n_8775);
  not g18684 (n_8776, n10273);
  not g18685 (n_8777, n10274);
  and g18686 (n10275, n_8776, n_8777);
  not g18687 (n_8778, n10016);
  and g18688 (n10276, n_8778, n10275);
  not g18689 (n_8779, n10275);
  and g18690 (n10277, n10016, n_8779);
  not g18691 (n_8780, n10276);
  not g18692 (n_8781, n10277);
  and g18693 (n10278, n_8780, n_8781);
  not g18694 (n_8782, n10015);
  and g18695 (n10279, n_8782, n10278);
  not g18696 (n_8783, n10279);
  and g18697 (n10280, n_8782, n_8783);
  and g18698 (n10281, n10278, n_8783);
  not g18699 (n_8784, n10280);
  not g18700 (n_8785, n10281);
  and g18701 (n10282, n_8784, n_8785);
  not g18702 (n_8786, n9920);
  not g18703 (n_8787, n10282);
  and g18704 (n10283, n_8786, n_8787);
  not g18705 (n_8788, n10283);
  and g18706 (n10284, n_8786, n_8788);
  and g18707 (n10285, n_8787, n_8788);
  not g18708 (n_8789, n10284);
  not g18709 (n_8790, n10285);
  and g18710 (n10286, n_8789, n_8790);
  and g18711 (n10287, \b[48] , n511);
  and g18712 (n10288, \b[46] , n541);
  and g18713 (n10289, \b[47] , n506);
  and g18719 (n10292, n514, n8009);
  not g18722 (n_8795, n10293);
  and g18723 (n10294, \a[8] , n_8795);
  not g18724 (n_8796, n10294);
  and g18725 (n10295, \a[8] , n_8796);
  and g18726 (n10296, n_8795, n_8796);
  not g18727 (n_8797, n10295);
  not g18728 (n_8798, n10296);
  and g18729 (n10297, n_8797, n_8798);
  not g18730 (n_8799, n10286);
  not g18731 (n_8800, n10297);
  and g18732 (n10298, n_8799, n_8800);
  not g18733 (n_8801, n10298);
  and g18734 (n10299, n_8799, n_8801);
  and g18735 (n10300, n_8800, n_8801);
  not g18736 (n_8802, n10299);
  not g18737 (n_8803, n10300);
  and g18738 (n10301, n_8802, n_8803);
  and g18739 (n10302, n_8482, n_8488);
  and g18740 (n10303, n10301, n10302);
  not g18741 (n_8804, n10301);
  not g18742 (n_8805, n10302);
  and g18743 (n10304, n_8804, n_8805);
  not g18744 (n_8806, n10303);
  not g18745 (n_8807, n10304);
  and g18746 (n10305, n_8806, n_8807);
  and g18747 (n10306, \b[51] , n362);
  and g18748 (n10307, \b[49] , n403);
  and g18749 (n10308, \b[50] , n357);
  and g18755 (n10311, n365, n8976);
  not g18758 (n_8812, n10312);
  and g18759 (n10313, \a[5] , n_8812);
  not g18760 (n_8813, n10313);
  and g18761 (n10314, \a[5] , n_8813);
  and g18762 (n10315, n_8812, n_8813);
  not g18763 (n_8814, n10314);
  not g18764 (n_8815, n10315);
  and g18765 (n10316, n_8814, n_8815);
  not g18766 (n_8816, n10305);
  and g18767 (n10317, n_8816, n10316);
  not g18768 (n_8817, n10316);
  and g18769 (n10318, n10305, n_8817);
  not g18770 (n_8818, n10317);
  not g18771 (n_8819, n10318);
  and g18772 (n10319, n_8818, n_8819);
  not g18773 (n_8820, n9958);
  and g18774 (n10320, n_8820, n10319);
  not g18775 (n_8821, n10319);
  and g18776 (n10321, n9958, n_8821);
  not g18777 (n_8822, n10320);
  not g18778 (n_8823, n10321);
  and g18779 (n10322, n_8822, n_8823);
  not g18780 (n_8824, n10004);
  and g18781 (n10323, n_8824, n10322);
  not g18782 (n_8825, n10322);
  and g18783 (n10324, n10004, n_8825);
  not g18784 (n_8826, n10323);
  not g18785 (n_8827, n10324);
  and g18786 (n10325, n_8826, n_8827);
  not g18787 (n_8828, n9986);
  and g18788 (n10326, n_8828, n10325);
  not g18789 (n_8829, n10325);
  and g18790 (n10327, n9986, n_8829);
  not g18791 (n_8830, n10326);
  not g18792 (n_8831, n10327);
  and g18793 (\f[54] , n_8830, n_8831);
  and g18794 (n10329, n_8826, n_8830);
  and g18795 (n10330, n_8819, n_8822);
  and g18796 (n10331, \b[52] , n362);
  and g18797 (n10332, \b[50] , n403);
  and g18798 (n10333, \b[51] , n357);
  and g18804 (n10336, n365, n9628);
  not g18807 (n_8836, n10337);
  and g18808 (n10338, \a[5] , n_8836);
  not g18809 (n_8837, n10338);
  and g18810 (n10339, \a[5] , n_8837);
  and g18811 (n10340, n_8836, n_8837);
  not g18812 (n_8838, n10339);
  not g18813 (n_8839, n10340);
  and g18814 (n10341, n_8838, n_8839);
  and g18815 (n10342, n_8801, n_8807);
  and g18816 (n10343, \b[49] , n511);
  and g18817 (n10344, \b[47] , n541);
  and g18818 (n10345, \b[48] , n506);
  and g18824 (n10348, n514, n8625);
  not g18827 (n_8844, n10349);
  and g18828 (n10350, \a[8] , n_8844);
  not g18829 (n_8845, n10350);
  and g18830 (n10351, \a[8] , n_8845);
  and g18831 (n10352, n_8844, n_8845);
  not g18832 (n_8846, n10351);
  not g18833 (n_8847, n10352);
  and g18834 (n10353, n_8846, n_8847);
  and g18835 (n10354, n_8783, n_8788);
  and g18836 (n10355, n_8777, n_8780);
  and g18837 (n10356, n_8679, n_8684);
  and g18838 (n10357, \b[16] , n5777);
  and g18839 (n10358, \b[14] , n6059);
  and g18840 (n10359, \b[15] , n5772);
  and g18846 (n10362, n1237, n5780);
  not g18849 (n_8852, n10363);
  and g18850 (n10364, \a[41] , n_8852);
  not g18851 (n_8853, n10364);
  and g18852 (n10365, \a[41] , n_8853);
  and g18853 (n10366, n_8852, n_8853);
  not g18854 (n_8854, n10365);
  not g18855 (n_8855, n10366);
  and g18856 (n10367, n_8854, n_8855);
  and g18857 (n10368, n_8663, n_8668);
  and g18858 (n10369, \b[13] , n6595);
  and g18859 (n10370, \b[11] , n6902);
  and g18860 (n10371, \b[12] , n6590);
  and g18866 (n10374, n1008, n6598);
  not g18869 (n_8860, n10375);
  and g18870 (n10376, \a[44] , n_8860);
  not g18871 (n_8861, n10376);
  and g18872 (n10377, \a[44] , n_8861);
  and g18873 (n10378, n_8860, n_8861);
  not g18874 (n_8862, n10377);
  not g18875 (n_8863, n10378);
  and g18876 (n10379, n_8862, n_8863);
  and g18877 (n10380, n_8655, n_8660);
  and g18878 (n10381, \b[10] , n7446);
  and g18879 (n10382, \b[8] , n7787);
  and g18880 (n10383, \b[9] , n7441);
  and g18886 (n10386, n738, n7449);
  not g18889 (n_8868, n10387);
  and g18890 (n10388, \a[47] , n_8868);
  not g18891 (n_8869, n10388);
  and g18892 (n10389, \a[47] , n_8869);
  and g18893 (n10390, n_8868, n_8869);
  not g18894 (n_8870, n10389);
  not g18895 (n_8871, n10390);
  and g18896 (n10391, n_8870, n_8871);
  and g18897 (n10392, n_8647, n_8652);
  and g18898 (n10393, \b[7] , n8362);
  and g18899 (n10394, \b[5] , n8715);
  and g18900 (n10395, \b[6] , n8357);
  and g18906 (n10398, n484, n8365);
  not g18909 (n_8876, n10399);
  and g18910 (n10400, \a[50] , n_8876);
  not g18911 (n_8877, n10400);
  and g18912 (n10401, \a[50] , n_8877);
  and g18913 (n10402, n_8876, n_8877);
  not g18914 (n_8878, n10401);
  not g18915 (n_8879, n10402);
  and g18916 (n10403, n_8878, n_8879);
  and g18917 (n10404, n9744, n10129);
  not g18918 (n_8880, n10404);
  and g18919 (n10405, n_8644, n_8880);
  and g18920 (n10406, \b[4] , n9339);
  and g18921 (n10407, \b[2] , n9732);
  and g18922 (n10408, \b[3] , n9334);
  and g18928 (n10411, n346, n9342);
  not g18931 (n_8885, n10412);
  and g18932 (n10413, \a[53] , n_8885);
  not g18933 (n_8886, n10413);
  and g18934 (n10414, \a[53] , n_8886);
  and g18935 (n10415, n_8885, n_8886);
  not g18936 (n_8887, n10414);
  not g18937 (n_8888, n10415);
  and g18938 (n10416, n_8887, n_8888);
  and g18939 (n10417, \a[56] , n_8631);
  and g18940 (n10418, n_8627, \a[55] );
  not g18941 (n_8891, \a[55] );
  and g18942 (n10419, \a[54] , n_8891);
  not g18943 (n_8892, n10418);
  not g18944 (n_8893, n10419);
  and g18945 (n10420, n_8892, n_8893);
  not g18946 (n_8894, n10420);
  and g18947 (n10421, n10128, n_8894);
  and g18948 (n10422, \b[0] , n10421);
  and g18949 (n10423, n_8891, \a[56] );
  not g18950 (n_8895, \a[56] );
  and g18951 (n10424, \a[55] , n_8895);
  not g18952 (n_8896, n10423);
  not g18953 (n_8897, n10424);
  and g18954 (n10425, n_8896, n_8897);
  and g18955 (n10426, n_8630, n10425);
  and g18956 (n10427, \b[1] , n10426);
  not g18957 (n_8898, n10422);
  not g18958 (n_8899, n10427);
  and g18959 (n10428, n_8898, n_8899);
  not g18960 (n_8900, n10425);
  and g18961 (n10429, n_8630, n_8900);
  and g18962 (n10430, n_21, n10429);
  not g18963 (n_8901, n10430);
  and g18964 (n10431, n10428, n_8901);
  not g18965 (n_8902, n10431);
  and g18966 (n10432, \a[56] , n_8902);
  not g18967 (n_8903, n10432);
  and g18968 (n10433, \a[56] , n_8903);
  and g18969 (n10434, n_8902, n_8903);
  not g18970 (n_8904, n10433);
  not g18971 (n_8905, n10434);
  and g18972 (n10435, n_8904, n_8905);
  not g18973 (n_8906, n10435);
  and g18974 (n10436, n10417, n_8906);
  not g18975 (n_8907, n10417);
  and g18976 (n10437, n_8907, n10435);
  not g18977 (n_8908, n10436);
  not g18978 (n_8909, n10437);
  and g18979 (n10438, n_8908, n_8909);
  not g18980 (n_8910, n10438);
  and g18981 (n10439, n10416, n_8910);
  not g18982 (n_8911, n10416);
  and g18983 (n10440, n_8911, n10438);
  not g18984 (n_8912, n10439);
  not g18985 (n_8913, n10440);
  and g18986 (n10441, n_8912, n_8913);
  not g18987 (n_8914, n10405);
  and g18988 (n10442, n_8914, n10441);
  not g18989 (n_8915, n10441);
  and g18990 (n10443, n10405, n_8915);
  not g18991 (n_8916, n10442);
  not g18992 (n_8917, n10443);
  and g18993 (n10444, n_8916, n_8917);
  not g18994 (n_8918, n10444);
  and g18995 (n10445, n10403, n_8918);
  not g18996 (n_8919, n10403);
  and g18997 (n10446, n_8919, n10444);
  not g18998 (n_8920, n10445);
  not g18999 (n_8921, n10446);
  and g19000 (n10447, n_8920, n_8921);
  not g19001 (n_8922, n10392);
  and g19002 (n10448, n_8922, n10447);
  not g19003 (n_8923, n10447);
  and g19004 (n10449, n10392, n_8923);
  not g19005 (n_8924, n10448);
  not g19006 (n_8925, n10449);
  and g19007 (n10450, n_8924, n_8925);
  not g19008 (n_8926, n10450);
  and g19009 (n10451, n10391, n_8926);
  not g19010 (n_8927, n10391);
  and g19011 (n10452, n_8927, n10450);
  not g19012 (n_8928, n10451);
  not g19013 (n_8929, n10452);
  and g19014 (n10453, n_8928, n_8929);
  not g19015 (n_8930, n10380);
  and g19016 (n10454, n_8930, n10453);
  not g19017 (n_8931, n10453);
  and g19018 (n10455, n10380, n_8931);
  not g19019 (n_8932, n10454);
  not g19020 (n_8933, n10455);
  and g19021 (n10456, n_8932, n_8933);
  not g19022 (n_8934, n10456);
  and g19023 (n10457, n10379, n_8934);
  not g19024 (n_8935, n10379);
  and g19025 (n10458, n_8935, n10456);
  not g19026 (n_8936, n10457);
  not g19027 (n_8937, n10458);
  and g19028 (n10459, n_8936, n_8937);
  not g19029 (n_8938, n10368);
  and g19030 (n10460, n_8938, n10459);
  not g19031 (n_8939, n10459);
  and g19032 (n10461, n10368, n_8939);
  not g19033 (n_8940, n10460);
  not g19034 (n_8941, n10461);
  and g19035 (n10462, n_8940, n_8941);
  not g19036 (n_8942, n10367);
  and g19037 (n10463, n_8942, n10462);
  not g19038 (n_8943, n10463);
  and g19039 (n10464, n10462, n_8943);
  and g19040 (n10465, n_8942, n_8943);
  not g19041 (n_8944, n10464);
  not g19042 (n_8945, n10465);
  and g19043 (n10466, n_8944, n_8945);
  and g19044 (n10467, n_8672, n_8676);
  and g19045 (n10468, n10466, n10467);
  not g19046 (n_8946, n10466);
  not g19047 (n_8947, n10467);
  and g19048 (n10469, n_8946, n_8947);
  not g19049 (n_8948, n10468);
  not g19050 (n_8949, n10469);
  and g19051 (n10470, n_8948, n_8949);
  and g19052 (n10471, \b[19] , n5035);
  and g19053 (n10472, \b[17] , n5277);
  and g19054 (n10473, \b[18] , n5030);
  and g19060 (n10476, n1708, n5038);
  not g19063 (n_8954, n10477);
  and g19064 (n10478, \a[38] , n_8954);
  not g19065 (n_8955, n10478);
  and g19066 (n10479, \a[38] , n_8955);
  and g19067 (n10480, n_8954, n_8955);
  not g19068 (n_8956, n10479);
  not g19069 (n_8957, n10480);
  and g19070 (n10481, n_8956, n_8957);
  not g19071 (n_8958, n10481);
  and g19072 (n10482, n10470, n_8958);
  not g19073 (n_8959, n10470);
  and g19074 (n10483, n_8959, n10481);
  not g19075 (n_8960, n10356);
  not g19076 (n_8961, n10483);
  and g19077 (n10484, n_8960, n_8961);
  not g19078 (n_8962, n10482);
  and g19079 (n10485, n_8962, n10484);
  not g19080 (n_8963, n10485);
  and g19081 (n10486, n_8960, n_8963);
  and g19082 (n10487, n_8962, n_8963);
  and g19083 (n10488, n_8961, n10487);
  not g19084 (n_8964, n10486);
  not g19085 (n_8965, n10488);
  and g19086 (n10489, n_8964, n_8965);
  and g19087 (n10490, \b[22] , n4287);
  and g19088 (n10491, \b[20] , n4532);
  and g19089 (n10492, \b[21] , n4282);
  and g19095 (n10495, n2145, n4290);
  not g19098 (n_8970, n10496);
  and g19099 (n10497, \a[35] , n_8970);
  not g19100 (n_8971, n10497);
  and g19101 (n10498, \a[35] , n_8971);
  and g19102 (n10499, n_8970, n_8971);
  not g19103 (n_8972, n10498);
  not g19104 (n_8973, n10499);
  and g19105 (n10500, n_8972, n_8973);
  not g19106 (n_8974, n10489);
  not g19107 (n_8975, n10500);
  and g19108 (n10501, n_8974, n_8975);
  not g19109 (n_8976, n10501);
  and g19110 (n10502, n_8974, n_8976);
  and g19111 (n10503, n_8975, n_8976);
  not g19112 (n_8977, n10502);
  not g19113 (n_8978, n10503);
  and g19114 (n10504, n_8977, n_8978);
  and g19115 (n10505, n_8688, n_8692);
  and g19116 (n10506, n10504, n10505);
  not g19117 (n_8979, n10504);
  not g19118 (n_8980, n10505);
  and g19119 (n10507, n_8979, n_8980);
  not g19120 (n_8981, n10506);
  not g19121 (n_8982, n10507);
  and g19122 (n10508, n_8981, n_8982);
  and g19123 (n10509, \b[25] , n3638);
  and g19124 (n10510, \b[23] , n3843);
  and g19125 (n10511, \b[24] , n3633);
  and g19131 (n10514, n2485, n3641);
  not g19134 (n_8987, n10515);
  and g19135 (n10516, \a[32] , n_8987);
  not g19136 (n_8988, n10516);
  and g19137 (n10517, \a[32] , n_8988);
  and g19138 (n10518, n_8987, n_8988);
  not g19139 (n_8989, n10517);
  not g19140 (n_8990, n10518);
  and g19141 (n10519, n_8989, n_8990);
  not g19142 (n_8991, n10519);
  and g19143 (n10520, n10508, n_8991);
  not g19144 (n_8992, n10520);
  and g19145 (n10521, n10508, n_8992);
  and g19146 (n10522, n_8991, n_8992);
  not g19147 (n_8993, n10521);
  not g19148 (n_8994, n10522);
  and g19149 (n10523, n_8993, n_8994);
  and g19150 (n10524, n_8696, n_8700);
  and g19151 (n10525, n10523, n10524);
  not g19152 (n_8995, n10523);
  not g19153 (n_8996, n10524);
  and g19154 (n10526, n_8995, n_8996);
  not g19155 (n_8997, n10525);
  not g19156 (n_8998, n10526);
  and g19157 (n10527, n_8997, n_8998);
  and g19158 (n10528, \b[28] , n3050);
  and g19159 (n10529, \b[26] , n3243);
  and g19160 (n10530, \b[27] , n3045);
  and g19166 (n10533, n3053, n3189);
  not g19169 (n_9003, n10534);
  and g19170 (n10535, \a[29] , n_9003);
  not g19171 (n_9004, n10535);
  and g19172 (n10536, \a[29] , n_9004);
  and g19173 (n10537, n_9003, n_9004);
  not g19174 (n_9005, n10536);
  not g19175 (n_9006, n10537);
  and g19176 (n10538, n_9005, n_9006);
  not g19177 (n_9007, n10538);
  and g19178 (n10539, n10527, n_9007);
  not g19179 (n_9008, n10539);
  and g19180 (n10540, n10527, n_9008);
  and g19181 (n10541, n_9007, n_9008);
  not g19182 (n_9009, n10540);
  not g19183 (n_9010, n10541);
  and g19184 (n10542, n_9009, n_9010);
  and g19185 (n10543, n_8704, n_8708);
  and g19186 (n10544, n10542, n10543);
  not g19187 (n_9011, n10542);
  not g19188 (n_9012, n10543);
  and g19189 (n10545, n_9011, n_9012);
  not g19190 (n_9013, n10544);
  not g19191 (n_9014, n10545);
  and g19192 (n10546, n_9013, n_9014);
  and g19193 (n10547, \b[31] , n2539);
  and g19194 (n10548, \b[29] , n2685);
  and g19195 (n10549, \b[30] , n2534);
  and g19201 (n10552, n2542, n3796);
  not g19204 (n_9019, n10553);
  and g19205 (n10554, \a[26] , n_9019);
  not g19206 (n_9020, n10554);
  and g19207 (n10555, \a[26] , n_9020);
  and g19208 (n10556, n_9019, n_9020);
  not g19209 (n_9021, n10555);
  not g19210 (n_9022, n10556);
  and g19211 (n10557, n_9021, n_9022);
  not g19212 (n_9023, n10557);
  and g19213 (n10558, n10546, n_9023);
  not g19214 (n_9024, n10558);
  and g19215 (n10559, n10546, n_9024);
  and g19216 (n10560, n_9023, n_9024);
  not g19217 (n_9025, n10559);
  not g19218 (n_9026, n10560);
  and g19219 (n10561, n_9025, n_9026);
  and g19220 (n10562, n_8712, n_8716);
  and g19221 (n10563, n10561, n10562);
  not g19222 (n_9027, n10561);
  not g19223 (n_9028, n10562);
  and g19224 (n10564, n_9027, n_9028);
  not g19225 (n_9029, n10563);
  not g19226 (n_9030, n10564);
  and g19227 (n10565, n_9029, n_9030);
  and g19228 (n10566, \b[34] , n2048);
  and g19229 (n10567, \b[32] , n2198);
  and g19230 (n10568, \b[33] , n2043);
  and g19236 (n10571, n2051, n4466);
  not g19239 (n_9035, n10572);
  and g19240 (n10573, \a[23] , n_9035);
  not g19241 (n_9036, n10573);
  and g19242 (n10574, \a[23] , n_9036);
  and g19243 (n10575, n_9035, n_9036);
  not g19244 (n_9037, n10574);
  not g19245 (n_9038, n10575);
  and g19246 (n10576, n_9037, n_9038);
  not g19247 (n_9039, n10576);
  and g19248 (n10577, n10565, n_9039);
  not g19249 (n_9040, n10577);
  and g19250 (n10578, n10565, n_9040);
  and g19251 (n10579, n_9039, n_9040);
  not g19252 (n_9041, n10578);
  not g19253 (n_9042, n10579);
  and g19254 (n10580, n_9041, n_9042);
  and g19255 (n10581, n_8730, n_8731);
  not g19256 (n_9043, n10581);
  and g19257 (n10582, n_8727, n_9043);
  and g19258 (n10583, n10580, n10582);
  not g19259 (n_9044, n10580);
  not g19260 (n_9045, n10582);
  and g19261 (n10584, n_9044, n_9045);
  not g19262 (n_9046, n10583);
  not g19263 (n_9047, n10584);
  and g19264 (n10585, n_9046, n_9047);
  and g19265 (n10586, \b[37] , n1627);
  and g19266 (n10587, \b[35] , n1763);
  and g19267 (n10588, \b[36] , n1622);
  and g19273 (n10591, n1630, n5181);
  not g19276 (n_9052, n10592);
  and g19277 (n10593, \a[20] , n_9052);
  not g19278 (n_9053, n10593);
  and g19279 (n10594, \a[20] , n_9053);
  and g19280 (n10595, n_9052, n_9053);
  not g19281 (n_9054, n10594);
  not g19282 (n_9055, n10595);
  and g19283 (n10596, n_9054, n_9055);
  not g19284 (n_9056, n10596);
  and g19285 (n10597, n10585, n_9056);
  not g19286 (n_9057, n10597);
  and g19287 (n10598, n10585, n_9057);
  and g19288 (n10599, n_9056, n_9057);
  not g19289 (n_9058, n10598);
  not g19290 (n_9059, n10599);
  and g19291 (n10600, n_9058, n_9059);
  and g19292 (n10601, n_8744, n_8749);
  and g19293 (n10602, n10600, n10601);
  not g19294 (n_9060, n10600);
  not g19295 (n_9061, n10601);
  and g19296 (n10603, n_9060, n_9061);
  not g19297 (n_9062, n10602);
  not g19298 (n_9063, n10603);
  and g19299 (n10604, n_9062, n_9063);
  and g19300 (n10605, \b[40] , n1302);
  and g19301 (n10606, \b[38] , n1391);
  and g19302 (n10607, \b[39] , n1297);
  and g19308 (n10610, n1305, n5955);
  not g19311 (n_9068, n10611);
  and g19312 (n10612, \a[17] , n_9068);
  not g19313 (n_9069, n10612);
  and g19314 (n10613, \a[17] , n_9069);
  and g19315 (n10614, n_9068, n_9069);
  not g19316 (n_9070, n10613);
  not g19317 (n_9071, n10614);
  and g19318 (n10615, n_9070, n_9071);
  not g19319 (n_9072, n10615);
  and g19320 (n10616, n10604, n_9072);
  not g19321 (n_9073, n10616);
  and g19322 (n10617, n10604, n_9073);
  and g19323 (n10618, n_9072, n_9073);
  not g19324 (n_9074, n10617);
  not g19325 (n_9075, n10618);
  and g19326 (n10619, n_9074, n_9075);
  and g19327 (n10620, n_8759, n_8765);
  and g19328 (n10621, n10619, n10620);
  not g19329 (n_9076, n10619);
  not g19330 (n_9077, n10620);
  and g19331 (n10622, n_9076, n_9077);
  not g19332 (n_9078, n10621);
  not g19333 (n_9079, n10622);
  and g19334 (n10623, n_9078, n_9079);
  and g19335 (n10624, \b[43] , n951);
  and g19336 (n10625, \b[41] , n1056);
  and g19337 (n10626, \b[42] , n946);
  and g19343 (n10629, n954, n6515);
  not g19346 (n_9084, n10630);
  and g19347 (n10631, \a[14] , n_9084);
  not g19348 (n_9085, n10631);
  and g19349 (n10632, \a[14] , n_9085);
  and g19350 (n10633, n_9084, n_9085);
  not g19351 (n_9086, n10632);
  not g19352 (n_9087, n10633);
  and g19353 (n10634, n_9086, n_9087);
  not g19354 (n_9088, n10634);
  and g19355 (n10635, n10623, n_9088);
  not g19356 (n_9089, n10623);
  and g19357 (n10636, n_9089, n10634);
  not g19358 (n_9090, n10355);
  not g19359 (n_9091, n10636);
  and g19360 (n10637, n_9090, n_9091);
  not g19361 (n_9092, n10635);
  and g19362 (n10638, n_9092, n10637);
  not g19363 (n_9093, n10638);
  and g19364 (n10639, n_9090, n_9093);
  and g19365 (n10640, n_9092, n_9093);
  and g19366 (n10641, n_9091, n10640);
  not g19367 (n_9094, n10639);
  not g19368 (n_9095, n10641);
  and g19369 (n10642, n_9094, n_9095);
  and g19370 (n10643, \b[46] , n700);
  and g19371 (n10644, \b[44] , n767);
  and g19372 (n10645, \b[45] , n695);
  and g19378 (n10648, n703, n7677);
  not g19381 (n_9100, n10649);
  and g19382 (n10650, \a[11] , n_9100);
  not g19383 (n_9101, n10650);
  and g19384 (n10651, \a[11] , n_9101);
  and g19385 (n10652, n_9100, n_9101);
  not g19386 (n_9102, n10651);
  not g19387 (n_9103, n10652);
  and g19388 (n10653, n_9102, n_9103);
  and g19389 (n10654, n10642, n10653);
  not g19390 (n_9104, n10642);
  not g19391 (n_9105, n10653);
  and g19392 (n10655, n_9104, n_9105);
  not g19393 (n_9106, n10654);
  not g19394 (n_9107, n10655);
  and g19395 (n10656, n_9106, n_9107);
  not g19396 (n_9108, n10354);
  and g19397 (n10657, n_9108, n10656);
  not g19398 (n_9109, n10656);
  and g19399 (n10658, n10354, n_9109);
  not g19400 (n_9110, n10657);
  not g19401 (n_9111, n10658);
  and g19402 (n10659, n_9110, n_9111);
  not g19403 (n_9112, n10659);
  and g19404 (n10660, n10353, n_9112);
  not g19405 (n_9113, n10353);
  and g19406 (n10661, n_9113, n10659);
  not g19407 (n_9114, n10660);
  not g19408 (n_9115, n10661);
  and g19409 (n10662, n_9114, n_9115);
  not g19410 (n_9116, n10342);
  and g19411 (n10663, n_9116, n10662);
  not g19412 (n_9117, n10662);
  and g19413 (n10664, n10342, n_9117);
  not g19414 (n_9118, n10663);
  not g19415 (n_9119, n10664);
  and g19416 (n10665, n_9118, n_9119);
  not g19417 (n_9120, n10341);
  and g19418 (n10666, n_9120, n10665);
  not g19419 (n_9121, n10666);
  and g19420 (n10667, n10665, n_9121);
  and g19421 (n10668, n_9120, n_9121);
  not g19422 (n_9122, n10667);
  not g19423 (n_9123, n10668);
  and g19424 (n10669, n_9122, n_9123);
  not g19425 (n_9124, n10330);
  and g19426 (n10670, n_9124, n10669);
  not g19427 (n_9125, n10669);
  and g19428 (n10671, n10330, n_9125);
  not g19429 (n_9126, n10670);
  not g19430 (n_9127, n10671);
  and g19431 (n10672, n_9126, n_9127);
  and g19432 (n10673, \b[55] , n266);
  and g19433 (n10674, \b[53] , n284);
  and g19434 (n10675, \b[54] , n261);
  and g19440 (n10678, n_8536, n_8539);
  not g19441 (n_9132, \b[55] );
  and g19442 (n10679, n_8534, n_9132);
  and g19443 (n10680, \b[54] , \b[55] );
  not g19444 (n_9133, n10679);
  not g19445 (n_9134, n10680);
  and g19446 (n10681, n_9133, n_9134);
  not g19447 (n_9135, n10678);
  and g19448 (n10682, n_9135, n10681);
  not g19449 (n_9136, n10681);
  and g19450 (n10683, n10678, n_9136);
  not g19451 (n_9137, n10682);
  not g19452 (n_9138, n10683);
  and g19453 (n10684, n_9137, n_9138);
  and g19454 (n10685, n269, n10684);
  not g19457 (n_9140, n10686);
  and g19458 (n10687, \a[2] , n_9140);
  not g19459 (n_9141, n10687);
  and g19460 (n10688, \a[2] , n_9141);
  and g19461 (n10689, n_9140, n_9141);
  not g19462 (n_9142, n10688);
  not g19463 (n_9143, n10689);
  and g19464 (n10690, n_9142, n_9143);
  not g19465 (n_9144, n10672);
  not g19466 (n_9145, n10690);
  and g19467 (n10691, n_9144, n_9145);
  and g19468 (n10692, n10672, n10690);
  not g19469 (n_9146, n10691);
  not g19470 (n_9147, n10692);
  and g19471 (n10693, n_9146, n_9147);
  not g19472 (n_9148, n10329);
  and g19473 (n10694, n_9148, n10693);
  not g19474 (n_9149, n10693);
  and g19475 (n10695, n10329, n_9149);
  not g19476 (n_9150, n10694);
  not g19477 (n_9151, n10695);
  and g19478 (\f[55] , n_9150, n_9151);
  and g19479 (n10697, \b[56] , n266);
  and g19480 (n10698, \b[54] , n284);
  and g19481 (n10699, \b[55] , n261);
  and g19487 (n10702, n_9134, n_9137);
  not g19488 (n_9156, \b[56] );
  and g19489 (n10703, n_9132, n_9156);
  and g19490 (n10704, \b[55] , \b[56] );
  not g19491 (n_9157, n10703);
  not g19492 (n_9158, n10704);
  and g19493 (n10705, n_9157, n_9158);
  not g19494 (n_9159, n10702);
  and g19495 (n10706, n_9159, n10705);
  not g19496 (n_9160, n10705);
  and g19497 (n10707, n10702, n_9160);
  not g19498 (n_9161, n10706);
  not g19499 (n_9162, n10707);
  and g19500 (n10708, n_9161, n_9162);
  and g19501 (n10709, n269, n10708);
  not g19504 (n_9164, n10710);
  and g19505 (n10711, \a[2] , n_9164);
  not g19506 (n_9165, n10711);
  and g19507 (n10712, \a[2] , n_9165);
  and g19508 (n10713, n_9164, n_9165);
  not g19509 (n_9166, n10712);
  not g19510 (n_9167, n10713);
  and g19511 (n10714, n_9166, n_9167);
  and g19512 (n10715, n_9124, n_9125);
  not g19513 (n_9168, n10715);
  and g19514 (n10716, n_9121, n_9168);
  and g19515 (n10717, n_9115, n_9118);
  and g19516 (n10718, \b[50] , n511);
  and g19517 (n10719, \b[48] , n541);
  and g19518 (n10720, \b[49] , n506);
  and g19524 (n10723, n514, n8949);
  not g19527 (n_9173, n10724);
  and g19528 (n10725, \a[8] , n_9173);
  not g19529 (n_9174, n10725);
  and g19530 (n10726, \a[8] , n_9174);
  and g19531 (n10727, n_9173, n_9174);
  not g19532 (n_9175, n10726);
  not g19533 (n_9176, n10727);
  and g19534 (n10728, n_9175, n_9176);
  and g19535 (n10729, n_9107, n_9110);
  and g19536 (n10730, \b[35] , n2048);
  and g19537 (n10731, \b[33] , n2198);
  and g19538 (n10732, \b[34] , n2043);
  and g19544 (n10735, n2051, n4696);
  not g19547 (n_9181, n10736);
  and g19548 (n10737, \a[23] , n_9181);
  not g19549 (n_9182, n10737);
  and g19550 (n10738, \a[23] , n_9182);
  and g19551 (n10739, n_9181, n_9182);
  not g19552 (n_9183, n10738);
  not g19553 (n_9184, n10739);
  and g19554 (n10740, n_9183, n_9184);
  and g19555 (n10741, n_9024, n_9030);
  and g19556 (n10742, \b[32] , n2539);
  and g19557 (n10743, \b[30] , n2685);
  and g19558 (n10744, \b[31] , n2534);
  and g19564 (n10747, n2542, n4013);
  not g19567 (n_9189, n10748);
  and g19568 (n10749, \a[26] , n_9189);
  not g19569 (n_9190, n10749);
  and g19570 (n10750, \a[26] , n_9190);
  and g19571 (n10751, n_9189, n_9190);
  not g19572 (n_9191, n10750);
  not g19573 (n_9192, n10751);
  and g19574 (n10752, n_9191, n_9192);
  and g19575 (n10753, n_9008, n_9014);
  and g19576 (n10754, n_8992, n_8998);
  and g19577 (n10755, n_8976, n_8982);
  and g19578 (n10756, n_8943, n_8949);
  and g19579 (n10757, \b[17] , n5777);
  and g19580 (n10758, \b[15] , n6059);
  and g19581 (n10759, \b[16] , n5772);
  and g19587 (n10762, n1356, n5780);
  not g19590 (n_9197, n10763);
  and g19591 (n10764, \a[41] , n_9197);
  not g19592 (n_9198, n10764);
  and g19593 (n10765, \a[41] , n_9198);
  and g19594 (n10766, n_9197, n_9198);
  not g19595 (n_9199, n10765);
  not g19596 (n_9200, n10766);
  and g19597 (n10767, n_9199, n_9200);
  and g19598 (n10768, n_8937, n_8940);
  and g19599 (n10769, \b[14] , n6595);
  and g19600 (n10770, \b[12] , n6902);
  and g19601 (n10771, \b[13] , n6590);
  and g19607 (n10774, n1034, n6598);
  not g19610 (n_9205, n10775);
  and g19611 (n10776, \a[44] , n_9205);
  not g19612 (n_9206, n10776);
  and g19613 (n10777, \a[44] , n_9206);
  and g19614 (n10778, n_9205, n_9206);
  not g19615 (n_9207, n10777);
  not g19616 (n_9208, n10778);
  and g19617 (n10779, n_9207, n_9208);
  and g19618 (n10780, n_8929, n_8932);
  and g19619 (n10781, \b[11] , n7446);
  and g19620 (n10782, \b[9] , n7787);
  and g19621 (n10783, \b[10] , n7441);
  and g19627 (n10786, n818, n7449);
  not g19630 (n_9213, n10787);
  and g19631 (n10788, \a[47] , n_9213);
  not g19632 (n_9214, n10788);
  and g19633 (n10789, \a[47] , n_9214);
  and g19634 (n10790, n_9213, n_9214);
  not g19635 (n_9215, n10789);
  not g19636 (n_9216, n10790);
  and g19637 (n10791, n_9215, n_9216);
  and g19638 (n10792, n_8921, n_8924);
  and g19639 (n10793, n_8913, n_8916);
  and g19640 (n10794, \b[2] , n10426);
  and g19641 (n10795, n10128, n_8900);
  and g19642 (n10796, n10420, n10795);
  and g19643 (n10797, \b[0] , n10796);
  and g19644 (n10798, \b[1] , n10421);
  and g19650 (n10801, n296, n10429);
  not g19653 (n_9221, n10802);
  and g19654 (n10803, \a[56] , n_9221);
  not g19655 (n_9222, n10803);
  and g19656 (n10804, \a[56] , n_9222);
  and g19657 (n10805, n_9221, n_9222);
  not g19658 (n_9223, n10804);
  not g19659 (n_9224, n10805);
  and g19660 (n10806, n_9223, n_9224);
  and g19661 (n10807, n_8908, n10806);
  not g19662 (n_9225, n10806);
  and g19663 (n10808, n10436, n_9225);
  not g19664 (n_9226, n10807);
  not g19665 (n_9227, n10808);
  and g19666 (n10809, n_9226, n_9227);
  and g19667 (n10810, \b[5] , n9339);
  and g19668 (n10811, \b[3] , n9732);
  and g19669 (n10812, \b[4] , n9334);
  and g19675 (n10815, n394, n9342);
  not g19678 (n_9232, n10816);
  and g19679 (n10817, \a[53] , n_9232);
  not g19680 (n_9233, n10817);
  and g19681 (n10818, \a[53] , n_9233);
  and g19682 (n10819, n_9232, n_9233);
  not g19683 (n_9234, n10818);
  not g19684 (n_9235, n10819);
  and g19685 (n10820, n_9234, n_9235);
  not g19686 (n_9236, n10820);
  and g19687 (n10821, n10809, n_9236);
  not g19688 (n_9237, n10809);
  and g19689 (n10822, n_9237, n10820);
  not g19690 (n_9238, n10793);
  not g19691 (n_9239, n10822);
  and g19692 (n10823, n_9238, n_9239);
  not g19693 (n_9240, n10821);
  and g19694 (n10824, n_9240, n10823);
  not g19695 (n_9241, n10824);
  and g19696 (n10825, n_9238, n_9241);
  and g19697 (n10826, n_9240, n_9241);
  and g19698 (n10827, n_9239, n10826);
  not g19699 (n_9242, n10825);
  not g19700 (n_9243, n10827);
  and g19701 (n10828, n_9242, n_9243);
  and g19702 (n10829, \b[8] , n8362);
  and g19703 (n10830, \b[6] , n8715);
  and g19704 (n10831, \b[7] , n8357);
  and g19710 (n10834, n585, n8365);
  not g19713 (n_9248, n10835);
  and g19714 (n10836, \a[50] , n_9248);
  not g19715 (n_9249, n10836);
  and g19716 (n10837, \a[50] , n_9249);
  and g19717 (n10838, n_9248, n_9249);
  not g19718 (n_9250, n10837);
  not g19719 (n_9251, n10838);
  and g19720 (n10839, n_9250, n_9251);
  and g19721 (n10840, n10828, n10839);
  not g19722 (n_9252, n10828);
  not g19723 (n_9253, n10839);
  and g19724 (n10841, n_9252, n_9253);
  not g19725 (n_9254, n10840);
  not g19726 (n_9255, n10841);
  and g19727 (n10842, n_9254, n_9255);
  not g19728 (n_9256, n10792);
  and g19729 (n10843, n_9256, n10842);
  not g19730 (n_9257, n10842);
  and g19731 (n10844, n10792, n_9257);
  not g19732 (n_9258, n10843);
  not g19733 (n_9259, n10844);
  and g19734 (n10845, n_9258, n_9259);
  not g19735 (n_9260, n10845);
  and g19736 (n10846, n10791, n_9260);
  not g19737 (n_9261, n10791);
  and g19738 (n10847, n_9261, n10845);
  not g19739 (n_9262, n10846);
  not g19740 (n_9263, n10847);
  and g19741 (n10848, n_9262, n_9263);
  not g19742 (n_9264, n10780);
  and g19743 (n10849, n_9264, n10848);
  not g19744 (n_9265, n10848);
  and g19745 (n10850, n10780, n_9265);
  not g19746 (n_9266, n10849);
  not g19747 (n_9267, n10850);
  and g19748 (n10851, n_9266, n_9267);
  not g19749 (n_9268, n10779);
  and g19750 (n10852, n_9268, n10851);
  not g19751 (n_9269, n10852);
  and g19752 (n10853, n10851, n_9269);
  and g19753 (n10854, n_9268, n_9269);
  not g19754 (n_9270, n10853);
  not g19755 (n_9271, n10854);
  and g19756 (n10855, n_9270, n_9271);
  not g19757 (n_9272, n10768);
  not g19758 (n_9273, n10855);
  and g19759 (n10856, n_9272, n_9273);
  and g19760 (n10857, n10768, n10855);
  not g19761 (n_9274, n10856);
  not g19762 (n_9275, n10857);
  and g19763 (n10858, n_9274, n_9275);
  not g19764 (n_9276, n10767);
  and g19765 (n10859, n_9276, n10858);
  not g19766 (n_9277, n10859);
  and g19767 (n10860, n_9276, n_9277);
  and g19768 (n10861, n10858, n_9277);
  not g19769 (n_9278, n10860);
  not g19770 (n_9279, n10861);
  and g19771 (n10862, n_9278, n_9279);
  not g19772 (n_9280, n10756);
  not g19773 (n_9281, n10862);
  and g19774 (n10863, n_9280, n_9281);
  not g19775 (n_9282, n10863);
  and g19776 (n10864, n_9280, n_9282);
  and g19777 (n10865, n_9281, n_9282);
  not g19778 (n_9283, n10864);
  not g19779 (n_9284, n10865);
  and g19780 (n10866, n_9283, n_9284);
  and g19781 (n10867, \b[20] , n5035);
  and g19782 (n10868, \b[18] , n5277);
  and g19783 (n10869, \b[19] , n5030);
  and g19789 (n10872, n1846, n5038);
  not g19792 (n_9289, n10873);
  and g19793 (n10874, \a[38] , n_9289);
  not g19794 (n_9290, n10874);
  and g19795 (n10875, \a[38] , n_9290);
  and g19796 (n10876, n_9289, n_9290);
  not g19797 (n_9291, n10875);
  not g19798 (n_9292, n10876);
  and g19799 (n10877, n_9291, n_9292);
  not g19800 (n_9293, n10866);
  not g19801 (n_9294, n10877);
  and g19802 (n10878, n_9293, n_9294);
  not g19803 (n_9295, n10878);
  and g19804 (n10879, n_9293, n_9295);
  and g19805 (n10880, n_9294, n_9295);
  not g19806 (n_9296, n10879);
  not g19807 (n_9297, n10880);
  and g19808 (n10881, n_9296, n_9297);
  not g19809 (n_9298, n10487);
  and g19810 (n10882, n_9298, n10881);
  not g19811 (n_9299, n10881);
  and g19812 (n10883, n10487, n_9299);
  not g19813 (n_9300, n10882);
  not g19814 (n_9301, n10883);
  and g19815 (n10884, n_9300, n_9301);
  and g19816 (n10885, \b[23] , n4287);
  and g19817 (n10886, \b[21] , n4532);
  and g19818 (n10887, \b[22] , n4282);
  and g19824 (n10890, n2300, n4290);
  not g19827 (n_9306, n10891);
  and g19828 (n10892, \a[35] , n_9306);
  not g19829 (n_9307, n10892);
  and g19830 (n10893, \a[35] , n_9307);
  and g19831 (n10894, n_9306, n_9307);
  not g19832 (n_9308, n10893);
  not g19833 (n_9309, n10894);
  and g19834 (n10895, n_9308, n_9309);
  not g19835 (n_9310, n10884);
  not g19836 (n_9311, n10895);
  and g19837 (n10896, n_9310, n_9311);
  and g19838 (n10897, n10884, n10895);
  not g19839 (n_9312, n10896);
  not g19840 (n_9313, n10897);
  and g19841 (n10898, n_9312, n_9313);
  not g19842 (n_9314, n10898);
  and g19843 (n10899, n10755, n_9314);
  not g19844 (n_9315, n10755);
  and g19845 (n10900, n_9315, n10898);
  not g19846 (n_9316, n10899);
  not g19847 (n_9317, n10900);
  and g19848 (n10901, n_9316, n_9317);
  and g19849 (n10902, \b[26] , n3638);
  and g19850 (n10903, \b[24] , n3843);
  and g19851 (n10904, \b[25] , n3633);
  and g19857 (n10907, n2813, n3641);
  not g19860 (n_9322, n10908);
  and g19861 (n10909, \a[32] , n_9322);
  not g19862 (n_9323, n10909);
  and g19863 (n10910, \a[32] , n_9323);
  and g19864 (n10911, n_9322, n_9323);
  not g19865 (n_9324, n10910);
  not g19866 (n_9325, n10911);
  and g19867 (n10912, n_9324, n_9325);
  not g19868 (n_9326, n10912);
  and g19869 (n10913, n10901, n_9326);
  not g19870 (n_9327, n10901);
  and g19871 (n10914, n_9327, n10912);
  not g19872 (n_9328, n10754);
  not g19873 (n_9329, n10914);
  and g19874 (n10915, n_9328, n_9329);
  not g19875 (n_9330, n10913);
  and g19876 (n10916, n_9330, n10915);
  not g19877 (n_9331, n10916);
  and g19878 (n10917, n_9328, n_9331);
  and g19879 (n10918, n_9330, n_9331);
  and g19880 (n10919, n_9329, n10918);
  not g19881 (n_9332, n10917);
  not g19882 (n_9333, n10919);
  and g19883 (n10920, n_9332, n_9333);
  and g19884 (n10921, \b[29] , n3050);
  and g19885 (n10922, \b[27] , n3243);
  and g19886 (n10923, \b[28] , n3045);
  and g19892 (n10926, n3053, n3383);
  not g19895 (n_9338, n10927);
  and g19896 (n10928, \a[29] , n_9338);
  not g19897 (n_9339, n10928);
  and g19898 (n10929, \a[29] , n_9339);
  and g19899 (n10930, n_9338, n_9339);
  not g19900 (n_9340, n10929);
  not g19901 (n_9341, n10930);
  and g19902 (n10931, n_9340, n_9341);
  and g19903 (n10932, n10920, n10931);
  not g19904 (n_9342, n10920);
  not g19905 (n_9343, n10931);
  and g19906 (n10933, n_9342, n_9343);
  not g19907 (n_9344, n10932);
  not g19908 (n_9345, n10933);
  and g19909 (n10934, n_9344, n_9345);
  not g19910 (n_9346, n10753);
  and g19911 (n10935, n_9346, n10934);
  not g19912 (n_9347, n10934);
  and g19913 (n10936, n10753, n_9347);
  not g19914 (n_9348, n10935);
  not g19915 (n_9349, n10936);
  and g19916 (n10937, n_9348, n_9349);
  not g19917 (n_9350, n10937);
  and g19918 (n10938, n10752, n_9350);
  not g19919 (n_9351, n10752);
  and g19920 (n10939, n_9351, n10937);
  not g19921 (n_9352, n10938);
  not g19922 (n_9353, n10939);
  and g19923 (n10940, n_9352, n_9353);
  not g19924 (n_9354, n10741);
  and g19925 (n10941, n_9354, n10940);
  not g19926 (n_9355, n10940);
  and g19927 (n10942, n10741, n_9355);
  not g19928 (n_9356, n10941);
  not g19929 (n_9357, n10942);
  and g19930 (n10943, n_9356, n_9357);
  not g19931 (n_9358, n10740);
  and g19932 (n10944, n_9358, n10943);
  not g19933 (n_9359, n10944);
  and g19934 (n10945, n10943, n_9359);
  and g19935 (n10946, n_9358, n_9359);
  not g19936 (n_9360, n10945);
  not g19937 (n_9361, n10946);
  and g19938 (n10947, n_9360, n_9361);
  and g19939 (n10948, n_9040, n_9047);
  and g19940 (n10949, n10947, n10948);
  not g19941 (n_9362, n10947);
  not g19942 (n_9363, n10948);
  and g19943 (n10950, n_9362, n_9363);
  not g19944 (n_9364, n10949);
  not g19945 (n_9365, n10950);
  and g19946 (n10951, n_9364, n_9365);
  and g19947 (n10952, \b[38] , n1627);
  and g19948 (n10953, \b[36] , n1763);
  and g19949 (n10954, \b[37] , n1622);
  and g19955 (n10957, n1630, n5205);
  not g19958 (n_9370, n10958);
  and g19959 (n10959, \a[20] , n_9370);
  not g19960 (n_9371, n10959);
  and g19961 (n10960, \a[20] , n_9371);
  and g19962 (n10961, n_9370, n_9371);
  not g19963 (n_9372, n10960);
  not g19964 (n_9373, n10961);
  and g19965 (n10962, n_9372, n_9373);
  not g19966 (n_9374, n10962);
  and g19967 (n10963, n10951, n_9374);
  not g19968 (n_9375, n10963);
  and g19969 (n10964, n10951, n_9375);
  and g19970 (n10965, n_9374, n_9375);
  not g19971 (n_9376, n10964);
  not g19972 (n_9377, n10965);
  and g19973 (n10966, n_9376, n_9377);
  and g19974 (n10967, n_9057, n_9063);
  and g19975 (n10968, n10966, n10967);
  not g19976 (n_9378, n10966);
  not g19977 (n_9379, n10967);
  and g19978 (n10969, n_9378, n_9379);
  not g19979 (n_9380, n10968);
  not g19980 (n_9381, n10969);
  and g19981 (n10970, n_9380, n_9381);
  and g19982 (n10971, \b[41] , n1302);
  and g19983 (n10972, \b[39] , n1391);
  and g19984 (n10973, \b[40] , n1297);
  and g19990 (n10976, n1305, n6219);
  not g19993 (n_9386, n10977);
  and g19994 (n10978, \a[17] , n_9386);
  not g19995 (n_9387, n10978);
  and g19996 (n10979, \a[17] , n_9387);
  and g19997 (n10980, n_9386, n_9387);
  not g19998 (n_9388, n10979);
  not g19999 (n_9389, n10980);
  and g20000 (n10981, n_9388, n_9389);
  not g20001 (n_9390, n10981);
  and g20002 (n10982, n10970, n_9390);
  not g20003 (n_9391, n10982);
  and g20004 (n10983, n10970, n_9391);
  and g20005 (n10984, n_9390, n_9391);
  not g20006 (n_9392, n10983);
  not g20007 (n_9393, n10984);
  and g20008 (n10985, n_9392, n_9393);
  and g20009 (n10986, n_9073, n_9079);
  and g20010 (n10987, n10985, n10986);
  not g20011 (n_9394, n10985);
  not g20012 (n_9395, n10986);
  and g20013 (n10988, n_9394, n_9395);
  not g20014 (n_9396, n10987);
  not g20015 (n_9397, n10988);
  and g20016 (n10989, n_9396, n_9397);
  and g20017 (n10990, \b[44] , n951);
  and g20018 (n10991, \b[42] , n1056);
  and g20019 (n10992, \b[43] , n946);
  and g20025 (n10995, n954, n7072);
  not g20028 (n_9402, n10996);
  and g20029 (n10997, \a[14] , n_9402);
  not g20030 (n_9403, n10997);
  and g20031 (n10998, \a[14] , n_9403);
  and g20032 (n10999, n_9402, n_9403);
  not g20033 (n_9404, n10998);
  not g20034 (n_9405, n10999);
  and g20035 (n11000, n_9404, n_9405);
  not g20036 (n_9406, n11000);
  and g20037 (n11001, n10989, n_9406);
  not g20038 (n_9407, n10989);
  and g20039 (n11002, n_9407, n11000);
  not g20040 (n_9408, n10640);
  not g20041 (n_9409, n11002);
  and g20042 (n11003, n_9408, n_9409);
  not g20043 (n_9410, n11001);
  and g20044 (n11004, n_9410, n11003);
  not g20045 (n_9411, n11004);
  and g20046 (n11005, n_9408, n_9411);
  and g20047 (n11006, n_9410, n_9411);
  and g20048 (n11007, n_9409, n11006);
  not g20049 (n_9412, n11005);
  not g20050 (n_9413, n11007);
  and g20051 (n11008, n_9412, n_9413);
  and g20052 (n11009, \b[47] , n700);
  and g20053 (n11010, \b[45] , n767);
  and g20054 (n11011, \b[46] , n695);
  and g20060 (n11014, n703, n7703);
  not g20063 (n_9418, n11015);
  and g20064 (n11016, \a[11] , n_9418);
  not g20065 (n_9419, n11016);
  and g20066 (n11017, \a[11] , n_9419);
  and g20067 (n11018, n_9418, n_9419);
  not g20068 (n_9420, n11017);
  not g20069 (n_9421, n11018);
  and g20070 (n11019, n_9420, n_9421);
  not g20071 (n_9422, n11008);
  not g20072 (n_9423, n11019);
  and g20073 (n11020, n_9422, n_9423);
  not g20074 (n_9424, n11020);
  and g20075 (n11021, n_9422, n_9424);
  and g20076 (n11022, n_9423, n_9424);
  not g20077 (n_9425, n11021);
  not g20078 (n_9426, n11022);
  and g20079 (n11023, n_9425, n_9426);
  not g20080 (n_9427, n10729);
  not g20081 (n_9428, n11023);
  and g20082 (n11024, n_9427, n_9428);
  and g20083 (n11025, n10729, n11023);
  not g20084 (n_9429, n11024);
  not g20085 (n_9430, n11025);
  and g20086 (n11026, n_9429, n_9430);
  not g20087 (n_9431, n10728);
  and g20088 (n11027, n_9431, n11026);
  not g20089 (n_9432, n11027);
  and g20090 (n11028, n_9431, n_9432);
  and g20091 (n11029, n11026, n_9432);
  not g20092 (n_9433, n11028);
  not g20093 (n_9434, n11029);
  and g20094 (n11030, n_9433, n_9434);
  not g20095 (n_9435, n10717);
  not g20096 (n_9436, n11030);
  and g20097 (n11031, n_9435, n_9436);
  not g20098 (n_9437, n11031);
  and g20099 (n11032, n_9435, n_9437);
  and g20100 (n11033, n_9436, n_9437);
  not g20101 (n_9438, n11032);
  not g20102 (n_9439, n11033);
  and g20103 (n11034, n_9438, n_9439);
  and g20104 (n11035, \b[53] , n362);
  and g20105 (n11036, \b[51] , n403);
  and g20106 (n11037, \b[52] , n357);
  and g20112 (n11040, n365, n9972);
  not g20115 (n_9444, n11041);
  and g20116 (n11042, \a[5] , n_9444);
  not g20117 (n_9445, n11042);
  and g20118 (n11043, \a[5] , n_9445);
  and g20119 (n11044, n_9444, n_9445);
  not g20120 (n_9446, n11043);
  not g20121 (n_9447, n11044);
  and g20122 (n11045, n_9446, n_9447);
  and g20123 (n11046, n11034, n11045);
  not g20124 (n_9448, n11034);
  not g20125 (n_9449, n11045);
  and g20126 (n11047, n_9448, n_9449);
  not g20127 (n_9450, n11046);
  not g20128 (n_9451, n11047);
  and g20129 (n11048, n_9450, n_9451);
  not g20130 (n_9452, n10716);
  and g20131 (n11049, n_9452, n11048);
  not g20132 (n_9453, n11048);
  and g20133 (n11050, n10716, n_9453);
  not g20134 (n_9454, n11049);
  not g20135 (n_9455, n11050);
  and g20136 (n11051, n_9454, n_9455);
  not g20137 (n_9456, n10714);
  and g20138 (n11052, n_9456, n11051);
  not g20139 (n_9457, n11052);
  and g20140 (n11053, n11051, n_9457);
  and g20141 (n11054, n_9456, n_9457);
  not g20142 (n_9458, n11053);
  not g20143 (n_9459, n11054);
  and g20144 (n11055, n_9458, n_9459);
  and g20145 (n11056, n_9146, n_9150);
  not g20146 (n_9460, n11055);
  not g20147 (n_9461, n11056);
  and g20148 (n11057, n_9460, n_9461);
  and g20149 (n11058, n11055, n11056);
  not g20150 (n_9462, n11057);
  not g20151 (n_9463, n11058);
  and g20152 (\f[56] , n_9462, n_9463);
  and g20153 (n11060, n_9451, n_9454);
  and g20154 (n11061, \b[54] , n362);
  and g20155 (n11062, \b[52] , n403);
  and g20156 (n11063, \b[53] , n357);
  and g20162 (n11066, n365, n9998);
  not g20165 (n_9468, n11067);
  and g20166 (n11068, \a[5] , n_9468);
  not g20167 (n_9469, n11068);
  and g20168 (n11069, \a[5] , n_9469);
  and g20169 (n11070, n_9468, n_9469);
  not g20170 (n_9470, n11069);
  not g20171 (n_9471, n11070);
  and g20172 (n11071, n_9470, n_9471);
  and g20173 (n11072, n_9432, n_9437);
  and g20174 (n11073, \b[51] , n511);
  and g20175 (n11074, \b[49] , n541);
  and g20176 (n11075, \b[50] , n506);
  and g20182 (n11078, n514, n8976);
  not g20185 (n_9476, n11079);
  and g20186 (n11080, \a[8] , n_9476);
  not g20187 (n_9477, n11080);
  and g20188 (n11081, \a[8] , n_9477);
  and g20189 (n11082, n_9476, n_9477);
  not g20190 (n_9478, n11081);
  not g20191 (n_9479, n11082);
  and g20192 (n11083, n_9478, n_9479);
  and g20193 (n11084, n_9424, n_9429);
  and g20194 (n11085, \b[48] , n700);
  and g20195 (n11086, \b[46] , n767);
  and g20196 (n11087, \b[47] , n695);
  and g20202 (n11090, n703, n8009);
  not g20205 (n_9484, n11091);
  and g20206 (n11092, \a[11] , n_9484);
  not g20207 (n_9485, n11092);
  and g20208 (n11093, \a[11] , n_9485);
  and g20209 (n11094, n_9484, n_9485);
  not g20210 (n_9486, n11093);
  not g20211 (n_9487, n11094);
  and g20212 (n11095, n_9486, n_9487);
  and g20213 (n11096, \b[45] , n951);
  and g20214 (n11097, \b[43] , n1056);
  and g20215 (n11098, \b[44] , n946);
  and g20221 (n11101, n954, n7361);
  not g20224 (n_9492, n11102);
  and g20225 (n11103, \a[14] , n_9492);
  not g20226 (n_9493, n11103);
  and g20227 (n11104, \a[14] , n_9493);
  and g20228 (n11105, n_9492, n_9493);
  not g20229 (n_9494, n11104);
  not g20230 (n_9495, n11105);
  and g20231 (n11106, n_9494, n_9495);
  and g20232 (n11107, n_9391, n_9397);
  and g20233 (n11108, n_9359, n_9365);
  and g20234 (n11109, n_9353, n_9356);
  and g20235 (n11110, n_9345, n_9348);
  and g20236 (n11111, \b[30] , n3050);
  and g20237 (n11112, \b[28] , n3243);
  and g20238 (n11113, \b[29] , n3045);
  and g20244 (n11116, n3053, n3577);
  not g20247 (n_9500, n11117);
  and g20248 (n11118, \a[29] , n_9500);
  not g20249 (n_9501, n11118);
  and g20250 (n11119, \a[29] , n_9501);
  and g20251 (n11120, n_9500, n_9501);
  not g20252 (n_9502, n11119);
  not g20253 (n_9503, n11120);
  and g20254 (n11121, n_9502, n_9503);
  and g20255 (n11122, n_9298, n_9299);
  not g20256 (n_9504, n11122);
  and g20257 (n11123, n_9295, n_9504);
  and g20258 (n11124, \b[21] , n5035);
  and g20259 (n11125, \b[19] , n5277);
  and g20260 (n11126, \b[20] , n5030);
  and g20266 (n11129, n1984, n5038);
  not g20269 (n_9509, n11130);
  and g20270 (n11131, \a[38] , n_9509);
  not g20271 (n_9510, n11131);
  and g20272 (n11132, \a[38] , n_9510);
  and g20273 (n11133, n_9509, n_9510);
  not g20274 (n_9511, n11132);
  not g20275 (n_9512, n11133);
  and g20276 (n11134, n_9511, n_9512);
  and g20277 (n11135, n_9277, n_9282);
  and g20278 (n11136, \b[18] , n5777);
  and g20279 (n11137, \b[16] , n6059);
  and g20280 (n11138, \b[17] , n5772);
  and g20286 (n11141, n1566, n5780);
  not g20289 (n_9517, n11142);
  and g20290 (n11143, \a[41] , n_9517);
  not g20291 (n_9518, n11143);
  and g20292 (n11144, \a[41] , n_9518);
  and g20293 (n11145, n_9517, n_9518);
  not g20294 (n_9519, n11144);
  not g20295 (n_9520, n11145);
  and g20296 (n11146, n_9519, n_9520);
  and g20297 (n11147, n_9269, n_9274);
  and g20298 (n11148, \b[15] , n6595);
  and g20299 (n11149, \b[13] , n6902);
  and g20300 (n11150, \b[14] , n6590);
  and g20306 (n11153, n1131, n6598);
  not g20309 (n_9525, n11154);
  and g20310 (n11155, \a[44] , n_9525);
  not g20311 (n_9526, n11155);
  and g20312 (n11156, \a[44] , n_9526);
  and g20313 (n11157, n_9525, n_9526);
  not g20314 (n_9527, n11156);
  not g20315 (n_9528, n11157);
  and g20316 (n11158, n_9527, n_9528);
  and g20317 (n11159, n_9263, n_9266);
  and g20318 (n11160, \b[12] , n7446);
  and g20319 (n11161, \b[10] , n7787);
  and g20320 (n11162, \b[11] , n7441);
  and g20326 (n11165, n842, n7449);
  not g20329 (n_9533, n11166);
  and g20330 (n11167, \a[47] , n_9533);
  not g20331 (n_9534, n11167);
  and g20332 (n11168, \a[47] , n_9534);
  and g20333 (n11169, n_9533, n_9534);
  not g20334 (n_9535, n11168);
  not g20335 (n_9536, n11169);
  and g20336 (n11170, n_9535, n_9536);
  and g20337 (n11171, n_9255, n_9258);
  and g20338 (n11172, \b[6] , n9339);
  and g20339 (n11173, \b[4] , n9732);
  and g20340 (n11174, \b[5] , n9334);
  and g20346 (n11177, n459, n9342);
  not g20349 (n_9541, n11178);
  and g20350 (n11179, \a[53] , n_9541);
  not g20351 (n_9542, n11179);
  and g20352 (n11180, \a[53] , n_9542);
  and g20353 (n11181, n_9541, n_9542);
  not g20354 (n_9543, n11180);
  not g20355 (n_9544, n11181);
  and g20356 (n11182, n_9543, n_9544);
  not g20357 (n_9546, \a[57] );
  and g20358 (n11183, \a[56] , n_9546);
  and g20359 (n11184, n_8895, \a[57] );
  not g20360 (n_9547, n11183);
  not g20361 (n_9548, n11184);
  and g20362 (n11185, n_9547, n_9548);
  not g20363 (n_9549, n11185);
  and g20364 (n11186, \b[0] , n_9549);
  and g20365 (n11187, n_9227, n11186);
  not g20366 (n_9550, n11186);
  and g20367 (n11188, n10808, n_9550);
  not g20368 (n_9551, n11187);
  not g20369 (n_9552, n11188);
  and g20370 (n11189, n_9551, n_9552);
  and g20371 (n11190, \b[3] , n10426);
  and g20372 (n11191, \b[1] , n10796);
  and g20373 (n11192, \b[2] , n10421);
  and g20379 (n11195, n318, n10429);
  not g20382 (n_9557, n11196);
  and g20383 (n11197, \a[56] , n_9557);
  not g20384 (n_9558, n11197);
  and g20385 (n11198, \a[56] , n_9558);
  and g20386 (n11199, n_9557, n_9558);
  not g20387 (n_9559, n11198);
  not g20388 (n_9560, n11199);
  and g20389 (n11200, n_9559, n_9560);
  not g20390 (n_9561, n11189);
  not g20391 (n_9562, n11200);
  and g20392 (n11201, n_9561, n_9562);
  and g20393 (n11202, n11189, n11200);
  not g20394 (n_9563, n11201);
  not g20395 (n_9564, n11202);
  and g20396 (n11203, n_9563, n_9564);
  not g20397 (n_9565, n11182);
  and g20398 (n11204, n_9565, n11203);
  not g20399 (n_9566, n11204);
  and g20400 (n11205, n11203, n_9566);
  and g20401 (n11206, n_9565, n_9566);
  not g20402 (n_9567, n11205);
  not g20403 (n_9568, n11206);
  and g20404 (n11207, n_9567, n_9568);
  not g20405 (n_9569, n10826);
  and g20406 (n11208, n_9569, n11207);
  not g20407 (n_9570, n11207);
  and g20408 (n11209, n10826, n_9570);
  not g20409 (n_9571, n11208);
  not g20410 (n_9572, n11209);
  and g20411 (n11210, n_9571, n_9572);
  and g20412 (n11211, \b[9] , n8362);
  and g20413 (n11212, \b[7] , n8715);
  and g20414 (n11213, \b[8] , n8357);
  and g20420 (n11216, n651, n8365);
  not g20423 (n_9577, n11217);
  and g20424 (n11218, \a[50] , n_9577);
  not g20425 (n_9578, n11218);
  and g20426 (n11219, \a[50] , n_9578);
  and g20427 (n11220, n_9577, n_9578);
  not g20428 (n_9579, n11219);
  not g20429 (n_9580, n11220);
  and g20430 (n11221, n_9579, n_9580);
  not g20431 (n_9581, n11210);
  not g20432 (n_9582, n11221);
  and g20433 (n11222, n_9581, n_9582);
  and g20434 (n11223, n11210, n11221);
  not g20435 (n_9583, n11222);
  not g20436 (n_9584, n11223);
  and g20437 (n11224, n_9583, n_9584);
  not g20438 (n_9585, n11171);
  and g20439 (n11225, n_9585, n11224);
  not g20440 (n_9586, n11224);
  and g20441 (n11226, n11171, n_9586);
  not g20442 (n_9587, n11225);
  not g20443 (n_9588, n11226);
  and g20444 (n11227, n_9587, n_9588);
  not g20445 (n_9589, n11227);
  and g20446 (n11228, n11170, n_9589);
  not g20447 (n_9590, n11170);
  and g20448 (n11229, n_9590, n11227);
  not g20449 (n_9591, n11228);
  not g20450 (n_9592, n11229);
  and g20451 (n11230, n_9591, n_9592);
  not g20452 (n_9593, n11159);
  and g20453 (n11231, n_9593, n11230);
  not g20454 (n_9594, n11230);
  and g20455 (n11232, n11159, n_9594);
  not g20456 (n_9595, n11231);
  not g20457 (n_9596, n11232);
  and g20458 (n11233, n_9595, n_9596);
  not g20459 (n_9597, n11158);
  and g20460 (n11234, n_9597, n11233);
  not g20461 (n_9598, n11233);
  and g20462 (n11235, n11158, n_9598);
  not g20463 (n_9599, n11234);
  not g20464 (n_9600, n11235);
  and g20465 (n11236, n_9599, n_9600);
  not g20466 (n_9601, n11147);
  and g20467 (n11237, n_9601, n11236);
  not g20468 (n_9602, n11236);
  and g20469 (n11238, n11147, n_9602);
  not g20470 (n_9603, n11237);
  not g20471 (n_9604, n11238);
  and g20472 (n11239, n_9603, n_9604);
  not g20473 (n_9605, n11146);
  and g20474 (n11240, n_9605, n11239);
  not g20475 (n_9606, n11240);
  and g20476 (n11241, n_9605, n_9606);
  and g20477 (n11242, n11239, n_9606);
  not g20478 (n_9607, n11241);
  not g20479 (n_9608, n11242);
  and g20480 (n11243, n_9607, n_9608);
  not g20481 (n_9609, n11135);
  not g20482 (n_9610, n11243);
  and g20483 (n11244, n_9609, n_9610);
  and g20484 (n11245, n11135, n_9608);
  and g20485 (n11246, n_9607, n11245);
  not g20486 (n_9611, n11244);
  not g20487 (n_9612, n11246);
  and g20488 (n11247, n_9611, n_9612);
  not g20489 (n_9613, n11134);
  and g20490 (n11248, n_9613, n11247);
  not g20491 (n_9614, n11247);
  and g20492 (n11249, n11134, n_9614);
  not g20493 (n_9615, n11248);
  not g20494 (n_9616, n11249);
  and g20495 (n11250, n_9615, n_9616);
  not g20496 (n_9617, n11123);
  and g20497 (n11251, n_9617, n11250);
  not g20498 (n_9618, n11250);
  and g20499 (n11252, n11123, n_9618);
  not g20500 (n_9619, n11251);
  not g20501 (n_9620, n11252);
  and g20502 (n11253, n_9619, n_9620);
  and g20503 (n11254, \b[24] , n4287);
  and g20504 (n11255, \b[22] , n4532);
  and g20505 (n11256, \b[23] , n4282);
  and g20511 (n11259, n2458, n4290);
  not g20514 (n_9625, n11260);
  and g20515 (n11261, \a[35] , n_9625);
  not g20516 (n_9626, n11261);
  and g20517 (n11262, \a[35] , n_9626);
  and g20518 (n11263, n_9625, n_9626);
  not g20519 (n_9627, n11262);
  not g20520 (n_9628, n11263);
  and g20521 (n11264, n_9627, n_9628);
  not g20522 (n_9629, n11264);
  and g20523 (n11265, n11253, n_9629);
  not g20524 (n_9630, n11265);
  and g20525 (n11266, n11253, n_9630);
  and g20526 (n11267, n_9629, n_9630);
  not g20527 (n_9631, n11266);
  not g20528 (n_9632, n11267);
  and g20529 (n11268, n_9631, n_9632);
  and g20530 (n11269, n_9312, n_9317);
  and g20531 (n11270, n11268, n11269);
  not g20532 (n_9633, n11268);
  not g20533 (n_9634, n11269);
  and g20534 (n11271, n_9633, n_9634);
  not g20535 (n_9635, n11270);
  not g20536 (n_9636, n11271);
  and g20537 (n11272, n_9635, n_9636);
  and g20538 (n11273, \b[27] , n3638);
  and g20539 (n11274, \b[25] , n3843);
  and g20540 (n11275, \b[26] , n3633);
  and g20546 (n11278, n2990, n3641);
  not g20549 (n_9641, n11279);
  and g20550 (n11280, \a[32] , n_9641);
  not g20551 (n_9642, n11280);
  and g20552 (n11281, \a[32] , n_9642);
  and g20553 (n11282, n_9641, n_9642);
  not g20554 (n_9643, n11281);
  not g20555 (n_9644, n11282);
  and g20556 (n11283, n_9643, n_9644);
  not g20557 (n_9645, n11272);
  and g20558 (n11284, n_9645, n11283);
  not g20559 (n_9646, n11283);
  and g20560 (n11285, n11272, n_9646);
  not g20561 (n_9647, n11284);
  not g20562 (n_9648, n11285);
  and g20563 (n11286, n_9647, n_9648);
  not g20564 (n_9649, n10918);
  and g20565 (n11287, n_9649, n11286);
  not g20566 (n_9650, n11286);
  and g20567 (n11288, n10918, n_9650);
  not g20568 (n_9651, n11287);
  not g20569 (n_9652, n11288);
  and g20570 (n11289, n_9651, n_9652);
  not g20571 (n_9653, n11121);
  and g20572 (n11290, n_9653, n11289);
  not g20573 (n_9654, n11289);
  and g20574 (n11291, n11121, n_9654);
  not g20575 (n_9655, n11290);
  not g20576 (n_9656, n11291);
  and g20577 (n11292, n_9655, n_9656);
  not g20578 (n_9657, n11110);
  and g20579 (n11293, n_9657, n11292);
  not g20580 (n_9658, n11292);
  and g20581 (n11294, n11110, n_9658);
  not g20582 (n_9659, n11293);
  not g20583 (n_9660, n11294);
  and g20584 (n11295, n_9659, n_9660);
  and g20585 (n11296, \b[33] , n2539);
  and g20586 (n11297, \b[31] , n2685);
  and g20587 (n11298, \b[32] , n2534);
  and g20593 (n11301, n2542, n4223);
  not g20596 (n_9665, n11302);
  and g20597 (n11303, \a[26] , n_9665);
  not g20598 (n_9666, n11303);
  and g20599 (n11304, \a[26] , n_9666);
  and g20600 (n11305, n_9665, n_9666);
  not g20601 (n_9667, n11304);
  not g20602 (n_9668, n11305);
  and g20603 (n11306, n_9667, n_9668);
  not g20604 (n_9669, n11306);
  and g20605 (n11307, n11295, n_9669);
  not g20606 (n_9670, n11307);
  and g20607 (n11308, n11295, n_9670);
  and g20608 (n11309, n_9669, n_9670);
  not g20609 (n_9671, n11308);
  not g20610 (n_9672, n11309);
  and g20611 (n11310, n_9671, n_9672);
  not g20612 (n_9673, n11109);
  and g20613 (n11311, n_9673, n11310);
  not g20614 (n_9674, n11310);
  and g20615 (n11312, n11109, n_9674);
  not g20616 (n_9675, n11311);
  not g20617 (n_9676, n11312);
  and g20618 (n11313, n_9675, n_9676);
  and g20619 (n11314, \b[36] , n2048);
  and g20620 (n11315, \b[34] , n2198);
  and g20621 (n11316, \b[35] , n2043);
  and g20627 (n11319, n2051, n4922);
  not g20630 (n_9681, n11320);
  and g20631 (n11321, \a[23] , n_9681);
  not g20632 (n_9682, n11321);
  and g20633 (n11322, \a[23] , n_9682);
  and g20634 (n11323, n_9681, n_9682);
  not g20635 (n_9683, n11322);
  not g20636 (n_9684, n11323);
  and g20637 (n11324, n_9683, n_9684);
  not g20638 (n_9685, n11313);
  not g20639 (n_9686, n11324);
  and g20640 (n11325, n_9685, n_9686);
  and g20641 (n11326, n11313, n11324);
  not g20642 (n_9687, n11325);
  not g20643 (n_9688, n11326);
  and g20644 (n11327, n_9687, n_9688);
  not g20645 (n_9689, n11327);
  and g20646 (n11328, n11108, n_9689);
  not g20647 (n_9690, n11108);
  and g20648 (n11329, n_9690, n11327);
  not g20649 (n_9691, n11328);
  not g20650 (n_9692, n11329);
  and g20651 (n11330, n_9691, n_9692);
  and g20652 (n11331, \b[39] , n1627);
  and g20653 (n11332, \b[37] , n1763);
  and g20654 (n11333, \b[38] , n1622);
  and g20660 (n11336, n1630, n5451);
  not g20663 (n_9697, n11337);
  and g20664 (n11338, \a[20] , n_9697);
  not g20665 (n_9698, n11338);
  and g20666 (n11339, \a[20] , n_9698);
  and g20667 (n11340, n_9697, n_9698);
  not g20668 (n_9699, n11339);
  not g20669 (n_9700, n11340);
  and g20670 (n11341, n_9699, n_9700);
  not g20671 (n_9701, n11341);
  and g20672 (n11342, n11330, n_9701);
  not g20673 (n_9702, n11342);
  and g20674 (n11343, n11330, n_9702);
  and g20675 (n11344, n_9701, n_9702);
  not g20676 (n_9703, n11343);
  not g20677 (n_9704, n11344);
  and g20678 (n11345, n_9703, n_9704);
  and g20679 (n11346, n_9375, n_9381);
  and g20680 (n11347, n11345, n11346);
  not g20681 (n_9705, n11345);
  not g20682 (n_9706, n11346);
  and g20683 (n11348, n_9705, n_9706);
  not g20684 (n_9707, n11347);
  not g20685 (n_9708, n11348);
  and g20686 (n11349, n_9707, n_9708);
  and g20687 (n11350, \b[42] , n1302);
  and g20688 (n11351, \b[40] , n1391);
  and g20689 (n11352, \b[41] , n1297);
  and g20695 (n11355, n1305, n6489);
  not g20698 (n_9713, n11356);
  and g20699 (n11357, \a[17] , n_9713);
  not g20700 (n_9714, n11357);
  and g20701 (n11358, \a[17] , n_9714);
  and g20702 (n11359, n_9713, n_9714);
  not g20703 (n_9715, n11358);
  not g20704 (n_9716, n11359);
  and g20705 (n11360, n_9715, n_9716);
  not g20706 (n_9717, n11349);
  and g20707 (n11361, n_9717, n11360);
  not g20708 (n_9718, n11360);
  and g20709 (n11362, n11349, n_9718);
  not g20710 (n_9719, n11361);
  not g20711 (n_9720, n11362);
  and g20712 (n11363, n_9719, n_9720);
  not g20713 (n_9721, n11107);
  and g20714 (n11364, n_9721, n11363);
  not g20715 (n_9722, n11363);
  and g20716 (n11365, n11107, n_9722);
  not g20717 (n_9723, n11364);
  not g20718 (n_9724, n11365);
  and g20719 (n11366, n_9723, n_9724);
  not g20720 (n_9725, n11106);
  and g20721 (n11367, n_9725, n11366);
  not g20722 (n_9726, n11367);
  and g20723 (n11368, n_9725, n_9726);
  and g20724 (n11369, n11366, n_9726);
  not g20725 (n_9727, n11368);
  not g20726 (n_9728, n11369);
  and g20727 (n11370, n_9727, n_9728);
  not g20728 (n_9729, n11006);
  not g20729 (n_9730, n11370);
  and g20730 (n11371, n_9729, n_9730);
  and g20731 (n11372, n11006, n_9728);
  and g20732 (n11373, n_9727, n11372);
  not g20733 (n_9731, n11371);
  not g20734 (n_9732, n11373);
  and g20735 (n11374, n_9731, n_9732);
  not g20736 (n_9733, n11095);
  and g20737 (n11375, n_9733, n11374);
  not g20738 (n_9734, n11375);
  and g20739 (n11376, n_9733, n_9734);
  and g20740 (n11377, n11374, n_9734);
  not g20741 (n_9735, n11376);
  not g20742 (n_9736, n11377);
  and g20743 (n11378, n_9735, n_9736);
  not g20744 (n_9737, n11084);
  not g20745 (n_9738, n11378);
  and g20746 (n11379, n_9737, n_9738);
  and g20747 (n11380, n11084, n_9736);
  and g20748 (n11381, n_9735, n11380);
  not g20749 (n_9739, n11379);
  not g20750 (n_9740, n11381);
  and g20751 (n11382, n_9739, n_9740);
  not g20752 (n_9741, n11083);
  and g20753 (n11383, n_9741, n11382);
  not g20754 (n_9742, n11383);
  and g20755 (n11384, n_9741, n_9742);
  and g20756 (n11385, n11382, n_9742);
  not g20757 (n_9743, n11384);
  not g20758 (n_9744, n11385);
  and g20759 (n11386, n_9743, n_9744);
  not g20760 (n_9745, n11072);
  not g20761 (n_9746, n11386);
  and g20762 (n11387, n_9745, n_9746);
  and g20763 (n11388, n11072, n_9744);
  and g20764 (n11389, n_9743, n11388);
  not g20765 (n_9747, n11387);
  not g20766 (n_9748, n11389);
  and g20767 (n11390, n_9747, n_9748);
  not g20768 (n_9749, n11071);
  and g20769 (n11391, n_9749, n11390);
  not g20770 (n_9750, n11391);
  and g20771 (n11392, n_9749, n_9750);
  and g20772 (n11393, n11390, n_9750);
  not g20773 (n_9751, n11392);
  not g20774 (n_9752, n11393);
  and g20775 (n11394, n_9751, n_9752);
  not g20776 (n_9753, n11060);
  not g20777 (n_9754, n11394);
  and g20778 (n11395, n_9753, n_9754);
  not g20779 (n_9755, n11395);
  and g20780 (n11396, n_9753, n_9755);
  and g20781 (n11397, n_9754, n_9755);
  not g20782 (n_9756, n11396);
  not g20783 (n_9757, n11397);
  and g20784 (n11398, n_9756, n_9757);
  and g20785 (n11399, \b[57] , n266);
  and g20786 (n11400, \b[55] , n284);
  and g20787 (n11401, \b[56] , n261);
  and g20793 (n11404, n_9158, n_9161);
  not g20794 (n_9762, \b[57] );
  and g20795 (n11405, n_9156, n_9762);
  and g20796 (n11406, \b[56] , \b[57] );
  not g20797 (n_9763, n11405);
  not g20798 (n_9764, n11406);
  and g20799 (n11407, n_9763, n_9764);
  not g20800 (n_9765, n11404);
  and g20801 (n11408, n_9765, n11407);
  not g20802 (n_9766, n11407);
  and g20803 (n11409, n11404, n_9766);
  not g20804 (n_9767, n11408);
  not g20805 (n_9768, n11409);
  and g20806 (n11410, n_9767, n_9768);
  and g20807 (n11411, n269, n11410);
  not g20810 (n_9770, n11412);
  and g20811 (n11413, \a[2] , n_9770);
  not g20812 (n_9771, n11413);
  and g20813 (n11414, \a[2] , n_9771);
  and g20814 (n11415, n_9770, n_9771);
  not g20815 (n_9772, n11414);
  not g20816 (n_9773, n11415);
  and g20817 (n11416, n_9772, n_9773);
  not g20818 (n_9774, n11398);
  not g20819 (n_9775, n11416);
  and g20820 (n11417, n_9774, n_9775);
  not g20821 (n_9776, n11417);
  and g20822 (n11418, n_9774, n_9776);
  and g20823 (n11419, n_9775, n_9776);
  not g20824 (n_9777, n11418);
  not g20825 (n_9778, n11419);
  and g20826 (n11420, n_9777, n_9778);
  and g20827 (n11421, n_9457, n_9462);
  not g20828 (n_9779, n11420);
  not g20829 (n_9780, n11421);
  and g20830 (n11422, n_9779, n_9780);
  and g20831 (n11423, n11420, n11421);
  not g20832 (n_9781, n11422);
  not g20833 (n_9782, n11423);
  and g20834 (\f[57] , n_9781, n_9782);
  and g20835 (n11425, \b[58] , n266);
  and g20836 (n11426, \b[56] , n284);
  and g20837 (n11427, \b[57] , n261);
  and g20843 (n11430, n_9764, n_9767);
  not g20844 (n_9787, \b[58] );
  and g20845 (n11431, n_9762, n_9787);
  and g20846 (n11432, \b[57] , \b[58] );
  not g20847 (n_9788, n11431);
  not g20848 (n_9789, n11432);
  and g20849 (n11433, n_9788, n_9789);
  not g20850 (n_9790, n11430);
  and g20851 (n11434, n_9790, n11433);
  not g20852 (n_9791, n11433);
  and g20853 (n11435, n11430, n_9791);
  not g20854 (n_9792, n11434);
  not g20855 (n_9793, n11435);
  and g20856 (n11436, n_9792, n_9793);
  and g20857 (n11437, n269, n11436);
  not g20860 (n_9795, n11438);
  and g20861 (n11439, \a[2] , n_9795);
  not g20862 (n_9796, n11439);
  and g20863 (n11440, \a[2] , n_9796);
  and g20864 (n11441, n_9795, n_9796);
  not g20865 (n_9797, n11440);
  not g20866 (n_9798, n11441);
  and g20867 (n11442, n_9797, n_9798);
  and g20868 (n11443, n_9750, n_9755);
  and g20869 (n11444, \b[55] , n362);
  and g20870 (n11445, \b[53] , n403);
  and g20871 (n11446, \b[54] , n357);
  and g20877 (n11449, n365, n10684);
  not g20880 (n_9803, n11450);
  and g20881 (n11451, \a[5] , n_9803);
  not g20882 (n_9804, n11451);
  and g20883 (n11452, \a[5] , n_9804);
  and g20884 (n11453, n_9803, n_9804);
  not g20885 (n_9805, n11452);
  not g20886 (n_9806, n11453);
  and g20887 (n11454, n_9805, n_9806);
  and g20888 (n11455, n_9742, n_9747);
  and g20889 (n11456, \b[52] , n511);
  and g20890 (n11457, \b[50] , n541);
  and g20891 (n11458, \b[51] , n506);
  and g20897 (n11461, n514, n9628);
  not g20900 (n_9811, n11462);
  and g20901 (n11463, \a[8] , n_9811);
  not g20902 (n_9812, n11463);
  and g20903 (n11464, \a[8] , n_9812);
  and g20904 (n11465, n_9811, n_9812);
  not g20905 (n_9813, n11464);
  not g20906 (n_9814, n11465);
  and g20907 (n11466, n_9813, n_9814);
  and g20908 (n11467, n_9734, n_9739);
  and g20909 (n11468, \b[49] , n700);
  and g20910 (n11469, \b[47] , n767);
  and g20911 (n11470, \b[48] , n695);
  and g20917 (n11473, n703, n8625);
  not g20920 (n_9819, n11474);
  and g20921 (n11475, \a[11] , n_9819);
  not g20922 (n_9820, n11475);
  and g20923 (n11476, \a[11] , n_9820);
  and g20924 (n11477, n_9819, n_9820);
  not g20925 (n_9821, n11476);
  not g20926 (n_9822, n11477);
  and g20927 (n11478, n_9821, n_9822);
  and g20928 (n11479, n_9726, n_9731);
  and g20929 (n11480, n_9720, n_9723);
  and g20930 (n11481, n_9655, n_9659);
  and g20931 (n11482, n_9648, n_9651);
  and g20932 (n11483, n_9606, n_9611);
  and g20933 (n11484, n_9592, n_9595);
  and g20934 (n11485, \b[10] , n8362);
  and g20935 (n11486, \b[8] , n8715);
  and g20936 (n11487, \b[9] , n8357);
  and g20942 (n11490, n738, n8365);
  not g20945 (n_9827, n11491);
  and g20946 (n11492, \a[50] , n_9827);
  not g20947 (n_9828, n11492);
  and g20948 (n11493, \a[50] , n_9828);
  and g20949 (n11494, n_9827, n_9828);
  not g20950 (n_9829, n11493);
  not g20951 (n_9830, n11494);
  and g20952 (n11495, n_9829, n_9830);
  and g20953 (n11496, n_9569, n_9570);
  not g20954 (n_9831, n11496);
  and g20955 (n11497, n_9566, n_9831);
  and g20956 (n11498, \b[7] , n9339);
  and g20957 (n11499, \b[5] , n9732);
  and g20958 (n11500, \b[6] , n9334);
  and g20964 (n11503, n484, n9342);
  not g20967 (n_9836, n11504);
  and g20968 (n11505, \a[53] , n_9836);
  not g20969 (n_9837, n11505);
  and g20970 (n11506, \a[53] , n_9837);
  and g20971 (n11507, n_9836, n_9837);
  not g20972 (n_9838, n11506);
  not g20973 (n_9839, n11507);
  and g20974 (n11508, n_9838, n_9839);
  and g20975 (n11509, n10808, n11186);
  not g20976 (n_9840, n11509);
  and g20977 (n11510, n_9563, n_9840);
  and g20978 (n11511, \b[4] , n10426);
  and g20979 (n11512, \b[2] , n10796);
  and g20980 (n11513, \b[3] , n10421);
  and g20986 (n11516, n346, n10429);
  not g20989 (n_9845, n11517);
  and g20990 (n11518, \a[56] , n_9845);
  not g20991 (n_9846, n11518);
  and g20992 (n11519, \a[56] , n_9846);
  and g20993 (n11520, n_9845, n_9846);
  not g20994 (n_9847, n11519);
  not g20995 (n_9848, n11520);
  and g20996 (n11521, n_9847, n_9848);
  and g20997 (n11522, \a[59] , n_9550);
  and g20998 (n11523, n_9546, \a[58] );
  not g20999 (n_9851, \a[58] );
  and g21000 (n11524, \a[57] , n_9851);
  not g21001 (n_9852, n11523);
  not g21002 (n_9853, n11524);
  and g21003 (n11525, n_9852, n_9853);
  not g21004 (n_9854, n11525);
  and g21005 (n11526, n11185, n_9854);
  and g21006 (n11527, \b[0] , n11526);
  and g21007 (n11528, n_9851, \a[59] );
  not g21008 (n_9855, \a[59] );
  and g21009 (n11529, \a[58] , n_9855);
  not g21010 (n_9856, n11528);
  not g21011 (n_9857, n11529);
  and g21012 (n11530, n_9856, n_9857);
  and g21013 (n11531, n_9549, n11530);
  and g21014 (n11532, \b[1] , n11531);
  not g21015 (n_9858, n11527);
  not g21016 (n_9859, n11532);
  and g21017 (n11533, n_9858, n_9859);
  not g21018 (n_9860, n11530);
  and g21019 (n11534, n_9549, n_9860);
  and g21020 (n11535, n_21, n11534);
  not g21021 (n_9861, n11535);
  and g21022 (n11536, n11533, n_9861);
  not g21023 (n_9862, n11536);
  and g21024 (n11537, \a[59] , n_9862);
  not g21025 (n_9863, n11537);
  and g21026 (n11538, \a[59] , n_9863);
  and g21027 (n11539, n_9862, n_9863);
  not g21028 (n_9864, n11538);
  not g21029 (n_9865, n11539);
  and g21030 (n11540, n_9864, n_9865);
  not g21031 (n_9866, n11540);
  and g21032 (n11541, n11522, n_9866);
  not g21033 (n_9867, n11522);
  and g21034 (n11542, n_9867, n11540);
  not g21035 (n_9868, n11541);
  not g21036 (n_9869, n11542);
  and g21037 (n11543, n_9868, n_9869);
  not g21038 (n_9870, n11543);
  and g21039 (n11544, n11521, n_9870);
  not g21040 (n_9871, n11521);
  and g21041 (n11545, n_9871, n11543);
  not g21042 (n_9872, n11544);
  not g21043 (n_9873, n11545);
  and g21044 (n11546, n_9872, n_9873);
  not g21045 (n_9874, n11510);
  and g21046 (n11547, n_9874, n11546);
  not g21047 (n_9875, n11546);
  and g21048 (n11548, n11510, n_9875);
  not g21049 (n_9876, n11547);
  not g21050 (n_9877, n11548);
  and g21051 (n11549, n_9876, n_9877);
  not g21052 (n_9878, n11549);
  and g21053 (n11550, n11508, n_9878);
  not g21054 (n_9879, n11508);
  and g21055 (n11551, n_9879, n11549);
  not g21056 (n_9880, n11550);
  not g21057 (n_9881, n11551);
  and g21058 (n11552, n_9880, n_9881);
  not g21059 (n_9882, n11497);
  and g21060 (n11553, n_9882, n11552);
  not g21061 (n_9883, n11552);
  and g21062 (n11554, n11497, n_9883);
  not g21063 (n_9884, n11553);
  not g21064 (n_9885, n11554);
  and g21065 (n11555, n_9884, n_9885);
  not g21066 (n_9886, n11495);
  and g21067 (n11556, n_9886, n11555);
  not g21068 (n_9887, n11556);
  and g21069 (n11557, n11555, n_9887);
  and g21070 (n11558, n_9886, n_9887);
  not g21071 (n_9888, n11557);
  not g21072 (n_9889, n11558);
  and g21073 (n11559, n_9888, n_9889);
  and g21074 (n11560, n_9583, n_9587);
  and g21075 (n11561, n11559, n11560);
  not g21076 (n_9890, n11559);
  not g21077 (n_9891, n11560);
  and g21078 (n11562, n_9890, n_9891);
  not g21079 (n_9892, n11561);
  not g21080 (n_9893, n11562);
  and g21081 (n11563, n_9892, n_9893);
  and g21082 (n11564, \b[13] , n7446);
  and g21083 (n11565, \b[11] , n7787);
  and g21084 (n11566, \b[12] , n7441);
  and g21090 (n11569, n1008, n7449);
  not g21093 (n_9898, n11570);
  and g21094 (n11571, \a[47] , n_9898);
  not g21095 (n_9899, n11571);
  and g21096 (n11572, \a[47] , n_9899);
  and g21097 (n11573, n_9898, n_9899);
  not g21098 (n_9900, n11572);
  not g21099 (n_9901, n11573);
  and g21100 (n11574, n_9900, n_9901);
  not g21101 (n_9902, n11574);
  and g21102 (n11575, n11563, n_9902);
  not g21103 (n_9903, n11563);
  and g21104 (n11576, n_9903, n11574);
  not g21105 (n_9904, n11484);
  not g21106 (n_9905, n11576);
  and g21107 (n11577, n_9904, n_9905);
  not g21108 (n_9906, n11575);
  and g21109 (n11578, n_9906, n11577);
  not g21110 (n_9907, n11578);
  and g21111 (n11579, n_9904, n_9907);
  and g21112 (n11580, n_9906, n_9907);
  and g21113 (n11581, n_9905, n11580);
  not g21114 (n_9908, n11579);
  not g21115 (n_9909, n11581);
  and g21116 (n11582, n_9908, n_9909);
  and g21117 (n11583, \b[16] , n6595);
  and g21118 (n11584, \b[14] , n6902);
  and g21119 (n11585, \b[15] , n6590);
  and g21125 (n11588, n1237, n6598);
  not g21128 (n_9914, n11589);
  and g21129 (n11590, \a[44] , n_9914);
  not g21130 (n_9915, n11590);
  and g21131 (n11591, \a[44] , n_9915);
  and g21132 (n11592, n_9914, n_9915);
  not g21133 (n_9916, n11591);
  not g21134 (n_9917, n11592);
  and g21135 (n11593, n_9916, n_9917);
  not g21136 (n_9918, n11582);
  not g21137 (n_9919, n11593);
  and g21138 (n11594, n_9918, n_9919);
  not g21139 (n_9920, n11594);
  and g21140 (n11595, n_9918, n_9920);
  and g21141 (n11596, n_9919, n_9920);
  not g21142 (n_9921, n11595);
  not g21143 (n_9922, n11596);
  and g21144 (n11597, n_9921, n_9922);
  and g21145 (n11598, n_9599, n_9603);
  and g21146 (n11599, n11597, n11598);
  not g21147 (n_9923, n11597);
  not g21148 (n_9924, n11598);
  and g21149 (n11600, n_9923, n_9924);
  not g21150 (n_9925, n11599);
  not g21151 (n_9926, n11600);
  and g21152 (n11601, n_9925, n_9926);
  and g21153 (n11602, \b[19] , n5777);
  and g21154 (n11603, \b[17] , n6059);
  and g21155 (n11604, \b[18] , n5772);
  and g21161 (n11607, n1708, n5780);
  not g21164 (n_9931, n11608);
  and g21165 (n11609, \a[41] , n_9931);
  not g21166 (n_9932, n11609);
  and g21167 (n11610, \a[41] , n_9932);
  and g21168 (n11611, n_9931, n_9932);
  not g21169 (n_9933, n11610);
  not g21170 (n_9934, n11611);
  and g21171 (n11612, n_9933, n_9934);
  not g21172 (n_9935, n11612);
  and g21173 (n11613, n11601, n_9935);
  not g21174 (n_9936, n11601);
  and g21175 (n11614, n_9936, n11612);
  not g21176 (n_9937, n11483);
  not g21177 (n_9938, n11614);
  and g21178 (n11615, n_9937, n_9938);
  not g21179 (n_9939, n11613);
  and g21180 (n11616, n_9939, n11615);
  not g21181 (n_9940, n11616);
  and g21182 (n11617, n_9937, n_9940);
  and g21183 (n11618, n_9939, n_9940);
  and g21184 (n11619, n_9938, n11618);
  not g21185 (n_9941, n11617);
  not g21186 (n_9942, n11619);
  and g21187 (n11620, n_9941, n_9942);
  and g21188 (n11621, \b[22] , n5035);
  and g21189 (n11622, \b[20] , n5277);
  and g21190 (n11623, \b[21] , n5030);
  and g21196 (n11626, n2145, n5038);
  not g21199 (n_9947, n11627);
  and g21200 (n11628, \a[38] , n_9947);
  not g21201 (n_9948, n11628);
  and g21202 (n11629, \a[38] , n_9948);
  and g21203 (n11630, n_9947, n_9948);
  not g21204 (n_9949, n11629);
  not g21205 (n_9950, n11630);
  and g21206 (n11631, n_9949, n_9950);
  not g21207 (n_9951, n11620);
  not g21208 (n_9952, n11631);
  and g21209 (n11632, n_9951, n_9952);
  not g21210 (n_9953, n11632);
  and g21211 (n11633, n_9951, n_9953);
  and g21212 (n11634, n_9952, n_9953);
  not g21213 (n_9954, n11633);
  not g21214 (n_9955, n11634);
  and g21215 (n11635, n_9954, n_9955);
  and g21216 (n11636, n_9615, n_9619);
  and g21217 (n11637, n11635, n11636);
  not g21218 (n_9956, n11635);
  not g21219 (n_9957, n11636);
  and g21220 (n11638, n_9956, n_9957);
  not g21221 (n_9958, n11637);
  not g21222 (n_9959, n11638);
  and g21223 (n11639, n_9958, n_9959);
  and g21224 (n11640, \b[25] , n4287);
  and g21225 (n11641, \b[23] , n4532);
  and g21226 (n11642, \b[24] , n4282);
  and g21232 (n11645, n2485, n4290);
  not g21235 (n_9964, n11646);
  and g21236 (n11647, \a[35] , n_9964);
  not g21237 (n_9965, n11647);
  and g21238 (n11648, \a[35] , n_9965);
  and g21239 (n11649, n_9964, n_9965);
  not g21240 (n_9966, n11648);
  not g21241 (n_9967, n11649);
  and g21242 (n11650, n_9966, n_9967);
  not g21243 (n_9968, n11650);
  and g21244 (n11651, n11639, n_9968);
  not g21245 (n_9969, n11651);
  and g21246 (n11652, n11639, n_9969);
  and g21247 (n11653, n_9968, n_9969);
  not g21248 (n_9970, n11652);
  not g21249 (n_9971, n11653);
  and g21250 (n11654, n_9970, n_9971);
  and g21251 (n11655, n_9630, n_9636);
  and g21252 (n11656, n11654, n11655);
  not g21253 (n_9972, n11654);
  not g21254 (n_9973, n11655);
  and g21255 (n11657, n_9972, n_9973);
  not g21256 (n_9974, n11656);
  not g21257 (n_9975, n11657);
  and g21258 (n11658, n_9974, n_9975);
  and g21259 (n11659, \b[28] , n3638);
  and g21260 (n11660, \b[26] , n3843);
  and g21261 (n11661, \b[27] , n3633);
  and g21267 (n11664, n3189, n3641);
  not g21270 (n_9980, n11665);
  and g21271 (n11666, \a[32] , n_9980);
  not g21272 (n_9981, n11666);
  and g21273 (n11667, \a[32] , n_9981);
  and g21274 (n11668, n_9980, n_9981);
  not g21275 (n_9982, n11667);
  not g21276 (n_9983, n11668);
  and g21277 (n11669, n_9982, n_9983);
  not g21278 (n_9984, n11669);
  and g21279 (n11670, n11658, n_9984);
  not g21280 (n_9985, n11670);
  and g21281 (n11671, n11658, n_9985);
  and g21282 (n11672, n_9984, n_9985);
  not g21283 (n_9986, n11671);
  not g21284 (n_9987, n11672);
  and g21285 (n11673, n_9986, n_9987);
  not g21286 (n_9988, n11482);
  and g21287 (n11674, n_9988, n11673);
  not g21288 (n_9989, n11673);
  and g21289 (n11675, n11482, n_9989);
  not g21290 (n_9990, n11674);
  not g21291 (n_9991, n11675);
  and g21292 (n11676, n_9990, n_9991);
  and g21293 (n11677, \b[31] , n3050);
  and g21294 (n11678, \b[29] , n3243);
  and g21295 (n11679, \b[30] , n3045);
  and g21301 (n11682, n3053, n3796);
  not g21304 (n_9996, n11683);
  and g21305 (n11684, \a[29] , n_9996);
  not g21306 (n_9997, n11684);
  and g21307 (n11685, \a[29] , n_9997);
  and g21308 (n11686, n_9996, n_9997);
  not g21309 (n_9998, n11685);
  not g21310 (n_9999, n11686);
  and g21311 (n11687, n_9998, n_9999);
  not g21312 (n_10000, n11676);
  not g21313 (n_10001, n11687);
  and g21314 (n11688, n_10000, n_10001);
  and g21315 (n11689, n11676, n11687);
  not g21316 (n_10002, n11688);
  not g21317 (n_10003, n11689);
  and g21318 (n11690, n_10002, n_10003);
  not g21319 (n_10004, n11690);
  and g21320 (n11691, n11481, n_10004);
  not g21321 (n_10005, n11481);
  and g21322 (n11692, n_10005, n11690);
  not g21323 (n_10006, n11691);
  not g21324 (n_10007, n11692);
  and g21325 (n11693, n_10006, n_10007);
  and g21326 (n11694, \b[34] , n2539);
  and g21327 (n11695, \b[32] , n2685);
  and g21328 (n11696, \b[33] , n2534);
  and g21334 (n11699, n2542, n4466);
  not g21337 (n_10012, n11700);
  and g21338 (n11701, \a[26] , n_10012);
  not g21339 (n_10013, n11701);
  and g21340 (n11702, \a[26] , n_10013);
  and g21341 (n11703, n_10012, n_10013);
  not g21342 (n_10014, n11702);
  not g21343 (n_10015, n11703);
  and g21344 (n11704, n_10014, n_10015);
  not g21345 (n_10016, n11704);
  and g21346 (n11705, n11693, n_10016);
  not g21347 (n_10017, n11705);
  and g21348 (n11706, n11693, n_10017);
  and g21349 (n11707, n_10016, n_10017);
  not g21350 (n_10018, n11706);
  not g21351 (n_10019, n11707);
  and g21352 (n11708, n_10018, n_10019);
  and g21353 (n11709, n_9673, n_9674);
  not g21354 (n_10020, n11709);
  and g21355 (n11710, n_9670, n_10020);
  and g21356 (n11711, n11708, n11710);
  not g21357 (n_10021, n11708);
  not g21358 (n_10022, n11710);
  and g21359 (n11712, n_10021, n_10022);
  not g21360 (n_10023, n11711);
  not g21361 (n_10024, n11712);
  and g21362 (n11713, n_10023, n_10024);
  and g21363 (n11714, \b[37] , n2048);
  and g21364 (n11715, \b[35] , n2198);
  and g21365 (n11716, \b[36] , n2043);
  and g21371 (n11719, n2051, n5181);
  not g21374 (n_10029, n11720);
  and g21375 (n11721, \a[23] , n_10029);
  not g21376 (n_10030, n11721);
  and g21377 (n11722, \a[23] , n_10030);
  and g21378 (n11723, n_10029, n_10030);
  not g21379 (n_10031, n11722);
  not g21380 (n_10032, n11723);
  and g21381 (n11724, n_10031, n_10032);
  not g21382 (n_10033, n11724);
  and g21383 (n11725, n11713, n_10033);
  not g21384 (n_10034, n11725);
  and g21385 (n11726, n11713, n_10034);
  and g21386 (n11727, n_10033, n_10034);
  not g21387 (n_10035, n11726);
  not g21388 (n_10036, n11727);
  and g21389 (n11728, n_10035, n_10036);
  and g21390 (n11729, n_9687, n_9692);
  and g21391 (n11730, n11728, n11729);
  not g21392 (n_10037, n11728);
  not g21393 (n_10038, n11729);
  and g21394 (n11731, n_10037, n_10038);
  not g21395 (n_10039, n11730);
  not g21396 (n_10040, n11731);
  and g21397 (n11732, n_10039, n_10040);
  and g21398 (n11733, \b[40] , n1627);
  and g21399 (n11734, \b[38] , n1763);
  and g21400 (n11735, \b[39] , n1622);
  and g21406 (n11738, n1630, n5955);
  not g21409 (n_10045, n11739);
  and g21410 (n11740, \a[20] , n_10045);
  not g21411 (n_10046, n11740);
  and g21412 (n11741, \a[20] , n_10046);
  and g21413 (n11742, n_10045, n_10046);
  not g21414 (n_10047, n11741);
  not g21415 (n_10048, n11742);
  and g21416 (n11743, n_10047, n_10048);
  not g21417 (n_10049, n11743);
  and g21418 (n11744, n11732, n_10049);
  not g21419 (n_10050, n11744);
  and g21420 (n11745, n11732, n_10050);
  and g21421 (n11746, n_10049, n_10050);
  not g21422 (n_10051, n11745);
  not g21423 (n_10052, n11746);
  and g21424 (n11747, n_10051, n_10052);
  and g21425 (n11748, n_9702, n_9708);
  and g21426 (n11749, n11747, n11748);
  not g21427 (n_10053, n11747);
  not g21428 (n_10054, n11748);
  and g21429 (n11750, n_10053, n_10054);
  not g21430 (n_10055, n11749);
  not g21431 (n_10056, n11750);
  and g21432 (n11751, n_10055, n_10056);
  and g21433 (n11752, \b[43] , n1302);
  and g21434 (n11753, \b[41] , n1391);
  and g21435 (n11754, \b[42] , n1297);
  and g21441 (n11757, n1305, n6515);
  not g21444 (n_10061, n11758);
  and g21445 (n11759, \a[17] , n_10061);
  not g21446 (n_10062, n11759);
  and g21447 (n11760, \a[17] , n_10062);
  and g21448 (n11761, n_10061, n_10062);
  not g21449 (n_10063, n11760);
  not g21450 (n_10064, n11761);
  and g21451 (n11762, n_10063, n_10064);
  not g21452 (n_10065, n11762);
  and g21453 (n11763, n11751, n_10065);
  not g21454 (n_10066, n11751);
  and g21455 (n11764, n_10066, n11762);
  not g21456 (n_10067, n11480);
  not g21457 (n_10068, n11764);
  and g21458 (n11765, n_10067, n_10068);
  not g21459 (n_10069, n11763);
  and g21460 (n11766, n_10069, n11765);
  not g21461 (n_10070, n11766);
  and g21462 (n11767, n_10067, n_10070);
  and g21463 (n11768, n_10069, n_10070);
  and g21464 (n11769, n_10068, n11768);
  not g21465 (n_10071, n11767);
  not g21466 (n_10072, n11769);
  and g21467 (n11770, n_10071, n_10072);
  and g21468 (n11771, \b[46] , n951);
  and g21469 (n11772, \b[44] , n1056);
  and g21470 (n11773, \b[45] , n946);
  and g21476 (n11776, n954, n7677);
  not g21479 (n_10077, n11777);
  and g21480 (n11778, \a[14] , n_10077);
  not g21481 (n_10078, n11778);
  and g21482 (n11779, \a[14] , n_10078);
  and g21483 (n11780, n_10077, n_10078);
  not g21484 (n_10079, n11779);
  not g21485 (n_10080, n11780);
  and g21486 (n11781, n_10079, n_10080);
  and g21487 (n11782, n11770, n11781);
  not g21488 (n_10081, n11770);
  not g21489 (n_10082, n11781);
  and g21490 (n11783, n_10081, n_10082);
  not g21491 (n_10083, n11782);
  not g21492 (n_10084, n11783);
  and g21493 (n11784, n_10083, n_10084);
  not g21494 (n_10085, n11479);
  and g21495 (n11785, n_10085, n11784);
  not g21496 (n_10086, n11784);
  and g21497 (n11786, n11479, n_10086);
  not g21498 (n_10087, n11785);
  not g21499 (n_10088, n11786);
  and g21500 (n11787, n_10087, n_10088);
  not g21501 (n_10089, n11787);
  and g21502 (n11788, n11478, n_10089);
  not g21503 (n_10090, n11478);
  and g21504 (n11789, n_10090, n11787);
  not g21505 (n_10091, n11788);
  not g21506 (n_10092, n11789);
  and g21507 (n11790, n_10091, n_10092);
  not g21508 (n_10093, n11467);
  and g21509 (n11791, n_10093, n11790);
  not g21510 (n_10094, n11790);
  and g21511 (n11792, n11467, n_10094);
  not g21512 (n_10095, n11791);
  not g21513 (n_10096, n11792);
  and g21514 (n11793, n_10095, n_10096);
  not g21515 (n_10097, n11793);
  and g21516 (n11794, n11466, n_10097);
  not g21517 (n_10098, n11466);
  and g21518 (n11795, n_10098, n11793);
  not g21519 (n_10099, n11794);
  not g21520 (n_10100, n11795);
  and g21521 (n11796, n_10099, n_10100);
  not g21522 (n_10101, n11455);
  and g21523 (n11797, n_10101, n11796);
  not g21524 (n_10102, n11796);
  and g21525 (n11798, n11455, n_10102);
  not g21526 (n_10103, n11797);
  not g21527 (n_10104, n11798);
  and g21528 (n11799, n_10103, n_10104);
  not g21529 (n_10105, n11799);
  and g21530 (n11800, n11454, n_10105);
  not g21531 (n_10106, n11454);
  and g21532 (n11801, n_10106, n11799);
  not g21533 (n_10107, n11800);
  not g21534 (n_10108, n11801);
  and g21535 (n11802, n_10107, n_10108);
  not g21536 (n_10109, n11443);
  and g21537 (n11803, n_10109, n11802);
  not g21538 (n_10110, n11802);
  and g21539 (n11804, n11443, n_10110);
  not g21540 (n_10111, n11803);
  not g21541 (n_10112, n11804);
  and g21542 (n11805, n_10111, n_10112);
  not g21543 (n_10113, n11442);
  and g21544 (n11806, n_10113, n11805);
  not g21545 (n_10114, n11806);
  and g21546 (n11807, n11805, n_10114);
  and g21547 (n11808, n_10113, n_10114);
  not g21548 (n_10115, n11807);
  not g21549 (n_10116, n11808);
  and g21550 (n11809, n_10115, n_10116);
  and g21551 (n11810, n_9776, n_9781);
  not g21552 (n_10117, n11809);
  not g21553 (n_10118, n11810);
  and g21554 (n11811, n_10117, n_10118);
  and g21555 (n11812, n11809, n11810);
  not g21556 (n_10119, n11811);
  not g21557 (n_10120, n11812);
  and g21558 (\f[58] , n_10119, n_10120);
  and g21559 (n11814, n_10114, n_10119);
  and g21560 (n11815, n_10108, n_10111);
  and g21561 (n11816, n_10100, n_10103);
  and g21562 (n11817, \b[53] , n511);
  and g21563 (n11818, \b[51] , n541);
  and g21564 (n11819, \b[52] , n506);
  and g21570 (n11822, n514, n9972);
  not g21573 (n_10125, n11823);
  and g21574 (n11824, \a[8] , n_10125);
  not g21575 (n_10126, n11824);
  and g21576 (n11825, \a[8] , n_10126);
  and g21577 (n11826, n_10125, n_10126);
  not g21578 (n_10127, n11825);
  not g21579 (n_10128, n11826);
  and g21580 (n11827, n_10127, n_10128);
  and g21581 (n11828, n_10092, n_10095);
  and g21582 (n11829, \b[50] , n700);
  and g21583 (n11830, \b[48] , n767);
  and g21584 (n11831, \b[49] , n695);
  and g21590 (n11834, n703, n8949);
  not g21593 (n_10133, n11835);
  and g21594 (n11836, \a[11] , n_10133);
  not g21595 (n_10134, n11836);
  and g21596 (n11837, \a[11] , n_10134);
  and g21597 (n11838, n_10133, n_10134);
  not g21598 (n_10135, n11837);
  not g21599 (n_10136, n11838);
  and g21600 (n11839, n_10135, n_10136);
  and g21601 (n11840, n_10084, n_10087);
  and g21602 (n11841, n_10050, n_10056);
  and g21603 (n11842, \b[35] , n2539);
  and g21604 (n11843, \b[33] , n2685);
  and g21605 (n11844, \b[34] , n2534);
  and g21611 (n11847, n2542, n4696);
  not g21614 (n_10141, n11848);
  and g21615 (n11849, \a[26] , n_10141);
  not g21616 (n_10142, n11849);
  and g21617 (n11850, \a[26] , n_10142);
  and g21618 (n11851, n_10141, n_10142);
  not g21619 (n_10143, n11850);
  not g21620 (n_10144, n11851);
  and g21621 (n11852, n_10143, n_10144);
  and g21622 (n11853, n_10002, n_10007);
  and g21623 (n11854, n_9988, n_9989);
  not g21624 (n_10145, n11854);
  and g21625 (n11855, n_9985, n_10145);
  and g21626 (n11856, n_9953, n_9959);
  and g21627 (n11857, n_9920, n_9926);
  and g21628 (n11858, \b[17] , n6595);
  and g21629 (n11859, \b[15] , n6902);
  and g21630 (n11860, \b[16] , n6590);
  and g21636 (n11863, n1356, n6598);
  not g21639 (n_10150, n11864);
  and g21640 (n11865, \a[44] , n_10150);
  not g21641 (n_10151, n11865);
  and g21642 (n11866, \a[44] , n_10151);
  and g21643 (n11867, n_10150, n_10151);
  not g21644 (n_10152, n11866);
  not g21645 (n_10153, n11867);
  and g21646 (n11868, n_10152, n_10153);
  and g21647 (n11869, \b[14] , n7446);
  and g21648 (n11870, \b[12] , n7787);
  and g21649 (n11871, \b[13] , n7441);
  and g21655 (n11874, n1034, n7449);
  not g21658 (n_10158, n11875);
  and g21659 (n11876, \a[47] , n_10158);
  not g21660 (n_10159, n11876);
  and g21661 (n11877, \a[47] , n_10159);
  and g21662 (n11878, n_10158, n_10159);
  not g21663 (n_10160, n11877);
  not g21664 (n_10161, n11878);
  and g21665 (n11879, n_10160, n_10161);
  and g21666 (n11880, n_9887, n_9893);
  and g21667 (n11881, \b[11] , n8362);
  and g21668 (n11882, \b[9] , n8715);
  and g21669 (n11883, \b[10] , n8357);
  and g21675 (n11886, n818, n8365);
  not g21678 (n_10166, n11887);
  and g21679 (n11888, \a[50] , n_10166);
  not g21680 (n_10167, n11888);
  and g21681 (n11889, \a[50] , n_10167);
  and g21682 (n11890, n_10166, n_10167);
  not g21683 (n_10168, n11889);
  not g21684 (n_10169, n11890);
  and g21685 (n11891, n_10168, n_10169);
  and g21686 (n11892, n_9881, n_9884);
  and g21687 (n11893, n_9873, n_9876);
  and g21688 (n11894, \b[2] , n11531);
  and g21689 (n11895, n11185, n_9860);
  and g21690 (n11896, n11525, n11895);
  and g21691 (n11897, \b[0] , n11896);
  and g21692 (n11898, \b[1] , n11526);
  and g21698 (n11901, n296, n11534);
  not g21701 (n_10174, n11902);
  and g21702 (n11903, \a[59] , n_10174);
  not g21703 (n_10175, n11903);
  and g21704 (n11904, \a[59] , n_10175);
  and g21705 (n11905, n_10174, n_10175);
  not g21706 (n_10176, n11904);
  not g21707 (n_10177, n11905);
  and g21708 (n11906, n_10176, n_10177);
  and g21709 (n11907, n_9868, n11906);
  not g21710 (n_10178, n11906);
  and g21711 (n11908, n11541, n_10178);
  not g21712 (n_10179, n11907);
  not g21713 (n_10180, n11908);
  and g21714 (n11909, n_10179, n_10180);
  and g21715 (n11910, \b[5] , n10426);
  and g21716 (n11911, \b[3] , n10796);
  and g21717 (n11912, \b[4] , n10421);
  and g21723 (n11915, n394, n10429);
  not g21726 (n_10185, n11916);
  and g21727 (n11917, \a[56] , n_10185);
  not g21728 (n_10186, n11917);
  and g21729 (n11918, \a[56] , n_10186);
  and g21730 (n11919, n_10185, n_10186);
  not g21731 (n_10187, n11918);
  not g21732 (n_10188, n11919);
  and g21733 (n11920, n_10187, n_10188);
  not g21734 (n_10189, n11920);
  and g21735 (n11921, n11909, n_10189);
  not g21736 (n_10190, n11909);
  and g21737 (n11922, n_10190, n11920);
  not g21738 (n_10191, n11893);
  not g21739 (n_10192, n11922);
  and g21740 (n11923, n_10191, n_10192);
  not g21741 (n_10193, n11921);
  and g21742 (n11924, n_10193, n11923);
  not g21743 (n_10194, n11924);
  and g21744 (n11925, n_10191, n_10194);
  and g21745 (n11926, n_10193, n_10194);
  and g21746 (n11927, n_10192, n11926);
  not g21747 (n_10195, n11925);
  not g21748 (n_10196, n11927);
  and g21749 (n11928, n_10195, n_10196);
  and g21750 (n11929, \b[8] , n9339);
  and g21751 (n11930, \b[6] , n9732);
  and g21752 (n11931, \b[7] , n9334);
  and g21758 (n11934, n585, n9342);
  not g21761 (n_10201, n11935);
  and g21762 (n11936, \a[53] , n_10201);
  not g21763 (n_10202, n11936);
  and g21764 (n11937, \a[53] , n_10202);
  and g21765 (n11938, n_10201, n_10202);
  not g21766 (n_10203, n11937);
  not g21767 (n_10204, n11938);
  and g21768 (n11939, n_10203, n_10204);
  and g21769 (n11940, n11928, n11939);
  not g21770 (n_10205, n11928);
  not g21771 (n_10206, n11939);
  and g21772 (n11941, n_10205, n_10206);
  not g21773 (n_10207, n11940);
  not g21774 (n_10208, n11941);
  and g21775 (n11942, n_10207, n_10208);
  not g21776 (n_10209, n11892);
  and g21777 (n11943, n_10209, n11942);
  not g21778 (n_10210, n11942);
  and g21779 (n11944, n11892, n_10210);
  not g21780 (n_10211, n11943);
  not g21781 (n_10212, n11944);
  and g21782 (n11945, n_10211, n_10212);
  not g21783 (n_10213, n11945);
  and g21784 (n11946, n11891, n_10213);
  not g21785 (n_10214, n11891);
  and g21786 (n11947, n_10214, n11945);
  not g21787 (n_10215, n11946);
  not g21788 (n_10216, n11947);
  and g21789 (n11948, n_10215, n_10216);
  not g21790 (n_10217, n11880);
  and g21791 (n11949, n_10217, n11948);
  not g21792 (n_10218, n11948);
  and g21793 (n11950, n11880, n_10218);
  not g21794 (n_10219, n11949);
  not g21795 (n_10220, n11950);
  and g21796 (n11951, n_10219, n_10220);
  not g21797 (n_10221, n11879);
  and g21798 (n11952, n_10221, n11951);
  not g21799 (n_10222, n11952);
  and g21800 (n11953, n11951, n_10222);
  and g21801 (n11954, n_10221, n_10222);
  not g21802 (n_10223, n11953);
  not g21803 (n_10224, n11954);
  and g21804 (n11955, n_10223, n_10224);
  not g21805 (n_10225, n11580);
  not g21806 (n_10226, n11955);
  and g21807 (n11956, n_10225, n_10226);
  and g21808 (n11957, n11580, n11955);
  not g21809 (n_10227, n11956);
  not g21810 (n_10228, n11957);
  and g21811 (n11958, n_10227, n_10228);
  not g21812 (n_10229, n11868);
  and g21813 (n11959, n_10229, n11958);
  not g21814 (n_10230, n11959);
  and g21815 (n11960, n_10229, n_10230);
  and g21816 (n11961, n11958, n_10230);
  not g21817 (n_10231, n11960);
  not g21818 (n_10232, n11961);
  and g21819 (n11962, n_10231, n_10232);
  not g21820 (n_10233, n11857);
  not g21821 (n_10234, n11962);
  and g21822 (n11963, n_10233, n_10234);
  not g21823 (n_10235, n11963);
  and g21824 (n11964, n_10233, n_10235);
  and g21825 (n11965, n_10234, n_10235);
  not g21826 (n_10236, n11964);
  not g21827 (n_10237, n11965);
  and g21828 (n11966, n_10236, n_10237);
  and g21829 (n11967, \b[20] , n5777);
  and g21830 (n11968, \b[18] , n6059);
  and g21831 (n11969, \b[19] , n5772);
  and g21837 (n11972, n1846, n5780);
  not g21840 (n_10242, n11973);
  and g21841 (n11974, \a[41] , n_10242);
  not g21842 (n_10243, n11974);
  and g21843 (n11975, \a[41] , n_10243);
  and g21844 (n11976, n_10242, n_10243);
  not g21845 (n_10244, n11975);
  not g21846 (n_10245, n11976);
  and g21847 (n11977, n_10244, n_10245);
  not g21848 (n_10246, n11966);
  not g21849 (n_10247, n11977);
  and g21850 (n11978, n_10246, n_10247);
  not g21851 (n_10248, n11978);
  and g21852 (n11979, n_10246, n_10248);
  and g21853 (n11980, n_10247, n_10248);
  not g21854 (n_10249, n11979);
  not g21855 (n_10250, n11980);
  and g21856 (n11981, n_10249, n_10250);
  not g21857 (n_10251, n11618);
  and g21858 (n11982, n_10251, n11981);
  not g21859 (n_10252, n11981);
  and g21860 (n11983, n11618, n_10252);
  not g21861 (n_10253, n11982);
  not g21862 (n_10254, n11983);
  and g21863 (n11984, n_10253, n_10254);
  and g21864 (n11985, \b[23] , n5035);
  and g21865 (n11986, \b[21] , n5277);
  and g21866 (n11987, \b[22] , n5030);
  and g21872 (n11990, n2300, n5038);
  not g21875 (n_10259, n11991);
  and g21876 (n11992, \a[38] , n_10259);
  not g21877 (n_10260, n11992);
  and g21878 (n11993, \a[38] , n_10260);
  and g21879 (n11994, n_10259, n_10260);
  not g21880 (n_10261, n11993);
  not g21881 (n_10262, n11994);
  and g21882 (n11995, n_10261, n_10262);
  not g21883 (n_10263, n11984);
  not g21884 (n_10264, n11995);
  and g21885 (n11996, n_10263, n_10264);
  and g21886 (n11997, n11984, n11995);
  not g21887 (n_10265, n11996);
  not g21888 (n_10266, n11997);
  and g21889 (n11998, n_10265, n_10266);
  not g21890 (n_10267, n11998);
  and g21891 (n11999, n11856, n_10267);
  not g21892 (n_10268, n11856);
  and g21893 (n12000, n_10268, n11998);
  not g21894 (n_10269, n11999);
  not g21895 (n_10270, n12000);
  and g21896 (n12001, n_10269, n_10270);
  and g21897 (n12002, \b[26] , n4287);
  and g21898 (n12003, \b[24] , n4532);
  and g21899 (n12004, \b[25] , n4282);
  and g21905 (n12007, n2813, n4290);
  not g21908 (n_10275, n12008);
  and g21909 (n12009, \a[35] , n_10275);
  not g21910 (n_10276, n12009);
  and g21911 (n12010, \a[35] , n_10276);
  and g21912 (n12011, n_10275, n_10276);
  not g21913 (n_10277, n12010);
  not g21914 (n_10278, n12011);
  and g21915 (n12012, n_10277, n_10278);
  not g21916 (n_10279, n12012);
  and g21917 (n12013, n12001, n_10279);
  not g21918 (n_10280, n12013);
  and g21919 (n12014, n12001, n_10280);
  and g21920 (n12015, n_10279, n_10280);
  not g21921 (n_10281, n12014);
  not g21922 (n_10282, n12015);
  and g21923 (n12016, n_10281, n_10282);
  and g21924 (n12017, n_9969, n_9975);
  and g21925 (n12018, n12016, n12017);
  not g21926 (n_10283, n12016);
  not g21927 (n_10284, n12017);
  and g21928 (n12019, n_10283, n_10284);
  not g21929 (n_10285, n12018);
  not g21930 (n_10286, n12019);
  and g21931 (n12020, n_10285, n_10286);
  and g21932 (n12021, \b[29] , n3638);
  and g21933 (n12022, \b[27] , n3843);
  and g21934 (n12023, \b[28] , n3633);
  and g21940 (n12026, n3383, n3641);
  not g21943 (n_10291, n12027);
  and g21944 (n12028, \a[32] , n_10291);
  not g21945 (n_10292, n12028);
  and g21946 (n12029, \a[32] , n_10292);
  and g21947 (n12030, n_10291, n_10292);
  not g21948 (n_10293, n12029);
  not g21949 (n_10294, n12030);
  and g21950 (n12031, n_10293, n_10294);
  not g21951 (n_10295, n12031);
  and g21952 (n12032, n12020, n_10295);
  not g21953 (n_10296, n12020);
  and g21954 (n12033, n_10296, n12031);
  not g21955 (n_10297, n11855);
  not g21956 (n_10298, n12033);
  and g21957 (n12034, n_10297, n_10298);
  not g21958 (n_10299, n12032);
  and g21959 (n12035, n_10299, n12034);
  not g21960 (n_10300, n12035);
  and g21961 (n12036, n_10297, n_10300);
  and g21962 (n12037, n_10299, n_10300);
  and g21963 (n12038, n_10298, n12037);
  not g21964 (n_10301, n12036);
  not g21965 (n_10302, n12038);
  and g21966 (n12039, n_10301, n_10302);
  and g21967 (n12040, \b[32] , n3050);
  and g21968 (n12041, \b[30] , n3243);
  and g21969 (n12042, \b[31] , n3045);
  and g21975 (n12045, n3053, n4013);
  not g21978 (n_10307, n12046);
  and g21979 (n12047, \a[29] , n_10307);
  not g21980 (n_10308, n12047);
  and g21981 (n12048, \a[29] , n_10308);
  and g21982 (n12049, n_10307, n_10308);
  not g21983 (n_10309, n12048);
  not g21984 (n_10310, n12049);
  and g21985 (n12050, n_10309, n_10310);
  and g21986 (n12051, n12039, n12050);
  not g21987 (n_10311, n12039);
  not g21988 (n_10312, n12050);
  and g21989 (n12052, n_10311, n_10312);
  not g21990 (n_10313, n12051);
  not g21991 (n_10314, n12052);
  and g21992 (n12053, n_10313, n_10314);
  not g21993 (n_10315, n11853);
  and g21994 (n12054, n_10315, n12053);
  not g21995 (n_10316, n12053);
  and g21996 (n12055, n11853, n_10316);
  not g21997 (n_10317, n12054);
  not g21998 (n_10318, n12055);
  and g21999 (n12056, n_10317, n_10318);
  not g22000 (n_10319, n11852);
  and g22001 (n12057, n_10319, n12056);
  not g22002 (n_10320, n12057);
  and g22003 (n12058, n12056, n_10320);
  and g22004 (n12059, n_10319, n_10320);
  not g22005 (n_10321, n12058);
  not g22006 (n_10322, n12059);
  and g22007 (n12060, n_10321, n_10322);
  and g22008 (n12061, n_10017, n_10024);
  and g22009 (n12062, n12060, n12061);
  not g22010 (n_10323, n12060);
  not g22011 (n_10324, n12061);
  and g22012 (n12063, n_10323, n_10324);
  not g22013 (n_10325, n12062);
  not g22014 (n_10326, n12063);
  and g22015 (n12064, n_10325, n_10326);
  and g22016 (n12065, \b[38] , n2048);
  and g22017 (n12066, \b[36] , n2198);
  and g22018 (n12067, \b[37] , n2043);
  and g22024 (n12070, n2051, n5205);
  not g22027 (n_10331, n12071);
  and g22028 (n12072, \a[23] , n_10331);
  not g22029 (n_10332, n12072);
  and g22030 (n12073, \a[23] , n_10332);
  and g22031 (n12074, n_10331, n_10332);
  not g22032 (n_10333, n12073);
  not g22033 (n_10334, n12074);
  and g22034 (n12075, n_10333, n_10334);
  not g22035 (n_10335, n12075);
  and g22036 (n12076, n12064, n_10335);
  not g22037 (n_10336, n12076);
  and g22038 (n12077, n12064, n_10336);
  and g22039 (n12078, n_10335, n_10336);
  not g22040 (n_10337, n12077);
  not g22041 (n_10338, n12078);
  and g22042 (n12079, n_10337, n_10338);
  and g22043 (n12080, n_10034, n_10040);
  and g22044 (n12081, n12079, n12080);
  not g22045 (n_10339, n12079);
  not g22046 (n_10340, n12080);
  and g22047 (n12082, n_10339, n_10340);
  not g22048 (n_10341, n12081);
  not g22049 (n_10342, n12082);
  and g22050 (n12083, n_10341, n_10342);
  and g22051 (n12084, \b[41] , n1627);
  and g22052 (n12085, \b[39] , n1763);
  and g22053 (n12086, \b[40] , n1622);
  and g22059 (n12089, n1630, n6219);
  not g22062 (n_10347, n12090);
  and g22063 (n12091, \a[20] , n_10347);
  not g22064 (n_10348, n12091);
  and g22065 (n12092, \a[20] , n_10348);
  and g22066 (n12093, n_10347, n_10348);
  not g22067 (n_10349, n12092);
  not g22068 (n_10350, n12093);
  and g22069 (n12094, n_10349, n_10350);
  not g22070 (n_10351, n12094);
  and g22071 (n12095, n12083, n_10351);
  not g22072 (n_10352, n12083);
  and g22073 (n12096, n_10352, n12094);
  not g22074 (n_10353, n11841);
  not g22075 (n_10354, n12096);
  and g22076 (n12097, n_10353, n_10354);
  not g22077 (n_10355, n12095);
  and g22078 (n12098, n_10355, n12097);
  not g22079 (n_10356, n12098);
  and g22080 (n12099, n_10353, n_10356);
  and g22081 (n12100, n_10355, n_10356);
  and g22082 (n12101, n_10354, n12100);
  not g22083 (n_10357, n12099);
  not g22084 (n_10358, n12101);
  and g22085 (n12102, n_10357, n_10358);
  and g22086 (n12103, \b[44] , n1302);
  and g22087 (n12104, \b[42] , n1391);
  and g22088 (n12105, \b[43] , n1297);
  and g22094 (n12108, n1305, n7072);
  not g22097 (n_10363, n12109);
  and g22098 (n12110, \a[17] , n_10363);
  not g22099 (n_10364, n12110);
  and g22100 (n12111, \a[17] , n_10364);
  and g22101 (n12112, n_10363, n_10364);
  not g22102 (n_10365, n12111);
  not g22103 (n_10366, n12112);
  and g22104 (n12113, n_10365, n_10366);
  not g22105 (n_10367, n12102);
  not g22106 (n_10368, n12113);
  and g22107 (n12114, n_10367, n_10368);
  not g22108 (n_10369, n12114);
  and g22109 (n12115, n_10367, n_10369);
  and g22110 (n12116, n_10368, n_10369);
  not g22111 (n_10370, n12115);
  not g22112 (n_10371, n12116);
  and g22113 (n12117, n_10370, n_10371);
  not g22114 (n_10372, n11768);
  and g22115 (n12118, n_10372, n12117);
  not g22116 (n_10373, n12117);
  and g22117 (n12119, n11768, n_10373);
  not g22118 (n_10374, n12118);
  not g22119 (n_10375, n12119);
  and g22120 (n12120, n_10374, n_10375);
  and g22121 (n12121, \b[47] , n951);
  and g22122 (n12122, \b[45] , n1056);
  and g22123 (n12123, \b[46] , n946);
  and g22129 (n12126, n954, n7703);
  not g22132 (n_10380, n12127);
  and g22133 (n12128, \a[14] , n_10380);
  not g22134 (n_10381, n12128);
  and g22135 (n12129, \a[14] , n_10381);
  and g22136 (n12130, n_10380, n_10381);
  not g22137 (n_10382, n12129);
  not g22138 (n_10383, n12130);
  and g22139 (n12131, n_10382, n_10383);
  not g22140 (n_10384, n12120);
  not g22141 (n_10385, n12131);
  and g22142 (n12132, n_10384, n_10385);
  and g22143 (n12133, n12120, n12131);
  not g22144 (n_10386, n12132);
  not g22145 (n_10387, n12133);
  and g22146 (n12134, n_10386, n_10387);
  not g22147 (n_10388, n11840);
  and g22148 (n12135, n_10388, n12134);
  not g22149 (n_10389, n12134);
  and g22150 (n12136, n11840, n_10389);
  not g22151 (n_10390, n12135);
  not g22152 (n_10391, n12136);
  and g22153 (n12137, n_10390, n_10391);
  not g22154 (n_10392, n11839);
  and g22155 (n12138, n_10392, n12137);
  not g22156 (n_10393, n12138);
  and g22157 (n12139, n12137, n_10393);
  and g22158 (n12140, n_10392, n_10393);
  not g22159 (n_10394, n12139);
  not g22160 (n_10395, n12140);
  and g22161 (n12141, n_10394, n_10395);
  not g22162 (n_10396, n11828);
  not g22163 (n_10397, n12141);
  and g22164 (n12142, n_10396, n_10397);
  and g22165 (n12143, n11828, n12141);
  not g22166 (n_10398, n12142);
  not g22167 (n_10399, n12143);
  and g22168 (n12144, n_10398, n_10399);
  not g22169 (n_10400, n11827);
  and g22170 (n12145, n_10400, n12144);
  not g22171 (n_10401, n12145);
  and g22172 (n12146, n_10400, n_10401);
  and g22173 (n12147, n12144, n_10401);
  not g22174 (n_10402, n12146);
  not g22175 (n_10403, n12147);
  and g22176 (n12148, n_10402, n_10403);
  not g22177 (n_10404, n11816);
  not g22178 (n_10405, n12148);
  and g22179 (n12149, n_10404, n_10405);
  not g22180 (n_10406, n12149);
  and g22181 (n12150, n_10404, n_10406);
  and g22182 (n12151, n_10405, n_10406);
  not g22183 (n_10407, n12150);
  not g22184 (n_10408, n12151);
  and g22185 (n12152, n_10407, n_10408);
  and g22186 (n12153, \b[56] , n362);
  and g22187 (n12154, \b[54] , n403);
  and g22188 (n12155, \b[55] , n357);
  and g22194 (n12158, n365, n10708);
  not g22197 (n_10413, n12159);
  and g22198 (n12160, \a[5] , n_10413);
  not g22199 (n_10414, n12160);
  and g22200 (n12161, \a[5] , n_10414);
  and g22201 (n12162, n_10413, n_10414);
  not g22202 (n_10415, n12161);
  not g22203 (n_10416, n12162);
  and g22204 (n12163, n_10415, n_10416);
  not g22205 (n_10417, n12152);
  not g22206 (n_10418, n12163);
  and g22207 (n12164, n_10417, n_10418);
  not g22208 (n_10419, n12164);
  and g22209 (n12165, n_10417, n_10419);
  and g22210 (n12166, n_10418, n_10419);
  not g22211 (n_10420, n12165);
  not g22212 (n_10421, n12166);
  and g22213 (n12167, n_10420, n_10421);
  and g22214 (n12168, \b[59] , n266);
  and g22215 (n12169, \b[57] , n284);
  and g22216 (n12170, \b[58] , n261);
  and g22222 (n12173, n_9789, n_9792);
  not g22223 (n_10426, \b[59] );
  and g22224 (n12174, n_9787, n_10426);
  and g22225 (n12175, \b[58] , \b[59] );
  not g22226 (n_10427, n12174);
  not g22227 (n_10428, n12175);
  and g22228 (n12176, n_10427, n_10428);
  not g22229 (n_10429, n12173);
  and g22230 (n12177, n_10429, n12176);
  not g22231 (n_10430, n12176);
  and g22232 (n12178, n12173, n_10430);
  not g22233 (n_10431, n12177);
  not g22234 (n_10432, n12178);
  and g22235 (n12179, n_10431, n_10432);
  and g22236 (n12180, n269, n12179);
  not g22239 (n_10434, n12181);
  and g22240 (n12182, \a[2] , n_10434);
  not g22241 (n_10435, n12182);
  and g22242 (n12183, \a[2] , n_10435);
  and g22243 (n12184, n_10434, n_10435);
  not g22244 (n_10436, n12183);
  not g22245 (n_10437, n12184);
  and g22246 (n12185, n_10436, n_10437);
  not g22247 (n_10438, n12167);
  and g22248 (n12186, n_10438, n12185);
  not g22249 (n_10439, n12185);
  and g22250 (n12187, n12167, n_10439);
  not g22251 (n_10440, n12186);
  not g22252 (n_10441, n12187);
  and g22253 (n12188, n_10440, n_10441);
  not g22254 (n_10442, n11815);
  not g22255 (n_10443, n12188);
  and g22256 (n12189, n_10442, n_10443);
  not g22257 (n_10444, n12189);
  and g22258 (n12190, n_10442, n_10444);
  and g22259 (n12191, n_10443, n_10444);
  not g22260 (n_10445, n12190);
  not g22261 (n_10446, n12191);
  and g22262 (n12192, n_10445, n_10446);
  not g22263 (n_10447, n11814);
  not g22264 (n_10448, n12192);
  and g22265 (n12193, n_10447, n_10448);
  and g22266 (n12194, n11814, n_10446);
  and g22267 (n12195, n_10445, n12194);
  not g22268 (n_10449, n12193);
  not g22269 (n_10450, n12195);
  and g22270 (\f[59] , n_10449, n_10450);
  and g22271 (n12197, n_10444, n_10449);
  and g22272 (n12198, n_10438, n_10439);
  not g22273 (n_10451, n12198);
  and g22274 (n12199, n_10419, n_10451);
  and g22275 (n12200, \b[60] , n266);
  and g22276 (n12201, \b[58] , n284);
  and g22277 (n12202, \b[59] , n261);
  and g22283 (n12205, n_10428, n_10431);
  not g22284 (n_10456, \b[60] );
  and g22285 (n12206, n_10426, n_10456);
  and g22286 (n12207, \b[59] , \b[60] );
  not g22287 (n_10457, n12206);
  not g22288 (n_10458, n12207);
  and g22289 (n12208, n_10457, n_10458);
  not g22290 (n_10459, n12205);
  and g22291 (n12209, n_10459, n12208);
  not g22292 (n_10460, n12208);
  and g22293 (n12210, n12205, n_10460);
  not g22294 (n_10461, n12209);
  not g22295 (n_10462, n12210);
  and g22296 (n12211, n_10461, n_10462);
  and g22297 (n12212, n269, n12211);
  not g22300 (n_10464, n12213);
  and g22301 (n12214, \a[2] , n_10464);
  not g22302 (n_10465, n12214);
  and g22303 (n12215, \a[2] , n_10465);
  and g22304 (n12216, n_10464, n_10465);
  not g22305 (n_10466, n12215);
  not g22306 (n_10467, n12216);
  and g22307 (n12217, n_10466, n_10467);
  and g22308 (n12218, \b[57] , n362);
  and g22309 (n12219, \b[55] , n403);
  and g22310 (n12220, \b[56] , n357);
  and g22316 (n12223, n365, n11410);
  not g22319 (n_10472, n12224);
  and g22320 (n12225, \a[5] , n_10472);
  not g22321 (n_10473, n12225);
  and g22322 (n12226, \a[5] , n_10473);
  and g22323 (n12227, n_10472, n_10473);
  not g22324 (n_10474, n12226);
  not g22325 (n_10475, n12227);
  and g22326 (n12228, n_10474, n_10475);
  and g22327 (n12229, n_10401, n_10406);
  and g22328 (n12230, \b[54] , n511);
  and g22329 (n12231, \b[52] , n541);
  and g22330 (n12232, \b[53] , n506);
  and g22336 (n12235, n514, n9998);
  not g22339 (n_10480, n12236);
  and g22340 (n12237, \a[8] , n_10480);
  not g22341 (n_10481, n12237);
  and g22342 (n12238, \a[8] , n_10481);
  and g22343 (n12239, n_10480, n_10481);
  not g22344 (n_10482, n12238);
  not g22345 (n_10483, n12239);
  and g22346 (n12240, n_10482, n_10483);
  and g22347 (n12241, n_10393, n_10398);
  and g22348 (n12242, \b[51] , n700);
  and g22349 (n12243, \b[49] , n767);
  and g22350 (n12244, \b[50] , n695);
  and g22356 (n12247, n703, n8976);
  not g22359 (n_10488, n12248);
  and g22360 (n12249, \a[11] , n_10488);
  not g22361 (n_10489, n12249);
  and g22362 (n12250, \a[11] , n_10489);
  and g22363 (n12251, n_10488, n_10489);
  not g22364 (n_10490, n12250);
  not g22365 (n_10491, n12251);
  and g22366 (n12252, n_10490, n_10491);
  and g22367 (n12253, n_10386, n_10390);
  and g22368 (n12254, \b[48] , n951);
  and g22369 (n12255, \b[46] , n1056);
  and g22370 (n12256, \b[47] , n946);
  and g22376 (n12259, n954, n8009);
  not g22379 (n_10496, n12260);
  and g22380 (n12261, \a[14] , n_10496);
  not g22381 (n_10497, n12261);
  and g22382 (n12262, \a[14] , n_10497);
  and g22383 (n12263, n_10496, n_10497);
  not g22384 (n_10498, n12262);
  not g22385 (n_10499, n12263);
  and g22386 (n12264, n_10498, n_10499);
  and g22387 (n12265, n_10372, n_10373);
  not g22388 (n_10500, n12265);
  and g22389 (n12266, n_10369, n_10500);
  and g22390 (n12267, \b[45] , n1302);
  and g22391 (n12268, \b[43] , n1391);
  and g22392 (n12269, \b[44] , n1297);
  and g22398 (n12272, n1305, n7361);
  not g22401 (n_10505, n12273);
  and g22402 (n12274, \a[17] , n_10505);
  not g22403 (n_10506, n12274);
  and g22404 (n12275, \a[17] , n_10506);
  and g22405 (n12276, n_10505, n_10506);
  not g22406 (n_10507, n12275);
  not g22407 (n_10508, n12276);
  and g22408 (n12277, n_10507, n_10508);
  and g22409 (n12278, n_10320, n_10326);
  and g22410 (n12279, n_10314, n_10317);
  and g22411 (n12280, \b[33] , n3050);
  and g22412 (n12281, \b[31] , n3243);
  and g22413 (n12282, \b[32] , n3045);
  and g22419 (n12285, n3053, n4223);
  not g22422 (n_10513, n12286);
  and g22423 (n12287, \a[29] , n_10513);
  not g22424 (n_10514, n12287);
  and g22425 (n12288, \a[29] , n_10514);
  and g22426 (n12289, n_10513, n_10514);
  not g22427 (n_10515, n12288);
  not g22428 (n_10516, n12289);
  and g22429 (n12290, n_10515, n_10516);
  and g22430 (n12291, n_10251, n_10252);
  not g22431 (n_10517, n12291);
  and g22432 (n12292, n_10248, n_10517);
  and g22433 (n12293, \b[21] , n5777);
  and g22434 (n12294, \b[19] , n6059);
  and g22435 (n12295, \b[20] , n5772);
  and g22441 (n12298, n1984, n5780);
  not g22444 (n_10522, n12299);
  and g22445 (n12300, \a[41] , n_10522);
  not g22446 (n_10523, n12300);
  and g22447 (n12301, \a[41] , n_10523);
  and g22448 (n12302, n_10522, n_10523);
  not g22449 (n_10524, n12301);
  not g22450 (n_10525, n12302);
  and g22451 (n12303, n_10524, n_10525);
  and g22452 (n12304, n_10230, n_10235);
  and g22453 (n12305, \b[18] , n6595);
  and g22454 (n12306, \b[16] , n6902);
  and g22455 (n12307, \b[17] , n6590);
  and g22461 (n12310, n1566, n6598);
  not g22464 (n_10530, n12311);
  and g22465 (n12312, \a[44] , n_10530);
  not g22466 (n_10531, n12312);
  and g22467 (n12313, \a[44] , n_10531);
  and g22468 (n12314, n_10530, n_10531);
  not g22469 (n_10532, n12313);
  not g22470 (n_10533, n12314);
  and g22471 (n12315, n_10532, n_10533);
  and g22472 (n12316, n_10222, n_10227);
  and g22473 (n12317, \b[15] , n7446);
  and g22474 (n12318, \b[13] , n7787);
  and g22475 (n12319, \b[14] , n7441);
  and g22481 (n12322, n1131, n7449);
  not g22484 (n_10538, n12323);
  and g22485 (n12324, \a[47] , n_10538);
  not g22486 (n_10539, n12324);
  and g22487 (n12325, \a[47] , n_10539);
  and g22488 (n12326, n_10538, n_10539);
  not g22489 (n_10540, n12325);
  not g22490 (n_10541, n12326);
  and g22491 (n12327, n_10540, n_10541);
  and g22492 (n12328, n_10216, n_10219);
  and g22493 (n12329, \b[12] , n8362);
  and g22494 (n12330, \b[10] , n8715);
  and g22495 (n12331, \b[11] , n8357);
  and g22501 (n12334, n842, n8365);
  not g22504 (n_10546, n12335);
  and g22505 (n12336, \a[50] , n_10546);
  not g22506 (n_10547, n12336);
  and g22507 (n12337, \a[50] , n_10547);
  and g22508 (n12338, n_10546, n_10547);
  not g22509 (n_10548, n12337);
  not g22510 (n_10549, n12338);
  and g22511 (n12339, n_10548, n_10549);
  and g22512 (n12340, n_10208, n_10211);
  and g22513 (n12341, \b[6] , n10426);
  and g22514 (n12342, \b[4] , n10796);
  and g22515 (n12343, \b[5] , n10421);
  and g22521 (n12346, n459, n10429);
  not g22524 (n_10554, n12347);
  and g22525 (n12348, \a[56] , n_10554);
  not g22526 (n_10555, n12348);
  and g22527 (n12349, \a[56] , n_10555);
  and g22528 (n12350, n_10554, n_10555);
  not g22529 (n_10556, n12349);
  not g22530 (n_10557, n12350);
  and g22531 (n12351, n_10556, n_10557);
  not g22532 (n_10559, \a[60] );
  and g22533 (n12352, \a[59] , n_10559);
  and g22534 (n12353, n_9855, \a[60] );
  not g22535 (n_10560, n12352);
  not g22536 (n_10561, n12353);
  and g22537 (n12354, n_10560, n_10561);
  not g22538 (n_10562, n12354);
  and g22539 (n12355, \b[0] , n_10562);
  and g22540 (n12356, n_10180, n12355);
  not g22541 (n_10563, n12355);
  and g22542 (n12357, n11908, n_10563);
  not g22543 (n_10564, n12356);
  not g22544 (n_10565, n12357);
  and g22545 (n12358, n_10564, n_10565);
  and g22546 (n12359, \b[3] , n11531);
  and g22547 (n12360, \b[1] , n11896);
  and g22548 (n12361, \b[2] , n11526);
  and g22554 (n12364, n318, n11534);
  not g22557 (n_10570, n12365);
  and g22558 (n12366, \a[59] , n_10570);
  not g22559 (n_10571, n12366);
  and g22560 (n12367, \a[59] , n_10571);
  and g22561 (n12368, n_10570, n_10571);
  not g22562 (n_10572, n12367);
  not g22563 (n_10573, n12368);
  and g22564 (n12369, n_10572, n_10573);
  not g22565 (n_10574, n12358);
  not g22566 (n_10575, n12369);
  and g22567 (n12370, n_10574, n_10575);
  and g22568 (n12371, n12358, n12369);
  not g22569 (n_10576, n12370);
  not g22570 (n_10577, n12371);
  and g22571 (n12372, n_10576, n_10577);
  not g22572 (n_10578, n12351);
  and g22573 (n12373, n_10578, n12372);
  not g22574 (n_10579, n12373);
  and g22575 (n12374, n12372, n_10579);
  and g22576 (n12375, n_10578, n_10579);
  not g22577 (n_10580, n12374);
  not g22578 (n_10581, n12375);
  and g22579 (n12376, n_10580, n_10581);
  not g22580 (n_10582, n11926);
  and g22581 (n12377, n_10582, n12376);
  not g22582 (n_10583, n12376);
  and g22583 (n12378, n11926, n_10583);
  not g22584 (n_10584, n12377);
  not g22585 (n_10585, n12378);
  and g22586 (n12379, n_10584, n_10585);
  and g22587 (n12380, \b[9] , n9339);
  and g22588 (n12381, \b[7] , n9732);
  and g22589 (n12382, \b[8] , n9334);
  and g22595 (n12385, n651, n9342);
  not g22598 (n_10590, n12386);
  and g22599 (n12387, \a[53] , n_10590);
  not g22600 (n_10591, n12387);
  and g22601 (n12388, \a[53] , n_10591);
  and g22602 (n12389, n_10590, n_10591);
  not g22603 (n_10592, n12388);
  not g22604 (n_10593, n12389);
  and g22605 (n12390, n_10592, n_10593);
  not g22606 (n_10594, n12379);
  not g22607 (n_10595, n12390);
  and g22608 (n12391, n_10594, n_10595);
  and g22609 (n12392, n12379, n12390);
  not g22610 (n_10596, n12391);
  not g22611 (n_10597, n12392);
  and g22612 (n12393, n_10596, n_10597);
  not g22613 (n_10598, n12340);
  and g22614 (n12394, n_10598, n12393);
  not g22615 (n_10599, n12393);
  and g22616 (n12395, n12340, n_10599);
  not g22617 (n_10600, n12394);
  not g22618 (n_10601, n12395);
  and g22619 (n12396, n_10600, n_10601);
  not g22620 (n_10602, n12396);
  and g22621 (n12397, n12339, n_10602);
  not g22622 (n_10603, n12339);
  and g22623 (n12398, n_10603, n12396);
  not g22624 (n_10604, n12397);
  not g22625 (n_10605, n12398);
  and g22626 (n12399, n_10604, n_10605);
  not g22627 (n_10606, n12328);
  and g22628 (n12400, n_10606, n12399);
  not g22629 (n_10607, n12399);
  and g22630 (n12401, n12328, n_10607);
  not g22631 (n_10608, n12400);
  not g22632 (n_10609, n12401);
  and g22633 (n12402, n_10608, n_10609);
  not g22634 (n_10610, n12327);
  and g22635 (n12403, n_10610, n12402);
  not g22636 (n_10611, n12402);
  and g22637 (n12404, n12327, n_10611);
  not g22638 (n_10612, n12403);
  not g22639 (n_10613, n12404);
  and g22640 (n12405, n_10612, n_10613);
  not g22641 (n_10614, n12316);
  and g22642 (n12406, n_10614, n12405);
  not g22643 (n_10615, n12405);
  and g22644 (n12407, n12316, n_10615);
  not g22645 (n_10616, n12406);
  not g22646 (n_10617, n12407);
  and g22647 (n12408, n_10616, n_10617);
  not g22648 (n_10618, n12315);
  and g22649 (n12409, n_10618, n12408);
  not g22650 (n_10619, n12409);
  and g22651 (n12410, n_10618, n_10619);
  and g22652 (n12411, n12408, n_10619);
  not g22653 (n_10620, n12410);
  not g22654 (n_10621, n12411);
  and g22655 (n12412, n_10620, n_10621);
  not g22656 (n_10622, n12304);
  not g22657 (n_10623, n12412);
  and g22658 (n12413, n_10622, n_10623);
  and g22659 (n12414, n12304, n_10621);
  and g22660 (n12415, n_10620, n12414);
  not g22661 (n_10624, n12413);
  not g22662 (n_10625, n12415);
  and g22663 (n12416, n_10624, n_10625);
  not g22664 (n_10626, n12303);
  and g22665 (n12417, n_10626, n12416);
  not g22666 (n_10627, n12416);
  and g22667 (n12418, n12303, n_10627);
  not g22668 (n_10628, n12417);
  not g22669 (n_10629, n12418);
  and g22670 (n12419, n_10628, n_10629);
  not g22671 (n_10630, n12292);
  and g22672 (n12420, n_10630, n12419);
  not g22673 (n_10631, n12419);
  and g22674 (n12421, n12292, n_10631);
  not g22675 (n_10632, n12420);
  not g22676 (n_10633, n12421);
  and g22677 (n12422, n_10632, n_10633);
  and g22678 (n12423, \b[24] , n5035);
  and g22679 (n12424, \b[22] , n5277);
  and g22680 (n12425, \b[23] , n5030);
  and g22686 (n12428, n2458, n5038);
  not g22689 (n_10638, n12429);
  and g22690 (n12430, \a[38] , n_10638);
  not g22691 (n_10639, n12430);
  and g22692 (n12431, \a[38] , n_10639);
  and g22693 (n12432, n_10638, n_10639);
  not g22694 (n_10640, n12431);
  not g22695 (n_10641, n12432);
  and g22696 (n12433, n_10640, n_10641);
  not g22697 (n_10642, n12433);
  and g22698 (n12434, n12422, n_10642);
  not g22699 (n_10643, n12434);
  and g22700 (n12435, n12422, n_10643);
  and g22701 (n12436, n_10642, n_10643);
  not g22702 (n_10644, n12435);
  not g22703 (n_10645, n12436);
  and g22704 (n12437, n_10644, n_10645);
  and g22705 (n12438, n_10265, n_10270);
  and g22706 (n12439, n12437, n12438);
  not g22707 (n_10646, n12437);
  not g22708 (n_10647, n12438);
  and g22709 (n12440, n_10646, n_10647);
  not g22710 (n_10648, n12439);
  not g22711 (n_10649, n12440);
  and g22712 (n12441, n_10648, n_10649);
  and g22713 (n12442, \b[27] , n4287);
  and g22714 (n12443, \b[25] , n4532);
  and g22715 (n12444, \b[26] , n4282);
  and g22721 (n12447, n2990, n4290);
  not g22724 (n_10654, n12448);
  and g22725 (n12449, \a[35] , n_10654);
  not g22726 (n_10655, n12449);
  and g22727 (n12450, \a[35] , n_10655);
  and g22728 (n12451, n_10654, n_10655);
  not g22729 (n_10656, n12450);
  not g22730 (n_10657, n12451);
  and g22731 (n12452, n_10656, n_10657);
  not g22732 (n_10658, n12452);
  and g22733 (n12453, n12441, n_10658);
  not g22734 (n_10659, n12453);
  and g22735 (n12454, n12441, n_10659);
  and g22736 (n12455, n_10658, n_10659);
  not g22737 (n_10660, n12454);
  not g22738 (n_10661, n12455);
  and g22739 (n12456, n_10660, n_10661);
  and g22740 (n12457, n_10280, n_10286);
  and g22741 (n12458, n12456, n12457);
  not g22742 (n_10662, n12456);
  not g22743 (n_10663, n12457);
  and g22744 (n12459, n_10662, n_10663);
  not g22745 (n_10664, n12458);
  not g22746 (n_10665, n12459);
  and g22747 (n12460, n_10664, n_10665);
  and g22748 (n12461, \b[30] , n3638);
  and g22749 (n12462, \b[28] , n3843);
  and g22750 (n12463, \b[29] , n3633);
  and g22756 (n12466, n3577, n3641);
  not g22759 (n_10670, n12467);
  and g22760 (n12468, \a[32] , n_10670);
  not g22761 (n_10671, n12468);
  and g22762 (n12469, \a[32] , n_10671);
  and g22763 (n12470, n_10670, n_10671);
  not g22764 (n_10672, n12469);
  not g22765 (n_10673, n12470);
  and g22766 (n12471, n_10672, n_10673);
  not g22767 (n_10674, n12460);
  and g22768 (n12472, n_10674, n12471);
  not g22769 (n_10675, n12471);
  and g22770 (n12473, n12460, n_10675);
  not g22771 (n_10676, n12472);
  not g22772 (n_10677, n12473);
  and g22773 (n12474, n_10676, n_10677);
  not g22774 (n_10678, n12037);
  and g22775 (n12475, n_10678, n12474);
  not g22776 (n_10679, n12474);
  and g22777 (n12476, n12037, n_10679);
  not g22778 (n_10680, n12475);
  not g22779 (n_10681, n12476);
  and g22780 (n12477, n_10680, n_10681);
  not g22781 (n_10682, n12290);
  and g22782 (n12478, n_10682, n12477);
  not g22783 (n_10683, n12478);
  and g22784 (n12479, n12477, n_10683);
  and g22785 (n12480, n_10682, n_10683);
  not g22786 (n_10684, n12479);
  not g22787 (n_10685, n12480);
  and g22788 (n12481, n_10684, n_10685);
  not g22789 (n_10686, n12279);
  and g22790 (n12482, n_10686, n12481);
  not g22791 (n_10687, n12481);
  and g22792 (n12483, n12279, n_10687);
  not g22793 (n_10688, n12482);
  not g22794 (n_10689, n12483);
  and g22795 (n12484, n_10688, n_10689);
  and g22796 (n12485, \b[36] , n2539);
  and g22797 (n12486, \b[34] , n2685);
  and g22798 (n12487, \b[35] , n2534);
  and g22804 (n12490, n2542, n4922);
  not g22807 (n_10694, n12491);
  and g22808 (n12492, \a[26] , n_10694);
  not g22809 (n_10695, n12492);
  and g22810 (n12493, \a[26] , n_10695);
  and g22811 (n12494, n_10694, n_10695);
  not g22812 (n_10696, n12493);
  not g22813 (n_10697, n12494);
  and g22814 (n12495, n_10696, n_10697);
  not g22815 (n_10698, n12484);
  not g22816 (n_10699, n12495);
  and g22817 (n12496, n_10698, n_10699);
  and g22818 (n12497, n12484, n12495);
  not g22819 (n_10700, n12496);
  not g22820 (n_10701, n12497);
  and g22821 (n12498, n_10700, n_10701);
  not g22822 (n_10702, n12498);
  and g22823 (n12499, n12278, n_10702);
  not g22824 (n_10703, n12278);
  and g22825 (n12500, n_10703, n12498);
  not g22826 (n_10704, n12499);
  not g22827 (n_10705, n12500);
  and g22828 (n12501, n_10704, n_10705);
  and g22829 (n12502, \b[39] , n2048);
  and g22830 (n12503, \b[37] , n2198);
  and g22831 (n12504, \b[38] , n2043);
  and g22837 (n12507, n2051, n5451);
  not g22840 (n_10710, n12508);
  and g22841 (n12509, \a[23] , n_10710);
  not g22842 (n_10711, n12509);
  and g22843 (n12510, \a[23] , n_10711);
  and g22844 (n12511, n_10710, n_10711);
  not g22845 (n_10712, n12510);
  not g22846 (n_10713, n12511);
  and g22847 (n12512, n_10712, n_10713);
  not g22848 (n_10714, n12512);
  and g22849 (n12513, n12501, n_10714);
  not g22850 (n_10715, n12513);
  and g22851 (n12514, n12501, n_10715);
  and g22852 (n12515, n_10714, n_10715);
  not g22853 (n_10716, n12514);
  not g22854 (n_10717, n12515);
  and g22855 (n12516, n_10716, n_10717);
  and g22856 (n12517, n_10336, n_10342);
  and g22857 (n12518, n12516, n12517);
  not g22858 (n_10718, n12516);
  not g22859 (n_10719, n12517);
  and g22860 (n12519, n_10718, n_10719);
  not g22861 (n_10720, n12518);
  not g22862 (n_10721, n12519);
  and g22863 (n12520, n_10720, n_10721);
  and g22864 (n12521, \b[42] , n1627);
  and g22865 (n12522, \b[40] , n1763);
  and g22866 (n12523, \b[41] , n1622);
  and g22872 (n12526, n1630, n6489);
  not g22875 (n_10726, n12527);
  and g22876 (n12528, \a[20] , n_10726);
  not g22877 (n_10727, n12528);
  and g22878 (n12529, \a[20] , n_10727);
  and g22879 (n12530, n_10726, n_10727);
  not g22880 (n_10728, n12529);
  not g22881 (n_10729, n12530);
  and g22882 (n12531, n_10728, n_10729);
  not g22883 (n_10730, n12520);
  and g22884 (n12532, n_10730, n12531);
  not g22885 (n_10731, n12531);
  and g22886 (n12533, n12520, n_10731);
  not g22887 (n_10732, n12532);
  not g22888 (n_10733, n12533);
  and g22889 (n12534, n_10732, n_10733);
  not g22890 (n_10734, n12100);
  and g22891 (n12535, n_10734, n12534);
  not g22892 (n_10735, n12534);
  and g22893 (n12536, n12100, n_10735);
  not g22894 (n_10736, n12535);
  not g22895 (n_10737, n12536);
  and g22896 (n12537, n_10736, n_10737);
  not g22897 (n_10738, n12277);
  and g22898 (n12538, n_10738, n12537);
  not g22899 (n_10739, n12538);
  and g22900 (n12539, n_10738, n_10739);
  and g22901 (n12540, n12537, n_10739);
  not g22902 (n_10740, n12539);
  not g22903 (n_10741, n12540);
  and g22904 (n12541, n_10740, n_10741);
  not g22905 (n_10742, n12266);
  not g22906 (n_10743, n12541);
  and g22907 (n12542, n_10742, n_10743);
  and g22908 (n12543, n12266, n_10741);
  and g22909 (n12544, n_10740, n12543);
  not g22910 (n_10744, n12542);
  not g22911 (n_10745, n12544);
  and g22912 (n12545, n_10744, n_10745);
  not g22913 (n_10746, n12264);
  and g22914 (n12546, n_10746, n12545);
  not g22915 (n_10747, n12546);
  and g22916 (n12547, n_10746, n_10747);
  and g22917 (n12548, n12545, n_10747);
  not g22918 (n_10748, n12547);
  not g22919 (n_10749, n12548);
  and g22920 (n12549, n_10748, n_10749);
  not g22921 (n_10750, n12253);
  not g22922 (n_10751, n12549);
  and g22923 (n12550, n_10750, n_10751);
  and g22924 (n12551, n12253, n_10749);
  and g22925 (n12552, n_10748, n12551);
  not g22926 (n_10752, n12550);
  not g22927 (n_10753, n12552);
  and g22928 (n12553, n_10752, n_10753);
  not g22929 (n_10754, n12252);
  and g22930 (n12554, n_10754, n12553);
  not g22931 (n_10755, n12554);
  and g22932 (n12555, n_10754, n_10755);
  and g22933 (n12556, n12553, n_10755);
  not g22934 (n_10756, n12555);
  not g22935 (n_10757, n12556);
  and g22936 (n12557, n_10756, n_10757);
  not g22937 (n_10758, n12241);
  not g22938 (n_10759, n12557);
  and g22939 (n12558, n_10758, n_10759);
  and g22940 (n12559, n12241, n_10757);
  and g22941 (n12560, n_10756, n12559);
  not g22942 (n_10760, n12558);
  not g22943 (n_10761, n12560);
  and g22944 (n12561, n_10760, n_10761);
  not g22945 (n_10762, n12240);
  and g22946 (n12562, n_10762, n12561);
  not g22947 (n_10763, n12561);
  and g22948 (n12563, n12240, n_10763);
  not g22949 (n_10764, n12562);
  not g22950 (n_10765, n12563);
  and g22951 (n12564, n_10764, n_10765);
  not g22952 (n_10766, n12229);
  and g22953 (n12565, n_10766, n12564);
  not g22954 (n_10767, n12564);
  and g22955 (n12566, n12229, n_10767);
  not g22956 (n_10768, n12565);
  not g22957 (n_10769, n12566);
  and g22958 (n12567, n_10768, n_10769);
  not g22959 (n_10770, n12228);
  and g22960 (n12568, n_10770, n12567);
  not g22961 (n_10771, n12567);
  and g22962 (n12569, n12228, n_10771);
  not g22963 (n_10772, n12568);
  not g22964 (n_10773, n12569);
  and g22965 (n12570, n_10772, n_10773);
  not g22966 (n_10774, n12217);
  and g22967 (n12571, n_10774, n12570);
  not g22968 (n_10775, n12570);
  and g22969 (n12572, n12217, n_10775);
  not g22970 (n_10776, n12571);
  not g22971 (n_10777, n12572);
  and g22972 (n12573, n_10776, n_10777);
  not g22973 (n_10778, n12199);
  and g22974 (n12574, n_10778, n12573);
  not g22975 (n_10779, n12573);
  and g22976 (n12575, n12199, n_10779);
  not g22977 (n_10780, n12574);
  not g22978 (n_10781, n12575);
  and g22979 (n12576, n_10780, n_10781);
  not g22980 (n_10782, n12197);
  and g22981 (n12577, n_10782, n12576);
  not g22982 (n_10783, n12576);
  and g22983 (n12578, n12197, n_10783);
  not g22984 (n_10784, n12577);
  not g22985 (n_10785, n12578);
  and g22986 (\f[60] , n_10784, n_10785);
  and g22987 (n12580, \b[55] , n511);
  and g22988 (n12581, \b[53] , n541);
  and g22989 (n12582, \b[54] , n506);
  and g22995 (n12585, n514, n10684);
  not g22998 (n_10790, n12586);
  and g22999 (n12587, \a[8] , n_10790);
  not g23000 (n_10791, n12587);
  and g23001 (n12588, \a[8] , n_10791);
  and g23002 (n12589, n_10790, n_10791);
  not g23003 (n_10792, n12588);
  not g23004 (n_10793, n12589);
  and g23005 (n12590, n_10792, n_10793);
  and g23006 (n12591, n_10755, n_10760);
  and g23007 (n12592, \b[52] , n700);
  and g23008 (n12593, \b[50] , n767);
  and g23009 (n12594, \b[51] , n695);
  and g23015 (n12597, n703, n9628);
  not g23018 (n_10798, n12598);
  and g23019 (n12599, \a[11] , n_10798);
  not g23020 (n_10799, n12599);
  and g23021 (n12600, \a[11] , n_10799);
  and g23022 (n12601, n_10798, n_10799);
  not g23023 (n_10800, n12600);
  not g23024 (n_10801, n12601);
  and g23025 (n12602, n_10800, n_10801);
  and g23026 (n12603, n_10747, n_10752);
  and g23027 (n12604, \b[49] , n951);
  and g23028 (n12605, \b[47] , n1056);
  and g23029 (n12606, \b[48] , n946);
  and g23035 (n12609, n954, n8625);
  not g23038 (n_10806, n12610);
  and g23039 (n12611, \a[14] , n_10806);
  not g23040 (n_10807, n12611);
  and g23041 (n12612, \a[14] , n_10807);
  and g23042 (n12613, n_10806, n_10807);
  not g23043 (n_10808, n12612);
  not g23044 (n_10809, n12613);
  and g23045 (n12614, n_10808, n_10809);
  and g23046 (n12615, n_10739, n_10744);
  and g23047 (n12616, n_10733, n_10736);
  and g23048 (n12617, n_10686, n_10687);
  not g23049 (n_10810, n12617);
  and g23050 (n12618, n_10683, n_10810);
  and g23051 (n12619, n_10677, n_10680);
  and g23052 (n12620, n_10619, n_10624);
  and g23053 (n12621, n_10605, n_10608);
  and g23054 (n12622, \b[10] , n9339);
  and g23055 (n12623, \b[8] , n9732);
  and g23056 (n12624, \b[9] , n9334);
  and g23062 (n12627, n738, n9342);
  not g23065 (n_10815, n12628);
  and g23066 (n12629, \a[53] , n_10815);
  not g23067 (n_10816, n12629);
  and g23068 (n12630, \a[53] , n_10816);
  and g23069 (n12631, n_10815, n_10816);
  not g23070 (n_10817, n12630);
  not g23071 (n_10818, n12631);
  and g23072 (n12632, n_10817, n_10818);
  and g23073 (n12633, n_10582, n_10583);
  not g23074 (n_10819, n12633);
  and g23075 (n12634, n_10579, n_10819);
  and g23076 (n12635, \b[7] , n10426);
  and g23077 (n12636, \b[5] , n10796);
  and g23078 (n12637, \b[6] , n10421);
  and g23084 (n12640, n484, n10429);
  not g23087 (n_10824, n12641);
  and g23088 (n12642, \a[56] , n_10824);
  not g23089 (n_10825, n12642);
  and g23090 (n12643, \a[56] , n_10825);
  and g23091 (n12644, n_10824, n_10825);
  not g23092 (n_10826, n12643);
  not g23093 (n_10827, n12644);
  and g23094 (n12645, n_10826, n_10827);
  and g23095 (n12646, n11908, n12355);
  not g23096 (n_10828, n12646);
  and g23097 (n12647, n_10576, n_10828);
  and g23098 (n12648, \b[4] , n11531);
  and g23099 (n12649, \b[2] , n11896);
  and g23100 (n12650, \b[3] , n11526);
  and g23106 (n12653, n346, n11534);
  not g23109 (n_10833, n12654);
  and g23110 (n12655, \a[59] , n_10833);
  not g23111 (n_10834, n12655);
  and g23112 (n12656, \a[59] , n_10834);
  and g23113 (n12657, n_10833, n_10834);
  not g23114 (n_10835, n12656);
  not g23115 (n_10836, n12657);
  and g23116 (n12658, n_10835, n_10836);
  and g23117 (n12659, \a[62] , n_10563);
  and g23118 (n12660, n_10559, \a[61] );
  not g23119 (n_10839, \a[61] );
  and g23120 (n12661, \a[60] , n_10839);
  not g23121 (n_10840, n12660);
  not g23122 (n_10841, n12661);
  and g23123 (n12662, n_10840, n_10841);
  not g23124 (n_10842, n12662);
  and g23125 (n12663, n12354, n_10842);
  and g23126 (n12664, \b[0] , n12663);
  and g23127 (n12665, n_10839, \a[62] );
  not g23128 (n_10843, \a[62] );
  and g23129 (n12666, \a[61] , n_10843);
  not g23130 (n_10844, n12665);
  not g23131 (n_10845, n12666);
  and g23132 (n12667, n_10844, n_10845);
  and g23133 (n12668, n_10562, n12667);
  and g23134 (n12669, \b[1] , n12668);
  not g23135 (n_10846, n12664);
  not g23136 (n_10847, n12669);
  and g23137 (n12670, n_10846, n_10847);
  not g23138 (n_10848, n12667);
  and g23139 (n12671, n_10562, n_10848);
  and g23140 (n12672, n_21, n12671);
  not g23141 (n_10849, n12672);
  and g23142 (n12673, n12670, n_10849);
  not g23143 (n_10850, n12673);
  and g23144 (n12674, \a[62] , n_10850);
  not g23145 (n_10851, n12674);
  and g23146 (n12675, \a[62] , n_10851);
  and g23147 (n12676, n_10850, n_10851);
  not g23148 (n_10852, n12675);
  not g23149 (n_10853, n12676);
  and g23150 (n12677, n_10852, n_10853);
  not g23151 (n_10854, n12677);
  and g23152 (n12678, n12659, n_10854);
  not g23153 (n_10855, n12659);
  and g23154 (n12679, n_10855, n12677);
  not g23155 (n_10856, n12678);
  not g23156 (n_10857, n12679);
  and g23157 (n12680, n_10856, n_10857);
  not g23158 (n_10858, n12680);
  and g23159 (n12681, n12658, n_10858);
  not g23160 (n_10859, n12658);
  and g23161 (n12682, n_10859, n12680);
  not g23162 (n_10860, n12681);
  not g23163 (n_10861, n12682);
  and g23164 (n12683, n_10860, n_10861);
  not g23165 (n_10862, n12647);
  and g23166 (n12684, n_10862, n12683);
  not g23167 (n_10863, n12683);
  and g23168 (n12685, n12647, n_10863);
  not g23169 (n_10864, n12684);
  not g23170 (n_10865, n12685);
  and g23171 (n12686, n_10864, n_10865);
  not g23172 (n_10866, n12686);
  and g23173 (n12687, n12645, n_10866);
  not g23174 (n_10867, n12645);
  and g23175 (n12688, n_10867, n12686);
  not g23176 (n_10868, n12687);
  not g23177 (n_10869, n12688);
  and g23178 (n12689, n_10868, n_10869);
  not g23179 (n_10870, n12634);
  and g23180 (n12690, n_10870, n12689);
  not g23181 (n_10871, n12689);
  and g23182 (n12691, n12634, n_10871);
  not g23183 (n_10872, n12690);
  not g23184 (n_10873, n12691);
  and g23185 (n12692, n_10872, n_10873);
  not g23186 (n_10874, n12632);
  and g23187 (n12693, n_10874, n12692);
  not g23188 (n_10875, n12693);
  and g23189 (n12694, n12692, n_10875);
  and g23190 (n12695, n_10874, n_10875);
  not g23191 (n_10876, n12694);
  not g23192 (n_10877, n12695);
  and g23193 (n12696, n_10876, n_10877);
  and g23194 (n12697, n_10596, n_10600);
  and g23195 (n12698, n12696, n12697);
  not g23196 (n_10878, n12696);
  not g23197 (n_10879, n12697);
  and g23198 (n12699, n_10878, n_10879);
  not g23199 (n_10880, n12698);
  not g23200 (n_10881, n12699);
  and g23201 (n12700, n_10880, n_10881);
  and g23202 (n12701, \b[13] , n8362);
  and g23203 (n12702, \b[11] , n8715);
  and g23204 (n12703, \b[12] , n8357);
  and g23210 (n12706, n1008, n8365);
  not g23213 (n_10886, n12707);
  and g23214 (n12708, \a[50] , n_10886);
  not g23215 (n_10887, n12708);
  and g23216 (n12709, \a[50] , n_10887);
  and g23217 (n12710, n_10886, n_10887);
  not g23218 (n_10888, n12709);
  not g23219 (n_10889, n12710);
  and g23220 (n12711, n_10888, n_10889);
  not g23221 (n_10890, n12711);
  and g23222 (n12712, n12700, n_10890);
  not g23223 (n_10891, n12700);
  and g23224 (n12713, n_10891, n12711);
  not g23225 (n_10892, n12621);
  not g23226 (n_10893, n12713);
  and g23227 (n12714, n_10892, n_10893);
  not g23228 (n_10894, n12712);
  and g23229 (n12715, n_10894, n12714);
  not g23230 (n_10895, n12715);
  and g23231 (n12716, n_10892, n_10895);
  and g23232 (n12717, n_10894, n_10895);
  and g23233 (n12718, n_10893, n12717);
  not g23234 (n_10896, n12716);
  not g23235 (n_10897, n12718);
  and g23236 (n12719, n_10896, n_10897);
  and g23237 (n12720, \b[16] , n7446);
  and g23238 (n12721, \b[14] , n7787);
  and g23239 (n12722, \b[15] , n7441);
  and g23245 (n12725, n1237, n7449);
  not g23248 (n_10902, n12726);
  and g23249 (n12727, \a[47] , n_10902);
  not g23250 (n_10903, n12727);
  and g23251 (n12728, \a[47] , n_10903);
  and g23252 (n12729, n_10902, n_10903);
  not g23253 (n_10904, n12728);
  not g23254 (n_10905, n12729);
  and g23255 (n12730, n_10904, n_10905);
  not g23256 (n_10906, n12719);
  not g23257 (n_10907, n12730);
  and g23258 (n12731, n_10906, n_10907);
  not g23259 (n_10908, n12731);
  and g23260 (n12732, n_10906, n_10908);
  and g23261 (n12733, n_10907, n_10908);
  not g23262 (n_10909, n12732);
  not g23263 (n_10910, n12733);
  and g23264 (n12734, n_10909, n_10910);
  and g23265 (n12735, n_10612, n_10616);
  and g23266 (n12736, n12734, n12735);
  not g23267 (n_10911, n12734);
  not g23268 (n_10912, n12735);
  and g23269 (n12737, n_10911, n_10912);
  not g23270 (n_10913, n12736);
  not g23271 (n_10914, n12737);
  and g23272 (n12738, n_10913, n_10914);
  and g23273 (n12739, \b[19] , n6595);
  and g23274 (n12740, \b[17] , n6902);
  and g23275 (n12741, \b[18] , n6590);
  and g23281 (n12744, n1708, n6598);
  not g23284 (n_10919, n12745);
  and g23285 (n12746, \a[44] , n_10919);
  not g23286 (n_10920, n12746);
  and g23287 (n12747, \a[44] , n_10920);
  and g23288 (n12748, n_10919, n_10920);
  not g23289 (n_10921, n12747);
  not g23290 (n_10922, n12748);
  and g23291 (n12749, n_10921, n_10922);
  not g23292 (n_10923, n12749);
  and g23293 (n12750, n12738, n_10923);
  not g23294 (n_10924, n12738);
  and g23295 (n12751, n_10924, n12749);
  not g23296 (n_10925, n12620);
  not g23297 (n_10926, n12751);
  and g23298 (n12752, n_10925, n_10926);
  not g23299 (n_10927, n12750);
  and g23300 (n12753, n_10927, n12752);
  not g23301 (n_10928, n12753);
  and g23302 (n12754, n_10925, n_10928);
  and g23303 (n12755, n_10927, n_10928);
  and g23304 (n12756, n_10926, n12755);
  not g23305 (n_10929, n12754);
  not g23306 (n_10930, n12756);
  and g23307 (n12757, n_10929, n_10930);
  and g23308 (n12758, \b[22] , n5777);
  and g23309 (n12759, \b[20] , n6059);
  and g23310 (n12760, \b[21] , n5772);
  and g23316 (n12763, n2145, n5780);
  not g23319 (n_10935, n12764);
  and g23320 (n12765, \a[41] , n_10935);
  not g23321 (n_10936, n12765);
  and g23322 (n12766, \a[41] , n_10936);
  and g23323 (n12767, n_10935, n_10936);
  not g23324 (n_10937, n12766);
  not g23325 (n_10938, n12767);
  and g23326 (n12768, n_10937, n_10938);
  not g23327 (n_10939, n12757);
  not g23328 (n_10940, n12768);
  and g23329 (n12769, n_10939, n_10940);
  not g23330 (n_10941, n12769);
  and g23331 (n12770, n_10939, n_10941);
  and g23332 (n12771, n_10940, n_10941);
  not g23333 (n_10942, n12770);
  not g23334 (n_10943, n12771);
  and g23335 (n12772, n_10942, n_10943);
  and g23336 (n12773, n_10628, n_10632);
  and g23337 (n12774, n12772, n12773);
  not g23338 (n_10944, n12772);
  not g23339 (n_10945, n12773);
  and g23340 (n12775, n_10944, n_10945);
  not g23341 (n_10946, n12774);
  not g23342 (n_10947, n12775);
  and g23343 (n12776, n_10946, n_10947);
  and g23344 (n12777, \b[25] , n5035);
  and g23345 (n12778, \b[23] , n5277);
  and g23346 (n12779, \b[24] , n5030);
  and g23352 (n12782, n2485, n5038);
  not g23355 (n_10952, n12783);
  and g23356 (n12784, \a[38] , n_10952);
  not g23357 (n_10953, n12784);
  and g23358 (n12785, \a[38] , n_10953);
  and g23359 (n12786, n_10952, n_10953);
  not g23360 (n_10954, n12785);
  not g23361 (n_10955, n12786);
  and g23362 (n12787, n_10954, n_10955);
  not g23363 (n_10956, n12787);
  and g23364 (n12788, n12776, n_10956);
  not g23365 (n_10957, n12788);
  and g23366 (n12789, n12776, n_10957);
  and g23367 (n12790, n_10956, n_10957);
  not g23368 (n_10958, n12789);
  not g23369 (n_10959, n12790);
  and g23370 (n12791, n_10958, n_10959);
  and g23371 (n12792, n_10643, n_10649);
  and g23372 (n12793, n12791, n12792);
  not g23373 (n_10960, n12791);
  not g23374 (n_10961, n12792);
  and g23375 (n12794, n_10960, n_10961);
  not g23376 (n_10962, n12793);
  not g23377 (n_10963, n12794);
  and g23378 (n12795, n_10962, n_10963);
  and g23379 (n12796, \b[28] , n4287);
  and g23380 (n12797, \b[26] , n4532);
  and g23381 (n12798, \b[27] , n4282);
  and g23387 (n12801, n3189, n4290);
  not g23390 (n_10968, n12802);
  and g23391 (n12803, \a[35] , n_10968);
  not g23392 (n_10969, n12803);
  and g23393 (n12804, \a[35] , n_10969);
  and g23394 (n12805, n_10968, n_10969);
  not g23395 (n_10970, n12804);
  not g23396 (n_10971, n12805);
  and g23397 (n12806, n_10970, n_10971);
  not g23398 (n_10972, n12806);
  and g23399 (n12807, n12795, n_10972);
  not g23400 (n_10973, n12807);
  and g23401 (n12808, n12795, n_10973);
  and g23402 (n12809, n_10972, n_10973);
  not g23403 (n_10974, n12808);
  not g23404 (n_10975, n12809);
  and g23405 (n12810, n_10974, n_10975);
  and g23406 (n12811, n_10659, n_10665);
  and g23407 (n12812, n12810, n12811);
  not g23408 (n_10976, n12810);
  not g23409 (n_10977, n12811);
  and g23410 (n12813, n_10976, n_10977);
  not g23411 (n_10978, n12812);
  not g23412 (n_10979, n12813);
  and g23413 (n12814, n_10978, n_10979);
  and g23414 (n12815, \b[31] , n3638);
  and g23415 (n12816, \b[29] , n3843);
  and g23416 (n12817, \b[30] , n3633);
  and g23422 (n12820, n3641, n3796);
  not g23425 (n_10984, n12821);
  and g23426 (n12822, \a[32] , n_10984);
  not g23427 (n_10985, n12822);
  and g23428 (n12823, \a[32] , n_10985);
  and g23429 (n12824, n_10984, n_10985);
  not g23430 (n_10986, n12823);
  not g23431 (n_10987, n12824);
  and g23432 (n12825, n_10986, n_10987);
  not g23433 (n_10988, n12825);
  and g23434 (n12826, n12814, n_10988);
  not g23435 (n_10989, n12826);
  and g23436 (n12827, n12814, n_10989);
  and g23437 (n12828, n_10988, n_10989);
  not g23438 (n_10990, n12827);
  not g23439 (n_10991, n12828);
  and g23440 (n12829, n_10990, n_10991);
  not g23441 (n_10992, n12619);
  and g23442 (n12830, n_10992, n12829);
  not g23443 (n_10993, n12829);
  and g23444 (n12831, n12619, n_10993);
  not g23445 (n_10994, n12830);
  not g23446 (n_10995, n12831);
  and g23447 (n12832, n_10994, n_10995);
  and g23448 (n12833, \b[34] , n3050);
  and g23449 (n12834, \b[32] , n3243);
  and g23450 (n12835, \b[33] , n3045);
  and g23456 (n12838, n3053, n4466);
  not g23459 (n_11000, n12839);
  and g23460 (n12840, \a[29] , n_11000);
  not g23461 (n_11001, n12840);
  and g23462 (n12841, \a[29] , n_11001);
  and g23463 (n12842, n_11000, n_11001);
  not g23464 (n_11002, n12841);
  not g23465 (n_11003, n12842);
  and g23466 (n12843, n_11002, n_11003);
  not g23467 (n_11004, n12832);
  not g23468 (n_11005, n12843);
  and g23469 (n12844, n_11004, n_11005);
  and g23470 (n12845, n12832, n12843);
  not g23471 (n_11006, n12844);
  not g23472 (n_11007, n12845);
  and g23473 (n12846, n_11006, n_11007);
  not g23474 (n_11008, n12846);
  and g23475 (n12847, n12618, n_11008);
  not g23476 (n_11009, n12618);
  and g23477 (n12848, n_11009, n12846);
  not g23478 (n_11010, n12847);
  not g23479 (n_11011, n12848);
  and g23480 (n12849, n_11010, n_11011);
  and g23481 (n12850, \b[37] , n2539);
  and g23482 (n12851, \b[35] , n2685);
  and g23483 (n12852, \b[36] , n2534);
  and g23489 (n12855, n2542, n5181);
  not g23492 (n_11016, n12856);
  and g23493 (n12857, \a[26] , n_11016);
  not g23494 (n_11017, n12857);
  and g23495 (n12858, \a[26] , n_11017);
  and g23496 (n12859, n_11016, n_11017);
  not g23497 (n_11018, n12858);
  not g23498 (n_11019, n12859);
  and g23499 (n12860, n_11018, n_11019);
  not g23500 (n_11020, n12860);
  and g23501 (n12861, n12849, n_11020);
  not g23502 (n_11021, n12861);
  and g23503 (n12862, n12849, n_11021);
  and g23504 (n12863, n_11020, n_11021);
  not g23505 (n_11022, n12862);
  not g23506 (n_11023, n12863);
  and g23507 (n12864, n_11022, n_11023);
  and g23508 (n12865, n_10700, n_10705);
  and g23509 (n12866, n12864, n12865);
  not g23510 (n_11024, n12864);
  not g23511 (n_11025, n12865);
  and g23512 (n12867, n_11024, n_11025);
  not g23513 (n_11026, n12866);
  not g23514 (n_11027, n12867);
  and g23515 (n12868, n_11026, n_11027);
  and g23516 (n12869, \b[40] , n2048);
  and g23517 (n12870, \b[38] , n2198);
  and g23518 (n12871, \b[39] , n2043);
  and g23524 (n12874, n2051, n5955);
  not g23527 (n_11032, n12875);
  and g23528 (n12876, \a[23] , n_11032);
  not g23529 (n_11033, n12876);
  and g23530 (n12877, \a[23] , n_11033);
  and g23531 (n12878, n_11032, n_11033);
  not g23532 (n_11034, n12877);
  not g23533 (n_11035, n12878);
  and g23534 (n12879, n_11034, n_11035);
  not g23535 (n_11036, n12879);
  and g23536 (n12880, n12868, n_11036);
  not g23537 (n_11037, n12880);
  and g23538 (n12881, n12868, n_11037);
  and g23539 (n12882, n_11036, n_11037);
  not g23540 (n_11038, n12881);
  not g23541 (n_11039, n12882);
  and g23542 (n12883, n_11038, n_11039);
  and g23543 (n12884, n_10715, n_10721);
  and g23544 (n12885, n12883, n12884);
  not g23545 (n_11040, n12883);
  not g23546 (n_11041, n12884);
  and g23547 (n12886, n_11040, n_11041);
  not g23548 (n_11042, n12885);
  not g23549 (n_11043, n12886);
  and g23550 (n12887, n_11042, n_11043);
  and g23551 (n12888, \b[43] , n1627);
  and g23552 (n12889, \b[41] , n1763);
  and g23553 (n12890, \b[42] , n1622);
  and g23559 (n12893, n1630, n6515);
  not g23562 (n_11048, n12894);
  and g23563 (n12895, \a[20] , n_11048);
  not g23564 (n_11049, n12895);
  and g23565 (n12896, \a[20] , n_11049);
  and g23566 (n12897, n_11048, n_11049);
  not g23567 (n_11050, n12896);
  not g23568 (n_11051, n12897);
  and g23569 (n12898, n_11050, n_11051);
  not g23570 (n_11052, n12898);
  and g23571 (n12899, n12887, n_11052);
  not g23572 (n_11053, n12887);
  and g23573 (n12900, n_11053, n12898);
  not g23574 (n_11054, n12616);
  not g23575 (n_11055, n12900);
  and g23576 (n12901, n_11054, n_11055);
  not g23577 (n_11056, n12899);
  and g23578 (n12902, n_11056, n12901);
  not g23579 (n_11057, n12902);
  and g23580 (n12903, n_11054, n_11057);
  and g23581 (n12904, n_11056, n_11057);
  and g23582 (n12905, n_11055, n12904);
  not g23583 (n_11058, n12903);
  not g23584 (n_11059, n12905);
  and g23585 (n12906, n_11058, n_11059);
  and g23586 (n12907, \b[46] , n1302);
  and g23587 (n12908, \b[44] , n1391);
  and g23588 (n12909, \b[45] , n1297);
  and g23594 (n12912, n1305, n7677);
  not g23597 (n_11064, n12913);
  and g23598 (n12914, \a[17] , n_11064);
  not g23599 (n_11065, n12914);
  and g23600 (n12915, \a[17] , n_11065);
  and g23601 (n12916, n_11064, n_11065);
  not g23602 (n_11066, n12915);
  not g23603 (n_11067, n12916);
  and g23604 (n12917, n_11066, n_11067);
  and g23605 (n12918, n12906, n12917);
  not g23606 (n_11068, n12906);
  not g23607 (n_11069, n12917);
  and g23608 (n12919, n_11068, n_11069);
  not g23609 (n_11070, n12918);
  not g23610 (n_11071, n12919);
  and g23611 (n12920, n_11070, n_11071);
  not g23612 (n_11072, n12615);
  and g23613 (n12921, n_11072, n12920);
  not g23614 (n_11073, n12920);
  and g23615 (n12922, n12615, n_11073);
  not g23616 (n_11074, n12921);
  not g23617 (n_11075, n12922);
  and g23618 (n12923, n_11074, n_11075);
  not g23619 (n_11076, n12923);
  and g23620 (n12924, n12614, n_11076);
  not g23621 (n_11077, n12614);
  and g23622 (n12925, n_11077, n12923);
  not g23623 (n_11078, n12924);
  not g23624 (n_11079, n12925);
  and g23625 (n12926, n_11078, n_11079);
  not g23626 (n_11080, n12603);
  and g23627 (n12927, n_11080, n12926);
  not g23628 (n_11081, n12926);
  and g23629 (n12928, n12603, n_11081);
  not g23630 (n_11082, n12927);
  not g23631 (n_11083, n12928);
  and g23632 (n12929, n_11082, n_11083);
  not g23633 (n_11084, n12929);
  and g23634 (n12930, n12602, n_11084);
  not g23635 (n_11085, n12602);
  and g23636 (n12931, n_11085, n12929);
  not g23637 (n_11086, n12930);
  not g23638 (n_11087, n12931);
  and g23639 (n12932, n_11086, n_11087);
  not g23640 (n_11088, n12591);
  and g23641 (n12933, n_11088, n12932);
  not g23642 (n_11089, n12932);
  and g23643 (n12934, n12591, n_11089);
  not g23644 (n_11090, n12933);
  not g23645 (n_11091, n12934);
  and g23646 (n12935, n_11090, n_11091);
  not g23647 (n_11092, n12590);
  and g23648 (n12936, n_11092, n12935);
  not g23649 (n_11093, n12936);
  and g23650 (n12937, n12935, n_11093);
  and g23651 (n12938, n_11092, n_11093);
  not g23652 (n_11094, n12937);
  not g23653 (n_11095, n12938);
  and g23654 (n12939, n_11094, n_11095);
  and g23655 (n12940, n_10764, n_10768);
  and g23656 (n12941, n12939, n12940);
  not g23657 (n_11096, n12939);
  not g23658 (n_11097, n12940);
  and g23659 (n12942, n_11096, n_11097);
  not g23660 (n_11098, n12941);
  not g23661 (n_11099, n12942);
  and g23662 (n12943, n_11098, n_11099);
  and g23663 (n12944, \b[58] , n362);
  and g23664 (n12945, \b[56] , n403);
  and g23665 (n12946, \b[57] , n357);
  and g23671 (n12949, n365, n11436);
  not g23674 (n_11104, n12950);
  and g23675 (n12951, \a[5] , n_11104);
  not g23676 (n_11105, n12951);
  and g23677 (n12952, \a[5] , n_11105);
  and g23678 (n12953, n_11104, n_11105);
  not g23679 (n_11106, n12952);
  not g23680 (n_11107, n12953);
  and g23681 (n12954, n_11106, n_11107);
  not g23682 (n_11108, n12943);
  and g23683 (n12955, n_11108, n12954);
  not g23684 (n_11109, n12954);
  and g23685 (n12956, n12943, n_11109);
  not g23686 (n_11110, n12955);
  not g23687 (n_11111, n12956);
  and g23688 (n12957, n_11110, n_11111);
  and g23689 (n12958, \b[61] , n266);
  and g23690 (n12959, \b[59] , n284);
  and g23691 (n12960, \b[60] , n261);
  and g23697 (n12963, n_10458, n_10461);
  not g23698 (n_11116, \b[61] );
  and g23699 (n12964, n_10456, n_11116);
  and g23700 (n12965, \b[60] , \b[61] );
  not g23701 (n_11117, n12964);
  not g23702 (n_11118, n12965);
  and g23703 (n12966, n_11117, n_11118);
  not g23704 (n_11119, n12963);
  and g23705 (n12967, n_11119, n12966);
  not g23706 (n_11120, n12966);
  and g23707 (n12968, n12963, n_11120);
  not g23708 (n_11121, n12967);
  not g23709 (n_11122, n12968);
  and g23710 (n12969, n_11121, n_11122);
  and g23711 (n12970, n269, n12969);
  not g23714 (n_11124, n12971);
  and g23715 (n12972, \a[2] , n_11124);
  not g23716 (n_11125, n12972);
  and g23717 (n12973, \a[2] , n_11125);
  and g23718 (n12974, n_11124, n_11125);
  not g23719 (n_11126, n12973);
  not g23720 (n_11127, n12974);
  and g23721 (n12975, n_11126, n_11127);
  not g23722 (n_11128, n12975);
  and g23723 (n12976, n12957, n_11128);
  not g23724 (n_11129, n12976);
  and g23725 (n12977, n12957, n_11129);
  and g23726 (n12978, n_11128, n_11129);
  not g23727 (n_11130, n12977);
  not g23728 (n_11131, n12978);
  and g23729 (n12979, n_11130, n_11131);
  and g23730 (n12980, n_10772, n_10776);
  and g23731 (n12981, n12979, n12980);
  not g23732 (n_11132, n12979);
  not g23733 (n_11133, n12980);
  and g23734 (n12982, n_11132, n_11133);
  not g23735 (n_11134, n12981);
  not g23736 (n_11135, n12982);
  and g23737 (n12983, n_11134, n_11135);
  and g23738 (n12984, n_10780, n_10784);
  not g23739 (n_11136, n12984);
  and g23740 (n12985, n12983, n_11136);
  not g23741 (n_11137, n12983);
  and g23742 (n12986, n_11137, n12984);
  not g23743 (n_11138, n12985);
  not g23744 (n_11139, n12986);
  and g23745 (\f[61] , n_11138, n_11139);
  and g23746 (n12988, n_11135, n_11138);
  and g23747 (n12989, n_11111, n_11129);
  and g23748 (n12990, n_11087, n_11090);
  and g23749 (n12991, n_11079, n_11082);
  and g23750 (n12992, \b[50] , n951);
  and g23751 (n12993, \b[48] , n1056);
  and g23752 (n12994, \b[49] , n946);
  and g23758 (n12997, n954, n8949);
  not g23761 (n_11144, n12998);
  and g23762 (n12999, \a[14] , n_11144);
  not g23763 (n_11145, n12999);
  and g23764 (n13000, \a[14] , n_11145);
  and g23765 (n13001, n_11144, n_11145);
  not g23766 (n_11146, n13000);
  not g23767 (n_11147, n13001);
  and g23768 (n13002, n_11146, n_11147);
  and g23769 (n13003, n_11071, n_11074);
  and g23770 (n13004, n_11037, n_11043);
  and g23771 (n13005, n_10992, n_10993);
  not g23772 (n_11148, n13005);
  and g23773 (n13006, n_10989, n_11148);
  and g23774 (n13007, n_10941, n_10947);
  and g23775 (n13008, n_10908, n_10914);
  and g23776 (n13009, \b[17] , n7446);
  and g23777 (n13010, \b[15] , n7787);
  and g23778 (n13011, \b[16] , n7441);
  and g23784 (n13014, n1356, n7449);
  not g23787 (n_11153, n13015);
  and g23788 (n13016, \a[47] , n_11153);
  not g23789 (n_11154, n13016);
  and g23790 (n13017, \a[47] , n_11154);
  and g23791 (n13018, n_11153, n_11154);
  not g23792 (n_11155, n13017);
  not g23793 (n_11156, n13018);
  and g23794 (n13019, n_11155, n_11156);
  and g23795 (n13020, \b[14] , n8362);
  and g23796 (n13021, \b[12] , n8715);
  and g23797 (n13022, \b[13] , n8357);
  and g23803 (n13025, n1034, n8365);
  not g23806 (n_11161, n13026);
  and g23807 (n13027, \a[50] , n_11161);
  not g23808 (n_11162, n13027);
  and g23809 (n13028, \a[50] , n_11162);
  and g23810 (n13029, n_11161, n_11162);
  not g23811 (n_11163, n13028);
  not g23812 (n_11164, n13029);
  and g23813 (n13030, n_11163, n_11164);
  and g23814 (n13031, n_10875, n_10881);
  and g23815 (n13032, \b[11] , n9339);
  and g23816 (n13033, \b[9] , n9732);
  and g23817 (n13034, \b[10] , n9334);
  and g23823 (n13037, n818, n9342);
  not g23826 (n_11169, n13038);
  and g23827 (n13039, \a[53] , n_11169);
  not g23828 (n_11170, n13039);
  and g23829 (n13040, \a[53] , n_11170);
  and g23830 (n13041, n_11169, n_11170);
  not g23831 (n_11171, n13040);
  not g23832 (n_11172, n13041);
  and g23833 (n13042, n_11171, n_11172);
  and g23834 (n13043, n_10869, n_10872);
  and g23835 (n13044, n_10861, n_10864);
  and g23836 (n13045, \b[2] , n12668);
  and g23837 (n13046, n12354, n_10848);
  and g23838 (n13047, n12662, n13046);
  and g23839 (n13048, \b[0] , n13047);
  and g23840 (n13049, \b[1] , n12663);
  and g23846 (n13052, n296, n12671);
  not g23849 (n_11177, n13053);
  and g23850 (n13054, \a[62] , n_11177);
  not g23851 (n_11178, n13054);
  and g23852 (n13055, \a[62] , n_11178);
  and g23853 (n13056, n_11177, n_11178);
  not g23854 (n_11179, n13055);
  not g23855 (n_11180, n13056);
  and g23856 (n13057, n_11179, n_11180);
  and g23857 (n13058, n_10856, n13057);
  not g23858 (n_11181, n13057);
  and g23859 (n13059, n12678, n_11181);
  not g23860 (n_11182, n13058);
  not g23861 (n_11183, n13059);
  and g23862 (n13060, n_11182, n_11183);
  and g23863 (n13061, \b[5] , n11531);
  and g23864 (n13062, \b[3] , n11896);
  and g23865 (n13063, \b[4] , n11526);
  and g23871 (n13066, n394, n11534);
  not g23874 (n_11188, n13067);
  and g23875 (n13068, \a[59] , n_11188);
  not g23876 (n_11189, n13068);
  and g23877 (n13069, \a[59] , n_11189);
  and g23878 (n13070, n_11188, n_11189);
  not g23879 (n_11190, n13069);
  not g23880 (n_11191, n13070);
  and g23881 (n13071, n_11190, n_11191);
  not g23882 (n_11192, n13071);
  and g23883 (n13072, n13060, n_11192);
  not g23884 (n_11193, n13060);
  and g23885 (n13073, n_11193, n13071);
  not g23886 (n_11194, n13044);
  not g23887 (n_11195, n13073);
  and g23888 (n13074, n_11194, n_11195);
  not g23889 (n_11196, n13072);
  and g23890 (n13075, n_11196, n13074);
  not g23891 (n_11197, n13075);
  and g23892 (n13076, n_11194, n_11197);
  and g23893 (n13077, n_11196, n_11197);
  and g23894 (n13078, n_11195, n13077);
  not g23895 (n_11198, n13076);
  not g23896 (n_11199, n13078);
  and g23897 (n13079, n_11198, n_11199);
  and g23898 (n13080, \b[8] , n10426);
  and g23899 (n13081, \b[6] , n10796);
  and g23900 (n13082, \b[7] , n10421);
  and g23906 (n13085, n585, n10429);
  not g23909 (n_11204, n13086);
  and g23910 (n13087, \a[56] , n_11204);
  not g23911 (n_11205, n13087);
  and g23912 (n13088, \a[56] , n_11205);
  and g23913 (n13089, n_11204, n_11205);
  not g23914 (n_11206, n13088);
  not g23915 (n_11207, n13089);
  and g23916 (n13090, n_11206, n_11207);
  and g23917 (n13091, n13079, n13090);
  not g23918 (n_11208, n13079);
  not g23919 (n_11209, n13090);
  and g23920 (n13092, n_11208, n_11209);
  not g23921 (n_11210, n13091);
  not g23922 (n_11211, n13092);
  and g23923 (n13093, n_11210, n_11211);
  not g23924 (n_11212, n13043);
  and g23925 (n13094, n_11212, n13093);
  not g23926 (n_11213, n13093);
  and g23927 (n13095, n13043, n_11213);
  not g23928 (n_11214, n13094);
  not g23929 (n_11215, n13095);
  and g23930 (n13096, n_11214, n_11215);
  not g23931 (n_11216, n13096);
  and g23932 (n13097, n13042, n_11216);
  not g23933 (n_11217, n13042);
  and g23934 (n13098, n_11217, n13096);
  not g23935 (n_11218, n13097);
  not g23936 (n_11219, n13098);
  and g23937 (n13099, n_11218, n_11219);
  not g23938 (n_11220, n13031);
  and g23939 (n13100, n_11220, n13099);
  not g23940 (n_11221, n13099);
  and g23941 (n13101, n13031, n_11221);
  not g23942 (n_11222, n13100);
  not g23943 (n_11223, n13101);
  and g23944 (n13102, n_11222, n_11223);
  not g23945 (n_11224, n13030);
  and g23946 (n13103, n_11224, n13102);
  not g23947 (n_11225, n13103);
  and g23948 (n13104, n13102, n_11225);
  and g23949 (n13105, n_11224, n_11225);
  not g23950 (n_11226, n13104);
  not g23951 (n_11227, n13105);
  and g23952 (n13106, n_11226, n_11227);
  not g23953 (n_11228, n12717);
  not g23954 (n_11229, n13106);
  and g23955 (n13107, n_11228, n_11229);
  and g23956 (n13108, n12717, n13106);
  not g23957 (n_11230, n13107);
  not g23958 (n_11231, n13108);
  and g23959 (n13109, n_11230, n_11231);
  not g23960 (n_11232, n13019);
  and g23961 (n13110, n_11232, n13109);
  not g23962 (n_11233, n13110);
  and g23963 (n13111, n_11232, n_11233);
  and g23964 (n13112, n13109, n_11233);
  not g23965 (n_11234, n13111);
  not g23966 (n_11235, n13112);
  and g23967 (n13113, n_11234, n_11235);
  not g23968 (n_11236, n13008);
  not g23969 (n_11237, n13113);
  and g23970 (n13114, n_11236, n_11237);
  not g23971 (n_11238, n13114);
  and g23972 (n13115, n_11236, n_11238);
  and g23973 (n13116, n_11237, n_11238);
  not g23974 (n_11239, n13115);
  not g23975 (n_11240, n13116);
  and g23976 (n13117, n_11239, n_11240);
  and g23977 (n13118, \b[20] , n6595);
  and g23978 (n13119, \b[18] , n6902);
  and g23979 (n13120, \b[19] , n6590);
  and g23985 (n13123, n1846, n6598);
  not g23988 (n_11245, n13124);
  and g23989 (n13125, \a[44] , n_11245);
  not g23990 (n_11246, n13125);
  and g23991 (n13126, \a[44] , n_11246);
  and g23992 (n13127, n_11245, n_11246);
  not g23993 (n_11247, n13126);
  not g23994 (n_11248, n13127);
  and g23995 (n13128, n_11247, n_11248);
  not g23996 (n_11249, n13117);
  not g23997 (n_11250, n13128);
  and g23998 (n13129, n_11249, n_11250);
  not g23999 (n_11251, n13129);
  and g24000 (n13130, n_11249, n_11251);
  and g24001 (n13131, n_11250, n_11251);
  not g24002 (n_11252, n13130);
  not g24003 (n_11253, n13131);
  and g24004 (n13132, n_11252, n_11253);
  not g24005 (n_11254, n12755);
  and g24006 (n13133, n_11254, n13132);
  not g24007 (n_11255, n13132);
  and g24008 (n13134, n12755, n_11255);
  not g24009 (n_11256, n13133);
  not g24010 (n_11257, n13134);
  and g24011 (n13135, n_11256, n_11257);
  and g24012 (n13136, \b[23] , n5777);
  and g24013 (n13137, \b[21] , n6059);
  and g24014 (n13138, \b[22] , n5772);
  and g24020 (n13141, n2300, n5780);
  not g24023 (n_11262, n13142);
  and g24024 (n13143, \a[41] , n_11262);
  not g24025 (n_11263, n13143);
  and g24026 (n13144, \a[41] , n_11263);
  and g24027 (n13145, n_11262, n_11263);
  not g24028 (n_11264, n13144);
  not g24029 (n_11265, n13145);
  and g24030 (n13146, n_11264, n_11265);
  not g24031 (n_11266, n13135);
  not g24032 (n_11267, n13146);
  and g24033 (n13147, n_11266, n_11267);
  and g24034 (n13148, n13135, n13146);
  not g24035 (n_11268, n13147);
  not g24036 (n_11269, n13148);
  and g24037 (n13149, n_11268, n_11269);
  not g24038 (n_11270, n13149);
  and g24039 (n13150, n13007, n_11270);
  not g24040 (n_11271, n13007);
  and g24041 (n13151, n_11271, n13149);
  not g24042 (n_11272, n13150);
  not g24043 (n_11273, n13151);
  and g24044 (n13152, n_11272, n_11273);
  and g24045 (n13153, \b[26] , n5035);
  and g24046 (n13154, \b[24] , n5277);
  and g24047 (n13155, \b[25] , n5030);
  and g24053 (n13158, n2813, n5038);
  not g24056 (n_11278, n13159);
  and g24057 (n13160, \a[38] , n_11278);
  not g24058 (n_11279, n13160);
  and g24059 (n13161, \a[38] , n_11279);
  and g24060 (n13162, n_11278, n_11279);
  not g24061 (n_11280, n13161);
  not g24062 (n_11281, n13162);
  and g24063 (n13163, n_11280, n_11281);
  not g24064 (n_11282, n13163);
  and g24065 (n13164, n13152, n_11282);
  not g24066 (n_11283, n13164);
  and g24067 (n13165, n13152, n_11283);
  and g24068 (n13166, n_11282, n_11283);
  not g24069 (n_11284, n13165);
  not g24070 (n_11285, n13166);
  and g24071 (n13167, n_11284, n_11285);
  and g24072 (n13168, n_10957, n_10963);
  and g24073 (n13169, n13167, n13168);
  not g24074 (n_11286, n13167);
  not g24075 (n_11287, n13168);
  and g24076 (n13170, n_11286, n_11287);
  not g24077 (n_11288, n13169);
  not g24078 (n_11289, n13170);
  and g24079 (n13171, n_11288, n_11289);
  and g24080 (n13172, \b[29] , n4287);
  and g24081 (n13173, \b[27] , n4532);
  and g24082 (n13174, \b[28] , n4282);
  and g24088 (n13177, n3383, n4290);
  not g24091 (n_11294, n13178);
  and g24092 (n13179, \a[35] , n_11294);
  not g24093 (n_11295, n13179);
  and g24094 (n13180, \a[35] , n_11295);
  and g24095 (n13181, n_11294, n_11295);
  not g24096 (n_11296, n13180);
  not g24097 (n_11297, n13181);
  and g24098 (n13182, n_11296, n_11297);
  not g24099 (n_11298, n13182);
  and g24100 (n13183, n13171, n_11298);
  not g24101 (n_11299, n13183);
  and g24102 (n13184, n13171, n_11299);
  and g24103 (n13185, n_11298, n_11299);
  not g24104 (n_11300, n13184);
  not g24105 (n_11301, n13185);
  and g24106 (n13186, n_11300, n_11301);
  and g24107 (n13187, n_10973, n_10979);
  and g24108 (n13188, n13186, n13187);
  not g24109 (n_11302, n13186);
  not g24110 (n_11303, n13187);
  and g24111 (n13189, n_11302, n_11303);
  not g24112 (n_11304, n13188);
  not g24113 (n_11305, n13189);
  and g24114 (n13190, n_11304, n_11305);
  and g24115 (n13191, \b[32] , n3638);
  and g24116 (n13192, \b[30] , n3843);
  and g24117 (n13193, \b[31] , n3633);
  and g24123 (n13196, n3641, n4013);
  not g24126 (n_11310, n13197);
  and g24127 (n13198, \a[32] , n_11310);
  not g24128 (n_11311, n13198);
  and g24129 (n13199, \a[32] , n_11311);
  and g24130 (n13200, n_11310, n_11311);
  not g24131 (n_11312, n13199);
  not g24132 (n_11313, n13200);
  and g24133 (n13201, n_11312, n_11313);
  not g24134 (n_11314, n13201);
  and g24135 (n13202, n13190, n_11314);
  not g24136 (n_11315, n13190);
  and g24137 (n13203, n_11315, n13201);
  not g24138 (n_11316, n13006);
  not g24139 (n_11317, n13203);
  and g24140 (n13204, n_11316, n_11317);
  not g24141 (n_11318, n13202);
  and g24142 (n13205, n_11318, n13204);
  not g24143 (n_11319, n13205);
  and g24144 (n13206, n_11316, n_11319);
  and g24145 (n13207, n_11318, n_11319);
  and g24146 (n13208, n_11317, n13207);
  not g24147 (n_11320, n13206);
  not g24148 (n_11321, n13208);
  and g24149 (n13209, n_11320, n_11321);
  and g24150 (n13210, \b[35] , n3050);
  and g24151 (n13211, \b[33] , n3243);
  and g24152 (n13212, \b[34] , n3045);
  and g24158 (n13215, n3053, n4696);
  not g24161 (n_11326, n13216);
  and g24162 (n13217, \a[29] , n_11326);
  not g24163 (n_11327, n13217);
  and g24164 (n13218, \a[29] , n_11327);
  and g24165 (n13219, n_11326, n_11327);
  not g24166 (n_11328, n13218);
  not g24167 (n_11329, n13219);
  and g24168 (n13220, n_11328, n_11329);
  not g24169 (n_11330, n13209);
  not g24170 (n_11331, n13220);
  and g24171 (n13221, n_11330, n_11331);
  not g24172 (n_11332, n13221);
  and g24173 (n13222, n_11330, n_11332);
  and g24174 (n13223, n_11331, n_11332);
  not g24175 (n_11333, n13222);
  not g24176 (n_11334, n13223);
  and g24177 (n13224, n_11333, n_11334);
  and g24178 (n13225, n_11006, n_11011);
  and g24179 (n13226, n13224, n13225);
  not g24180 (n_11335, n13224);
  not g24181 (n_11336, n13225);
  and g24182 (n13227, n_11335, n_11336);
  not g24183 (n_11337, n13226);
  not g24184 (n_11338, n13227);
  and g24185 (n13228, n_11337, n_11338);
  and g24186 (n13229, \b[38] , n2539);
  and g24187 (n13230, \b[36] , n2685);
  and g24188 (n13231, \b[37] , n2534);
  and g24194 (n13234, n2542, n5205);
  not g24197 (n_11343, n13235);
  and g24198 (n13236, \a[26] , n_11343);
  not g24199 (n_11344, n13236);
  and g24200 (n13237, \a[26] , n_11344);
  and g24201 (n13238, n_11343, n_11344);
  not g24202 (n_11345, n13237);
  not g24203 (n_11346, n13238);
  and g24204 (n13239, n_11345, n_11346);
  not g24205 (n_11347, n13239);
  and g24206 (n13240, n13228, n_11347);
  not g24207 (n_11348, n13240);
  and g24208 (n13241, n13228, n_11348);
  and g24209 (n13242, n_11347, n_11348);
  not g24210 (n_11349, n13241);
  not g24211 (n_11350, n13242);
  and g24212 (n13243, n_11349, n_11350);
  and g24213 (n13244, n_11021, n_11027);
  and g24214 (n13245, n13243, n13244);
  not g24215 (n_11351, n13243);
  not g24216 (n_11352, n13244);
  and g24217 (n13246, n_11351, n_11352);
  not g24218 (n_11353, n13245);
  not g24219 (n_11354, n13246);
  and g24220 (n13247, n_11353, n_11354);
  and g24221 (n13248, \b[41] , n2048);
  and g24222 (n13249, \b[39] , n2198);
  and g24223 (n13250, \b[40] , n2043);
  and g24229 (n13253, n2051, n6219);
  not g24232 (n_11359, n13254);
  and g24233 (n13255, \a[23] , n_11359);
  not g24234 (n_11360, n13255);
  and g24235 (n13256, \a[23] , n_11360);
  and g24236 (n13257, n_11359, n_11360);
  not g24237 (n_11361, n13256);
  not g24238 (n_11362, n13257);
  and g24239 (n13258, n_11361, n_11362);
  not g24240 (n_11363, n13258);
  and g24241 (n13259, n13247, n_11363);
  not g24242 (n_11364, n13247);
  and g24243 (n13260, n_11364, n13258);
  not g24244 (n_11365, n13004);
  not g24245 (n_11366, n13260);
  and g24246 (n13261, n_11365, n_11366);
  not g24247 (n_11367, n13259);
  and g24248 (n13262, n_11367, n13261);
  not g24249 (n_11368, n13262);
  and g24250 (n13263, n_11365, n_11368);
  and g24251 (n13264, n_11367, n_11368);
  and g24252 (n13265, n_11366, n13264);
  not g24253 (n_11369, n13263);
  not g24254 (n_11370, n13265);
  and g24255 (n13266, n_11369, n_11370);
  and g24256 (n13267, \b[44] , n1627);
  and g24257 (n13268, \b[42] , n1763);
  and g24258 (n13269, \b[43] , n1622);
  and g24264 (n13272, n1630, n7072);
  not g24267 (n_11375, n13273);
  and g24268 (n13274, \a[20] , n_11375);
  not g24269 (n_11376, n13274);
  and g24270 (n13275, \a[20] , n_11376);
  and g24271 (n13276, n_11375, n_11376);
  not g24272 (n_11377, n13275);
  not g24273 (n_11378, n13276);
  and g24274 (n13277, n_11377, n_11378);
  not g24275 (n_11379, n13266);
  not g24276 (n_11380, n13277);
  and g24277 (n13278, n_11379, n_11380);
  not g24278 (n_11381, n13278);
  and g24279 (n13279, n_11379, n_11381);
  and g24280 (n13280, n_11380, n_11381);
  not g24281 (n_11382, n13279);
  not g24282 (n_11383, n13280);
  and g24283 (n13281, n_11382, n_11383);
  not g24284 (n_11384, n12904);
  and g24285 (n13282, n_11384, n13281);
  not g24286 (n_11385, n13281);
  and g24287 (n13283, n12904, n_11385);
  not g24288 (n_11386, n13282);
  not g24289 (n_11387, n13283);
  and g24290 (n13284, n_11386, n_11387);
  and g24291 (n13285, \b[47] , n1302);
  and g24292 (n13286, \b[45] , n1391);
  and g24293 (n13287, \b[46] , n1297);
  and g24299 (n13290, n1305, n7703);
  not g24302 (n_11392, n13291);
  and g24303 (n13292, \a[17] , n_11392);
  not g24304 (n_11393, n13292);
  and g24305 (n13293, \a[17] , n_11393);
  and g24306 (n13294, n_11392, n_11393);
  not g24307 (n_11394, n13293);
  not g24308 (n_11395, n13294);
  and g24309 (n13295, n_11394, n_11395);
  not g24310 (n_11396, n13284);
  not g24311 (n_11397, n13295);
  and g24312 (n13296, n_11396, n_11397);
  and g24313 (n13297, n13284, n13295);
  not g24314 (n_11398, n13296);
  not g24315 (n_11399, n13297);
  and g24316 (n13298, n_11398, n_11399);
  not g24317 (n_11400, n13003);
  and g24318 (n13299, n_11400, n13298);
  not g24319 (n_11401, n13298);
  and g24320 (n13300, n13003, n_11401);
  not g24321 (n_11402, n13299);
  not g24322 (n_11403, n13300);
  and g24323 (n13301, n_11402, n_11403);
  not g24324 (n_11404, n13002);
  and g24325 (n13302, n_11404, n13301);
  not g24326 (n_11405, n13302);
  and g24327 (n13303, n13301, n_11405);
  and g24328 (n13304, n_11404, n_11405);
  not g24329 (n_11406, n13303);
  not g24330 (n_11407, n13304);
  and g24331 (n13305, n_11406, n_11407);
  not g24332 (n_11408, n12991);
  and g24333 (n13306, n_11408, n13305);
  not g24334 (n_11409, n13305);
  and g24335 (n13307, n12991, n_11409);
  not g24336 (n_11410, n13306);
  not g24337 (n_11411, n13307);
  and g24338 (n13308, n_11410, n_11411);
  and g24339 (n13309, \b[53] , n700);
  and g24340 (n13310, \b[51] , n767);
  and g24341 (n13311, \b[52] , n695);
  and g24347 (n13314, n703, n9972);
  not g24350 (n_11416, n13315);
  and g24351 (n13316, \a[11] , n_11416);
  not g24352 (n_11417, n13316);
  and g24353 (n13317, \a[11] , n_11417);
  and g24354 (n13318, n_11416, n_11417);
  not g24355 (n_11418, n13317);
  not g24356 (n_11419, n13318);
  and g24357 (n13319, n_11418, n_11419);
  not g24358 (n_11420, n13308);
  not g24359 (n_11421, n13319);
  and g24360 (n13320, n_11420, n_11421);
  and g24361 (n13321, n13308, n13319);
  not g24362 (n_11422, n13320);
  not g24363 (n_11423, n13321);
  and g24364 (n13322, n_11422, n_11423);
  not g24365 (n_11424, n12990);
  and g24366 (n13323, n_11424, n13322);
  not g24367 (n_11425, n13322);
  and g24368 (n13324, n12990, n_11425);
  not g24369 (n_11426, n13323);
  not g24370 (n_11427, n13324);
  and g24371 (n13325, n_11426, n_11427);
  and g24372 (n13326, \b[56] , n511);
  and g24373 (n13327, \b[54] , n541);
  and g24374 (n13328, \b[55] , n506);
  and g24380 (n13331, n514, n10708);
  not g24383 (n_11432, n13332);
  and g24384 (n13333, \a[8] , n_11432);
  not g24385 (n_11433, n13333);
  and g24386 (n13334, \a[8] , n_11433);
  and g24387 (n13335, n_11432, n_11433);
  not g24388 (n_11434, n13334);
  not g24389 (n_11435, n13335);
  and g24390 (n13336, n_11434, n_11435);
  not g24391 (n_11436, n13325);
  and g24392 (n13337, n_11436, n13336);
  not g24393 (n_11437, n13336);
  and g24394 (n13338, n13325, n_11437);
  not g24395 (n_11438, n13337);
  not g24396 (n_11439, n13338);
  and g24397 (n13339, n_11438, n_11439);
  and g24398 (n13340, \b[59] , n362);
  and g24399 (n13341, \b[57] , n403);
  and g24400 (n13342, \b[58] , n357);
  and g24406 (n13345, n365, n12179);
  not g24409 (n_11444, n13346);
  and g24410 (n13347, \a[5] , n_11444);
  not g24411 (n_11445, n13347);
  and g24412 (n13348, \a[5] , n_11445);
  and g24413 (n13349, n_11444, n_11445);
  not g24414 (n_11446, n13348);
  not g24415 (n_11447, n13349);
  and g24416 (n13350, n_11446, n_11447);
  not g24417 (n_11448, n13350);
  and g24418 (n13351, n13339, n_11448);
  not g24419 (n_11449, n13351);
  and g24420 (n13352, n13339, n_11449);
  and g24421 (n13353, n_11448, n_11449);
  not g24422 (n_11450, n13352);
  not g24423 (n_11451, n13353);
  and g24424 (n13354, n_11450, n_11451);
  and g24425 (n13355, n_11093, n_11099);
  and g24426 (n13356, n13354, n13355);
  not g24427 (n_11452, n13354);
  not g24428 (n_11453, n13355);
  and g24429 (n13357, n_11452, n_11453);
  not g24430 (n_11454, n13356);
  not g24431 (n_11455, n13357);
  and g24432 (n13358, n_11454, n_11455);
  and g24433 (n13359, \b[62] , n266);
  and g24434 (n13360, \b[60] , n284);
  and g24435 (n13361, \b[61] , n261);
  and g24441 (n13364, n_11118, n_11121);
  not g24442 (n_11460, \b[62] );
  and g24443 (n13365, n_11116, n_11460);
  and g24444 (n13366, \b[61] , \b[62] );
  not g24445 (n_11461, n13365);
  not g24446 (n_11462, n13366);
  and g24447 (n13367, n_11461, n_11462);
  not g24448 (n_11463, n13364);
  and g24449 (n13368, n_11463, n13367);
  not g24450 (n_11464, n13367);
  and g24451 (n13369, n13364, n_11464);
  not g24452 (n_11465, n13368);
  not g24453 (n_11466, n13369);
  and g24454 (n13370, n_11465, n_11466);
  and g24455 (n13371, n269, n13370);
  not g24458 (n_11468, n13372);
  and g24459 (n13373, \a[2] , n_11468);
  not g24460 (n_11469, n13373);
  and g24461 (n13374, \a[2] , n_11469);
  and g24462 (n13375, n_11468, n_11469);
  not g24463 (n_11470, n13374);
  not g24464 (n_11471, n13375);
  and g24465 (n13376, n_11470, n_11471);
  not g24466 (n_11472, n13358);
  and g24467 (n13377, n_11472, n13376);
  not g24468 (n_11473, n13376);
  and g24469 (n13378, n13358, n_11473);
  not g24470 (n_11474, n13377);
  not g24471 (n_11475, n13378);
  and g24472 (n13379, n_11474, n_11475);
  not g24473 (n_11476, n12989);
  and g24474 (n13380, n_11476, n13379);
  not g24475 (n_11477, n13379);
  and g24476 (n13381, n12989, n_11477);
  not g24477 (n_11478, n13380);
  not g24478 (n_11479, n13381);
  and g24479 (n13382, n_11478, n_11479);
  not g24480 (n_11480, n12988);
  and g24481 (n13383, n_11480, n13382);
  not g24482 (n_11481, n13382);
  and g24483 (n13384, n12988, n_11481);
  not g24484 (n_11482, n13383);
  not g24485 (n_11483, n13384);
  and g24486 (\f[62] , n_11482, n_11483);
  and g24487 (n13386, n_11408, n_11409);
  not g24488 (n_11484, n13386);
  and g24489 (n13387, n_11405, n_11484);
  and g24490 (n13388, \b[51] , n951);
  and g24491 (n13389, \b[49] , n1056);
  and g24492 (n13390, \b[50] , n946);
  and g24498 (n13393, n954, n8976);
  not g24501 (n_11489, n13394);
  and g24502 (n13395, \a[14] , n_11489);
  not g24503 (n_11490, n13395);
  and g24504 (n13396, \a[14] , n_11490);
  and g24505 (n13397, n_11489, n_11490);
  not g24506 (n_11491, n13396);
  not g24507 (n_11492, n13397);
  and g24508 (n13398, n_11491, n_11492);
  and g24509 (n13399, n_11398, n_11402);
  and g24510 (n13400, \b[48] , n1302);
  and g24511 (n13401, \b[46] , n1391);
  and g24512 (n13402, \b[47] , n1297);
  and g24518 (n13405, n1305, n8009);
  not g24521 (n_11497, n13406);
  and g24522 (n13407, \a[17] , n_11497);
  not g24523 (n_11498, n13407);
  and g24524 (n13408, \a[17] , n_11498);
  and g24525 (n13409, n_11497, n_11498);
  not g24526 (n_11499, n13408);
  not g24527 (n_11500, n13409);
  and g24528 (n13410, n_11499, n_11500);
  and g24529 (n13411, n_11384, n_11385);
  not g24530 (n_11501, n13411);
  and g24531 (n13412, n_11381, n_11501);
  and g24532 (n13413, \b[45] , n1627);
  and g24533 (n13414, \b[43] , n1763);
  and g24534 (n13415, \b[44] , n1622);
  and g24540 (n13418, n1630, n7361);
  not g24543 (n_11506, n13419);
  and g24544 (n13420, \a[20] , n_11506);
  not g24545 (n_11507, n13420);
  and g24546 (n13421, \a[20] , n_11507);
  and g24547 (n13422, n_11506, n_11507);
  not g24548 (n_11508, n13421);
  not g24549 (n_11509, n13422);
  and g24550 (n13423, n_11508, n_11509);
  and g24551 (n13424, \b[42] , n2048);
  and g24552 (n13425, \b[40] , n2198);
  and g24553 (n13426, \b[41] , n2043);
  and g24559 (n13429, n2051, n6489);
  not g24562 (n_11514, n13430);
  and g24563 (n13431, \a[23] , n_11514);
  not g24564 (n_11515, n13431);
  and g24565 (n13432, \a[23] , n_11515);
  and g24566 (n13433, n_11514, n_11515);
  not g24567 (n_11516, n13432);
  not g24568 (n_11517, n13433);
  and g24569 (n13434, n_11516, n_11517);
  and g24570 (n13435, n_11348, n_11354);
  and g24571 (n13436, n_11332, n_11338);
  and g24572 (n13437, \b[33] , n3638);
  and g24573 (n13438, \b[31] , n3843);
  and g24574 (n13439, \b[32] , n3633);
  and g24580 (n13442, n3641, n4223);
  not g24583 (n_11522, n13443);
  and g24584 (n13444, \a[32] , n_11522);
  not g24585 (n_11523, n13444);
  and g24586 (n13445, \a[32] , n_11523);
  and g24587 (n13446, n_11522, n_11523);
  not g24588 (n_11524, n13445);
  not g24589 (n_11525, n13446);
  and g24590 (n13447, n_11524, n_11525);
  and g24591 (n13448, n_11254, n_11255);
  not g24592 (n_11526, n13448);
  and g24593 (n13449, n_11251, n_11526);
  and g24594 (n13450, \b[21] , n6595);
  and g24595 (n13451, \b[19] , n6902);
  and g24596 (n13452, \b[20] , n6590);
  and g24602 (n13455, n1984, n6598);
  not g24605 (n_11531, n13456);
  and g24606 (n13457, \a[44] , n_11531);
  not g24607 (n_11532, n13457);
  and g24608 (n13458, \a[44] , n_11532);
  and g24609 (n13459, n_11531, n_11532);
  not g24610 (n_11533, n13458);
  not g24611 (n_11534, n13459);
  and g24612 (n13460, n_11533, n_11534);
  and g24613 (n13461, n_11233, n_11238);
  and g24614 (n13462, \b[15] , n8362);
  and g24615 (n13463, \b[13] , n8715);
  and g24616 (n13464, \b[14] , n8357);
  and g24622 (n13467, n1131, n8365);
  not g24625 (n_11539, n13468);
  and g24626 (n13469, \a[50] , n_11539);
  not g24627 (n_11540, n13469);
  and g24628 (n13470, \a[50] , n_11540);
  and g24629 (n13471, n_11539, n_11540);
  not g24630 (n_11541, n13470);
  not g24631 (n_11542, n13471);
  and g24632 (n13472, n_11541, n_11542);
  and g24633 (n13473, n_11219, n_11222);
  and g24634 (n13474, n_11211, n_11214);
  and g24635 (n13475, \b[9] , n10426);
  and g24636 (n13476, \b[7] , n10796);
  and g24637 (n13477, \b[8] , n10421);
  and g24643 (n13480, n651, n10429);
  not g24646 (n_11547, n13481);
  and g24647 (n13482, \a[56] , n_11547);
  not g24648 (n_11548, n13482);
  and g24649 (n13483, \a[56] , n_11548);
  and g24650 (n13484, n_11547, n_11548);
  not g24651 (n_11549, n13483);
  not g24652 (n_11550, n13484);
  and g24653 (n13485, n_11549, n_11550);
  not g24654 (n_11552, \a[63] );
  and g24655 (n13486, \a[62] , n_11552);
  and g24656 (n13487, n_10843, \a[63] );
  not g24657 (n_11553, n13486);
  not g24658 (n_11554, n13487);
  and g24659 (n13488, n_11553, n_11554);
  not g24660 (n_11555, n13488);
  and g24661 (n13489, \b[0] , n_11555);
  and g24662 (n13490, n13059, n13489);
  not g24663 (n_11556, n13490);
  and g24664 (n13491, n13059, n_11556);
  and g24665 (n13492, n13489, n_11556);
  not g24666 (n_11557, n13491);
  not g24667 (n_11558, n13492);
  and g24668 (n13493, n_11557, n_11558);
  and g24669 (n13494, \b[3] , n12668);
  and g24670 (n13495, \b[1] , n13047);
  and g24671 (n13496, \b[2] , n12663);
  and g24677 (n13499, n318, n12671);
  not g24680 (n_11563, n13500);
  and g24681 (n13501, \a[62] , n_11563);
  not g24682 (n_11564, n13501);
  and g24683 (n13502, \a[62] , n_11564);
  and g24684 (n13503, n_11563, n_11564);
  not g24685 (n_11565, n13502);
  not g24686 (n_11566, n13503);
  and g24687 (n13504, n_11565, n_11566);
  not g24688 (n_11567, n13493);
  not g24689 (n_11568, n13504);
  and g24690 (n13505, n_11567, n_11568);
  not g24691 (n_11569, n13505);
  and g24692 (n13506, n_11567, n_11569);
  and g24693 (n13507, n_11568, n_11569);
  not g24694 (n_11570, n13506);
  not g24695 (n_11571, n13507);
  and g24696 (n13508, n_11570, n_11571);
  and g24697 (n13509, \b[6] , n11531);
  and g24698 (n13510, \b[4] , n11896);
  and g24699 (n13511, \b[5] , n11526);
  and g24705 (n13514, n459, n11534);
  not g24708 (n_11576, n13515);
  and g24709 (n13516, \a[59] , n_11576);
  not g24710 (n_11577, n13516);
  and g24711 (n13517, \a[59] , n_11577);
  and g24712 (n13518, n_11576, n_11577);
  not g24713 (n_11578, n13517);
  not g24714 (n_11579, n13518);
  and g24715 (n13519, n_11578, n_11579);
  and g24716 (n13520, n13508, n13519);
  not g24717 (n_11580, n13508);
  not g24718 (n_11581, n13519);
  and g24719 (n13521, n_11580, n_11581);
  not g24720 (n_11582, n13520);
  not g24721 (n_11583, n13521);
  and g24722 (n13522, n_11582, n_11583);
  not g24723 (n_11584, n13077);
  and g24724 (n13523, n_11584, n13522);
  not g24725 (n_11585, n13522);
  and g24726 (n13524, n13077, n_11585);
  not g24727 (n_11586, n13523);
  not g24728 (n_11587, n13524);
  and g24729 (n13525, n_11586, n_11587);
  not g24730 (n_11588, n13485);
  and g24731 (n13526, n_11588, n13525);
  not g24732 (n_11589, n13526);
  and g24733 (n13527, n13525, n_11589);
  and g24734 (n13528, n_11588, n_11589);
  not g24735 (n_11590, n13527);
  not g24736 (n_11591, n13528);
  and g24737 (n13529, n_11590, n_11591);
  not g24738 (n_11592, n13474);
  and g24739 (n13530, n_11592, n13529);
  not g24740 (n_11593, n13529);
  and g24741 (n13531, n13474, n_11593);
  not g24742 (n_11594, n13530);
  not g24743 (n_11595, n13531);
  and g24744 (n13532, n_11594, n_11595);
  and g24745 (n13533, \b[12] , n9339);
  and g24746 (n13534, \b[10] , n9732);
  and g24747 (n13535, \b[11] , n9334);
  and g24753 (n13538, n842, n9342);
  not g24756 (n_11600, n13539);
  and g24757 (n13540, \a[53] , n_11600);
  not g24758 (n_11601, n13540);
  and g24759 (n13541, \a[53] , n_11601);
  and g24760 (n13542, n_11600, n_11601);
  not g24761 (n_11602, n13541);
  not g24762 (n_11603, n13542);
  and g24763 (n13543, n_11602, n_11603);
  and g24764 (n13544, n13532, n13543);
  not g24765 (n_11604, n13532);
  not g24766 (n_11605, n13543);
  and g24767 (n13545, n_11604, n_11605);
  not g24768 (n_11606, n13544);
  not g24769 (n_11607, n13545);
  and g24770 (n13546, n_11606, n_11607);
  not g24771 (n_11608, n13473);
  and g24772 (n13547, n_11608, n13546);
  not g24773 (n_11609, n13546);
  and g24774 (n13548, n13473, n_11609);
  not g24775 (n_11610, n13547);
  not g24776 (n_11611, n13548);
  and g24777 (n13549, n_11610, n_11611);
  not g24778 (n_11612, n13472);
  and g24779 (n13550, n_11612, n13549);
  not g24780 (n_11613, n13550);
  and g24781 (n13551, n13549, n_11613);
  and g24782 (n13552, n_11612, n_11613);
  not g24783 (n_11614, n13551);
  not g24784 (n_11615, n13552);
  and g24785 (n13553, n_11614, n_11615);
  and g24786 (n13554, n_11225, n_11230);
  and g24787 (n13555, n13553, n13554);
  not g24788 (n_11616, n13553);
  not g24789 (n_11617, n13554);
  and g24790 (n13556, n_11616, n_11617);
  not g24791 (n_11618, n13555);
  not g24792 (n_11619, n13556);
  and g24793 (n13557, n_11618, n_11619);
  and g24794 (n13558, \b[18] , n7446);
  and g24795 (n13559, \b[16] , n7787);
  and g24796 (n13560, \b[17] , n7441);
  and g24802 (n13563, n1566, n7449);
  not g24805 (n_11624, n13564);
  and g24806 (n13565, \a[47] , n_11624);
  not g24807 (n_11625, n13565);
  and g24808 (n13566, \a[47] , n_11625);
  and g24809 (n13567, n_11624, n_11625);
  not g24810 (n_11626, n13566);
  not g24811 (n_11627, n13567);
  and g24812 (n13568, n_11626, n_11627);
  not g24813 (n_11628, n13557);
  and g24814 (n13569, n_11628, n13568);
  not g24815 (n_11629, n13568);
  and g24816 (n13570, n13557, n_11629);
  not g24817 (n_11630, n13569);
  not g24818 (n_11631, n13570);
  and g24819 (n13571, n_11630, n_11631);
  not g24820 (n_11632, n13461);
  and g24821 (n13572, n_11632, n13571);
  not g24822 (n_11633, n13571);
  and g24823 (n13573, n13461, n_11633);
  not g24824 (n_11634, n13572);
  not g24825 (n_11635, n13573);
  and g24826 (n13574, n_11634, n_11635);
  not g24827 (n_11636, n13460);
  and g24828 (n13575, n_11636, n13574);
  not g24829 (n_11637, n13574);
  and g24830 (n13576, n13460, n_11637);
  not g24831 (n_11638, n13575);
  not g24832 (n_11639, n13576);
  and g24833 (n13577, n_11638, n_11639);
  not g24834 (n_11640, n13449);
  and g24835 (n13578, n_11640, n13577);
  not g24836 (n_11641, n13577);
  and g24837 (n13579, n13449, n_11641);
  not g24838 (n_11642, n13578);
  not g24839 (n_11643, n13579);
  and g24840 (n13580, n_11642, n_11643);
  and g24841 (n13581, \b[24] , n5777);
  and g24842 (n13582, \b[22] , n6059);
  and g24843 (n13583, \b[23] , n5772);
  and g24849 (n13586, n2458, n5780);
  not g24852 (n_11648, n13587);
  and g24853 (n13588, \a[41] , n_11648);
  not g24854 (n_11649, n13588);
  and g24855 (n13589, \a[41] , n_11649);
  and g24856 (n13590, n_11648, n_11649);
  not g24857 (n_11650, n13589);
  not g24858 (n_11651, n13590);
  and g24859 (n13591, n_11650, n_11651);
  not g24860 (n_11652, n13591);
  and g24861 (n13592, n13580, n_11652);
  not g24862 (n_11653, n13592);
  and g24863 (n13593, n13580, n_11653);
  and g24864 (n13594, n_11652, n_11653);
  not g24865 (n_11654, n13593);
  not g24866 (n_11655, n13594);
  and g24867 (n13595, n_11654, n_11655);
  and g24868 (n13596, n_11268, n_11273);
  and g24869 (n13597, n13595, n13596);
  not g24870 (n_11656, n13595);
  not g24871 (n_11657, n13596);
  and g24872 (n13598, n_11656, n_11657);
  not g24873 (n_11658, n13597);
  not g24874 (n_11659, n13598);
  and g24875 (n13599, n_11658, n_11659);
  and g24876 (n13600, \b[27] , n5035);
  and g24877 (n13601, \b[25] , n5277);
  and g24878 (n13602, \b[26] , n5030);
  and g24884 (n13605, n2990, n5038);
  not g24887 (n_11664, n13606);
  and g24888 (n13607, \a[38] , n_11664);
  not g24889 (n_11665, n13607);
  and g24890 (n13608, \a[38] , n_11665);
  and g24891 (n13609, n_11664, n_11665);
  not g24892 (n_11666, n13608);
  not g24893 (n_11667, n13609);
  and g24894 (n13610, n_11666, n_11667);
  not g24895 (n_11668, n13610);
  and g24896 (n13611, n13599, n_11668);
  not g24897 (n_11669, n13611);
  and g24898 (n13612, n13599, n_11669);
  and g24899 (n13613, n_11668, n_11669);
  not g24900 (n_11670, n13612);
  not g24901 (n_11671, n13613);
  and g24902 (n13614, n_11670, n_11671);
  and g24903 (n13615, n_11283, n_11289);
  and g24904 (n13616, n13614, n13615);
  not g24905 (n_11672, n13614);
  not g24906 (n_11673, n13615);
  and g24907 (n13617, n_11672, n_11673);
  not g24908 (n_11674, n13616);
  not g24909 (n_11675, n13617);
  and g24910 (n13618, n_11674, n_11675);
  and g24911 (n13619, \b[30] , n4287);
  and g24912 (n13620, \b[28] , n4532);
  and g24913 (n13621, \b[29] , n4282);
  and g24919 (n13624, n3577, n4290);
  not g24922 (n_11680, n13625);
  and g24923 (n13626, \a[35] , n_11680);
  not g24924 (n_11681, n13626);
  and g24925 (n13627, \a[35] , n_11681);
  and g24926 (n13628, n_11680, n_11681);
  not g24927 (n_11682, n13627);
  not g24928 (n_11683, n13628);
  and g24929 (n13629, n_11682, n_11683);
  not g24930 (n_11684, n13618);
  and g24931 (n13630, n_11684, n13629);
  not g24932 (n_11685, n13629);
  and g24933 (n13631, n13618, n_11685);
  not g24934 (n_11686, n13630);
  not g24935 (n_11687, n13631);
  and g24936 (n13632, n_11686, n_11687);
  and g24937 (n13633, n_11299, n_11305);
  not g24938 (n_11688, n13633);
  and g24939 (n13634, n13632, n_11688);
  not g24940 (n_11689, n13632);
  and g24941 (n13635, n_11689, n13633);
  not g24942 (n_11690, n13634);
  not g24943 (n_11691, n13635);
  and g24944 (n13636, n_11690, n_11691);
  not g24945 (n_11692, n13447);
  and g24946 (n13637, n_11692, n13636);
  not g24947 (n_11693, n13637);
  and g24948 (n13638, n13636, n_11693);
  and g24949 (n13639, n_11692, n_11693);
  not g24950 (n_11694, n13638);
  not g24951 (n_11695, n13639);
  and g24952 (n13640, n_11694, n_11695);
  not g24953 (n_11696, n13207);
  and g24954 (n13641, n_11696, n13640);
  not g24955 (n_11697, n13640);
  and g24956 (n13642, n13207, n_11697);
  not g24957 (n_11698, n13641);
  not g24958 (n_11699, n13642);
  and g24959 (n13643, n_11698, n_11699);
  and g24960 (n13644, \b[36] , n3050);
  and g24961 (n13645, \b[34] , n3243);
  and g24962 (n13646, \b[35] , n3045);
  and g24968 (n13649, n3053, n4922);
  not g24971 (n_11704, n13650);
  and g24972 (n13651, \a[29] , n_11704);
  not g24973 (n_11705, n13651);
  and g24974 (n13652, \a[29] , n_11705);
  and g24975 (n13653, n_11704, n_11705);
  not g24976 (n_11706, n13652);
  not g24977 (n_11707, n13653);
  and g24978 (n13654, n_11706, n_11707);
  not g24979 (n_11708, n13643);
  not g24980 (n_11709, n13654);
  and g24981 (n13655, n_11708, n_11709);
  and g24982 (n13656, n13643, n13654);
  not g24983 (n_11710, n13655);
  not g24984 (n_11711, n13656);
  and g24985 (n13657, n_11710, n_11711);
  not g24986 (n_11712, n13657);
  and g24987 (n13658, n13436, n_11712);
  not g24988 (n_11713, n13436);
  and g24989 (n13659, n_11713, n13657);
  not g24990 (n_11714, n13658);
  not g24991 (n_11715, n13659);
  and g24992 (n13660, n_11714, n_11715);
  and g24993 (n13661, \b[39] , n2539);
  and g24994 (n13662, \b[37] , n2685);
  and g24995 (n13663, \b[38] , n2534);
  and g25001 (n13666, n2542, n5451);
  not g25004 (n_11720, n13667);
  and g25005 (n13668, \a[26] , n_11720);
  not g25006 (n_11721, n13668);
  and g25007 (n13669, \a[26] , n_11721);
  and g25008 (n13670, n_11720, n_11721);
  not g25009 (n_11722, n13669);
  not g25010 (n_11723, n13670);
  and g25011 (n13671, n_11722, n_11723);
  not g25012 (n_11724, n13660);
  and g25013 (n13672, n_11724, n13671);
  not g25014 (n_11725, n13671);
  and g25015 (n13673, n13660, n_11725);
  not g25016 (n_11726, n13672);
  not g25017 (n_11727, n13673);
  and g25018 (n13674, n_11726, n_11727);
  not g25019 (n_11728, n13435);
  and g25020 (n13675, n_11728, n13674);
  not g25021 (n_11729, n13674);
  and g25022 (n13676, n13435, n_11729);
  not g25023 (n_11730, n13675);
  not g25024 (n_11731, n13676);
  and g25025 (n13677, n_11730, n_11731);
  not g25026 (n_11732, n13434);
  and g25027 (n13678, n_11732, n13677);
  not g25028 (n_11733, n13678);
  and g25029 (n13679, n_11732, n_11733);
  and g25030 (n13680, n13677, n_11733);
  not g25031 (n_11734, n13679);
  not g25032 (n_11735, n13680);
  and g25033 (n13681, n_11734, n_11735);
  not g25034 (n_11736, n13264);
  not g25035 (n_11737, n13681);
  and g25036 (n13682, n_11736, n_11737);
  and g25037 (n13683, n13264, n_11735);
  and g25038 (n13684, n_11734, n13683);
  not g25039 (n_11738, n13682);
  not g25040 (n_11739, n13684);
  and g25041 (n13685, n_11738, n_11739);
  not g25042 (n_11740, n13423);
  and g25043 (n13686, n_11740, n13685);
  not g25044 (n_11741, n13686);
  and g25045 (n13687, n_11740, n_11741);
  and g25046 (n13688, n13685, n_11741);
  not g25047 (n_11742, n13687);
  not g25048 (n_11743, n13688);
  and g25049 (n13689, n_11742, n_11743);
  not g25050 (n_11744, n13412);
  not g25051 (n_11745, n13689);
  and g25052 (n13690, n_11744, n_11745);
  and g25053 (n13691, n13412, n_11743);
  and g25054 (n13692, n_11742, n13691);
  not g25055 (n_11746, n13690);
  not g25056 (n_11747, n13692);
  and g25057 (n13693, n_11746, n_11747);
  not g25058 (n_11748, n13410);
  and g25059 (n13694, n_11748, n13693);
  not g25060 (n_11749, n13694);
  and g25061 (n13695, n_11748, n_11749);
  and g25062 (n13696, n13693, n_11749);
  not g25063 (n_11750, n13695);
  not g25064 (n_11751, n13696);
  and g25065 (n13697, n_11750, n_11751);
  not g25066 (n_11752, n13399);
  not g25067 (n_11753, n13697);
  and g25068 (n13698, n_11752, n_11753);
  and g25069 (n13699, n13399, n_11751);
  and g25070 (n13700, n_11750, n13699);
  not g25071 (n_11754, n13698);
  not g25072 (n_11755, n13700);
  and g25073 (n13701, n_11754, n_11755);
  not g25074 (n_11756, n13398);
  and g25075 (n13702, n_11756, n13701);
  not g25076 (n_11757, n13701);
  and g25077 (n13703, n13398, n_11757);
  not g25078 (n_11758, n13702);
  not g25079 (n_11759, n13703);
  and g25080 (n13704, n_11758, n_11759);
  not g25081 (n_11760, n13387);
  and g25082 (n13705, n_11760, n13704);
  not g25083 (n_11761, n13704);
  and g25084 (n13706, n13387, n_11761);
  not g25085 (n_11762, n13705);
  not g25086 (n_11763, n13706);
  and g25087 (n13707, n_11762, n_11763);
  and g25088 (n13708, \b[54] , n700);
  and g25089 (n13709, \b[52] , n767);
  and g25090 (n13710, \b[53] , n695);
  and g25096 (n13713, n703, n9998);
  not g25099 (n_11768, n13714);
  and g25100 (n13715, \a[11] , n_11768);
  not g25101 (n_11769, n13715);
  and g25102 (n13716, \a[11] , n_11769);
  and g25103 (n13717, n_11768, n_11769);
  not g25104 (n_11770, n13716);
  not g25105 (n_11771, n13717);
  and g25106 (n13718, n_11770, n_11771);
  not g25107 (n_11772, n13718);
  and g25108 (n13719, n13707, n_11772);
  not g25109 (n_11773, n13719);
  and g25110 (n13720, n13707, n_11773);
  and g25111 (n13721, n_11772, n_11773);
  not g25112 (n_11774, n13720);
  not g25113 (n_11775, n13721);
  and g25114 (n13722, n_11774, n_11775);
  and g25115 (n13723, n_11422, n_11426);
  and g25116 (n13724, n13722, n13723);
  not g25117 (n_11776, n13722);
  not g25118 (n_11777, n13723);
  and g25119 (n13725, n_11776, n_11777);
  not g25120 (n_11778, n13724);
  not g25121 (n_11779, n13725);
  and g25122 (n13726, n_11778, n_11779);
  and g25123 (n13727, \b[57] , n511);
  and g25124 (n13728, \b[55] , n541);
  and g25125 (n13729, \b[56] , n506);
  and g25131 (n13732, n514, n11410);
  not g25134 (n_11784, n13733);
  and g25135 (n13734, \a[8] , n_11784);
  not g25136 (n_11785, n13734);
  and g25137 (n13735, \a[8] , n_11785);
  and g25138 (n13736, n_11784, n_11785);
  not g25139 (n_11786, n13735);
  not g25140 (n_11787, n13736);
  and g25141 (n13737, n_11786, n_11787);
  not g25142 (n_11788, n13737);
  and g25143 (n13738, n13726, n_11788);
  not g25144 (n_11789, n13738);
  and g25145 (n13739, n13726, n_11789);
  and g25146 (n13740, n_11788, n_11789);
  not g25147 (n_11790, n13739);
  not g25148 (n_11791, n13740);
  and g25149 (n13741, n_11790, n_11791);
  and g25150 (n13742, \b[60] , n362);
  and g25151 (n13743, \b[58] , n403);
  and g25152 (n13744, \b[59] , n357);
  and g25158 (n13747, n365, n12211);
  not g25161 (n_11796, n13748);
  and g25162 (n13749, \a[5] , n_11796);
  not g25163 (n_11797, n13749);
  and g25164 (n13750, \a[5] , n_11797);
  and g25165 (n13751, n_11796, n_11797);
  not g25166 (n_11798, n13750);
  not g25167 (n_11799, n13751);
  and g25168 (n13752, n_11798, n_11799);
  not g25169 (n_11800, n13741);
  and g25170 (n13753, n_11800, n13752);
  not g25171 (n_11801, n13752);
  and g25172 (n13754, n13741, n_11801);
  not g25173 (n_11802, n13753);
  not g25174 (n_11803, n13754);
  and g25175 (n13755, n_11802, n_11803);
  and g25176 (n13756, n_11439, n_11449);
  and g25177 (n13757, n13755, n13756);
  not g25178 (n_11804, n13755);
  not g25179 (n_11805, n13756);
  and g25180 (n13758, n_11804, n_11805);
  not g25181 (n_11806, n13757);
  not g25182 (n_11807, n13758);
  and g25183 (n13759, n_11806, n_11807);
  and g25184 (n13760, \b[63] , n266);
  and g25185 (n13761, \b[61] , n284);
  and g25186 (n13762, \b[62] , n261);
  and g25192 (n13765, n_11462, n_11465);
  not g25193 (n_11812, \b[63] );
  and g25194 (n13766, \b[62] , n_11812);
  and g25195 (n13767, n_11460, \b[63] );
  not g25196 (n_11813, n13766);
  not g25197 (n_11814, n13767);
  and g25198 (n13768, n_11813, n_11814);
  not g25199 (n_11815, n13765);
  not g25200 (n_11816, n13768);
  and g25201 (n13769, n_11815, n_11816);
  and g25202 (n13770, n13765, n13768);
  not g25203 (n_11817, n13769);
  not g25204 (n_11818, n13770);
  and g25205 (n13771, n_11817, n_11818);
  and g25206 (n13772, n269, n13771);
  not g25209 (n_11820, n13773);
  and g25210 (n13774, \a[2] , n_11820);
  not g25211 (n_11821, n13774);
  and g25212 (n13775, \a[2] , n_11821);
  and g25213 (n13776, n_11820, n_11821);
  not g25214 (n_11822, n13775);
  not g25215 (n_11823, n13776);
  and g25216 (n13777, n_11822, n_11823);
  not g25217 (n_11824, n13777);
  and g25218 (n13778, n13759, n_11824);
  not g25219 (n_11825, n13778);
  and g25220 (n13779, n13759, n_11825);
  and g25221 (n13780, n_11824, n_11825);
  not g25222 (n_11826, n13779);
  not g25223 (n_11827, n13780);
  and g25224 (n13781, n_11826, n_11827);
  and g25225 (n13782, n_11455, n_11475);
  not g25226 (n_11828, n13781);
  not g25227 (n_11829, n13782);
  and g25228 (n13783, n_11828, n_11829);
  not g25229 (n_11830, n13783);
  and g25230 (n13784, n_11828, n_11830);
  and g25231 (n13785, n_11829, n_11830);
  not g25232 (n_11831, n13784);
  not g25233 (n_11832, n13785);
  and g25234 (n13786, n_11831, n_11832);
  and g25235 (n13787, n_11478, n_11482);
  not g25236 (n_11833, n13786);
  not g25237 (n_11834, n13787);
  and g25238 (n13788, n_11833, n_11834);
  and g25239 (n13789, n13786, n13787);
  not g25240 (n_11835, n13788);
  not g25241 (n_11836, n13789);
  and g25242 (\f[63] , n_11835, n_11836);
  and g25243 (n13791, n_11830, n_11835);
  and g25244 (n13792, n_11807, n_11825);
  and g25245 (n13793, \b[62] , n284);
  and g25246 (n13794, \b[63] , n261);
  not g25247 (n_11837, n13793);
  not g25248 (n_11838, n13794);
  and g25249 (n13795, n_11837, n_11838);
  and g25250 (n13796, n_11460, n_11817);
  not g25251 (n_11839, n13796);
  and g25252 (n13797, \b[63] , n_11839);
  not g25253 (n_11840, n13797);
  and g25254 (n13798, \b[63] , n_11840);
  and g25255 (n13799, n_11815, n13766);
  not g25256 (n_11841, n13798);
  not g25257 (n_11842, n13799);
  and g25258 (n13800, n_11841, n_11842);
  not g25259 (n_11843, n13800);
  and g25260 (n13801, n269, n_11843);
  not g25261 (n_11844, n13801);
  and g25262 (n13802, n13795, n_11844);
  not g25263 (n_11845, n13802);
  and g25264 (n13803, \a[2] , n_11845);
  not g25265 (n_11846, n13803);
  and g25266 (n13804, \a[2] , n_11846);
  and g25267 (n13805, n_11845, n_11846);
  not g25268 (n_11847, n13804);
  not g25269 (n_11848, n13805);
  and g25270 (n13806, n_11847, n_11848);
  and g25271 (n13807, n_11800, n_11801);
  not g25272 (n_11849, n13807);
  and g25273 (n13808, n_11789, n_11849);
  and g25274 (n13809, n_11773, n_11779);
  and g25275 (n13810, \b[55] , n700);
  and g25276 (n13811, \b[53] , n767);
  and g25277 (n13812, \b[54] , n695);
  and g25283 (n13815, n703, n10684);
  not g25286 (n_11854, n13816);
  and g25287 (n13817, \a[11] , n_11854);
  not g25288 (n_11855, n13817);
  and g25289 (n13818, \a[11] , n_11855);
  and g25290 (n13819, n_11854, n_11855);
  not g25291 (n_11856, n13818);
  not g25292 (n_11857, n13819);
  and g25293 (n13820, n_11856, n_11857);
  and g25294 (n13821, n_11758, n_11762);
  and g25295 (n13822, \b[52] , n951);
  and g25296 (n13823, \b[50] , n1056);
  and g25297 (n13824, \b[51] , n946);
  and g25303 (n13827, n954, n9628);
  not g25306 (n_11862, n13828);
  and g25307 (n13829, \a[14] , n_11862);
  not g25308 (n_11863, n13829);
  and g25309 (n13830, \a[14] , n_11863);
  and g25310 (n13831, n_11862, n_11863);
  not g25311 (n_11864, n13830);
  not g25312 (n_11865, n13831);
  and g25313 (n13832, n_11864, n_11865);
  and g25314 (n13833, n_11749, n_11754);
  and g25315 (n13834, \b[49] , n1302);
  and g25316 (n13835, \b[47] , n1391);
  and g25317 (n13836, \b[48] , n1297);
  and g25323 (n13839, n1305, n8625);
  not g25326 (n_11870, n13840);
  and g25327 (n13841, \a[17] , n_11870);
  not g25328 (n_11871, n13841);
  and g25329 (n13842, \a[17] , n_11871);
  and g25330 (n13843, n_11870, n_11871);
  not g25331 (n_11872, n13842);
  not g25332 (n_11873, n13843);
  and g25333 (n13844, n_11872, n_11873);
  and g25334 (n13845, n_11741, n_11746);
  and g25335 (n13846, \b[46] , n1627);
  and g25336 (n13847, \b[44] , n1763);
  and g25337 (n13848, \b[45] , n1622);
  and g25343 (n13851, n1630, n7677);
  not g25346 (n_11878, n13852);
  and g25347 (n13853, \a[20] , n_11878);
  not g25348 (n_11879, n13853);
  and g25349 (n13854, \a[20] , n_11879);
  and g25350 (n13855, n_11878, n_11879);
  not g25351 (n_11880, n13854);
  not g25352 (n_11881, n13855);
  and g25353 (n13856, n_11880, n_11881);
  and g25354 (n13857, n_11733, n_11738);
  and g25355 (n13858, \b[34] , n3638);
  and g25356 (n13859, \b[32] , n3843);
  and g25357 (n13860, \b[33] , n3633);
  and g25363 (n13863, n3641, n4466);
  not g25366 (n_11886, n13864);
  and g25367 (n13865, \a[32] , n_11886);
  not g25368 (n_11887, n13865);
  and g25369 (n13866, \a[32] , n_11887);
  and g25370 (n13867, n_11886, n_11887);
  not g25371 (n_11888, n13866);
  not g25372 (n_11889, n13867);
  and g25373 (n13868, n_11888, n_11889);
  and g25374 (n13869, \b[22] , n6595);
  and g25375 (n13870, \b[20] , n6902);
  and g25376 (n13871, \b[21] , n6590);
  and g25382 (n13874, n2145, n6598);
  not g25385 (n_11894, n13875);
  and g25386 (n13876, \a[44] , n_11894);
  not g25387 (n_11895, n13876);
  and g25388 (n13877, \a[44] , n_11895);
  and g25389 (n13878, n_11894, n_11895);
  not g25390 (n_11896, n13877);
  not g25391 (n_11897, n13878);
  and g25392 (n13879, n_11896, n_11897);
  and g25393 (n13880, \b[16] , n8362);
  and g25394 (n13881, \b[14] , n8715);
  and g25395 (n13882, \b[15] , n8357);
  and g25401 (n13885, n1237, n8365);
  not g25404 (n_11902, n13886);
  and g25405 (n13887, \a[50] , n_11902);
  not g25406 (n_11903, n13887);
  and g25407 (n13888, \a[50] , n_11903);
  and g25408 (n13889, n_11902, n_11903);
  not g25409 (n_11904, n13888);
  not g25410 (n_11905, n13889);
  and g25411 (n13890, n_11904, n_11905);
  and g25412 (n13891, \b[10] , n10426);
  and g25413 (n13892, \b[8] , n10796);
  and g25414 (n13893, \b[9] , n10421);
  and g25420 (n13896, n738, n10429);
  not g25423 (n_11910, n13897);
  and g25424 (n13898, \a[56] , n_11910);
  not g25425 (n_11911, n13898);
  and g25426 (n13899, \a[56] , n_11911);
  and g25427 (n13900, n_11910, n_11911);
  not g25428 (n_11912, n13899);
  not g25429 (n_11913, n13900);
  and g25430 (n13901, n_11912, n_11913);
  and g25431 (n13902, n_11583, n_11586);
  and g25432 (n13903, \a[63] , n13488);
  and g25433 (n13904, \b[0] , n13903);
  and g25434 (n13905, \b[1] , n_11555);
  not g25435 (n_11914, n13904);
  not g25436 (n_11915, n13905);
  and g25437 (n13906, n_11914, n_11915);
  and g25438 (n13907, \b[4] , n12668);
  and g25439 (n13908, \b[2] , n13047);
  and g25440 (n13909, \b[3] , n12663);
  and g25446 (n13912, n346, n12671);
  not g25449 (n_11920, n13913);
  and g25450 (n13914, \a[62] , n_11920);
  not g25451 (n_11921, n13914);
  and g25452 (n13915, \a[62] , n_11921);
  and g25453 (n13916, n_11920, n_11921);
  not g25454 (n_11922, n13915);
  not g25455 (n_11923, n13916);
  and g25456 (n13917, n_11922, n_11923);
  not g25457 (n_11924, n13906);
  not g25458 (n_11925, n13917);
  and g25459 (n13918, n_11924, n_11925);
  not g25460 (n_11926, n13918);
  and g25461 (n13919, n_11924, n_11926);
  and g25462 (n13920, n_11925, n_11926);
  not g25463 (n_11927, n13919);
  not g25464 (n_11928, n13920);
  and g25465 (n13921, n_11927, n_11928);
  and g25466 (n13922, n_11556, n_11569);
  and g25467 (n13923, n13921, n13922);
  not g25468 (n_11929, n13921);
  not g25469 (n_11930, n13922);
  and g25470 (n13924, n_11929, n_11930);
  not g25471 (n_11931, n13923);
  not g25472 (n_11932, n13924);
  and g25473 (n13925, n_11931, n_11932);
  and g25474 (n13926, \b[7] , n11531);
  and g25475 (n13927, \b[5] , n11896);
  and g25476 (n13928, \b[6] , n11526);
  and g25482 (n13931, n484, n11534);
  not g25485 (n_11937, n13932);
  and g25486 (n13933, \a[59] , n_11937);
  not g25487 (n_11938, n13933);
  and g25488 (n13934, \a[59] , n_11938);
  and g25489 (n13935, n_11937, n_11938);
  not g25490 (n_11939, n13934);
  not g25491 (n_11940, n13935);
  and g25492 (n13936, n_11939, n_11940);
  not g25493 (n_11941, n13925);
  and g25494 (n13937, n_11941, n13936);
  not g25495 (n_11942, n13936);
  and g25496 (n13938, n13925, n_11942);
  not g25497 (n_11943, n13937);
  not g25498 (n_11944, n13938);
  and g25499 (n13939, n_11943, n_11944);
  not g25500 (n_11945, n13902);
  and g25501 (n13940, n_11945, n13939);
  not g25502 (n_11946, n13939);
  and g25503 (n13941, n13902, n_11946);
  not g25504 (n_11947, n13940);
  not g25505 (n_11948, n13941);
  and g25506 (n13942, n_11947, n_11948);
  not g25507 (n_11949, n13901);
  and g25508 (n13943, n_11949, n13942);
  not g25509 (n_11950, n13943);
  and g25510 (n13944, n13942, n_11950);
  and g25511 (n13945, n_11949, n_11950);
  not g25512 (n_11951, n13944);
  not g25513 (n_11952, n13945);
  and g25514 (n13946, n_11951, n_11952);
  and g25515 (n13947, n_11592, n_11593);
  not g25516 (n_11953, n13947);
  and g25517 (n13948, n_11589, n_11953);
  and g25518 (n13949, n13946, n13948);
  not g25519 (n_11954, n13946);
  not g25520 (n_11955, n13948);
  and g25521 (n13950, n_11954, n_11955);
  not g25522 (n_11956, n13949);
  not g25523 (n_11957, n13950);
  and g25524 (n13951, n_11956, n_11957);
  and g25525 (n13952, \b[13] , n9339);
  and g25526 (n13953, \b[11] , n9732);
  and g25527 (n13954, \b[12] , n9334);
  and g25533 (n13957, n1008, n9342);
  not g25536 (n_11962, n13958);
  and g25537 (n13959, \a[53] , n_11962);
  not g25538 (n_11963, n13959);
  and g25539 (n13960, \a[53] , n_11963);
  and g25540 (n13961, n_11962, n_11963);
  not g25541 (n_11964, n13960);
  not g25542 (n_11965, n13961);
  and g25543 (n13962, n_11964, n_11965);
  not g25544 (n_11966, n13951);
  and g25545 (n13963, n_11966, n13962);
  not g25546 (n_11967, n13962);
  and g25547 (n13964, n13951, n_11967);
  not g25548 (n_11968, n13963);
  not g25549 (n_11969, n13964);
  and g25550 (n13965, n_11968, n_11969);
  and g25551 (n13966, n_11607, n_11610);
  not g25552 (n_11970, n13966);
  and g25553 (n13967, n13965, n_11970);
  not g25554 (n_11971, n13965);
  and g25555 (n13968, n_11971, n13966);
  not g25556 (n_11972, n13967);
  not g25557 (n_11973, n13968);
  and g25558 (n13969, n_11972, n_11973);
  not g25559 (n_11974, n13890);
  and g25560 (n13970, n_11974, n13969);
  not g25561 (n_11975, n13970);
  and g25562 (n13971, n13969, n_11975);
  and g25563 (n13972, n_11974, n_11975);
  not g25564 (n_11976, n13971);
  not g25565 (n_11977, n13972);
  and g25566 (n13973, n_11976, n_11977);
  and g25567 (n13974, n_11613, n_11619);
  and g25568 (n13975, n13973, n13974);
  not g25569 (n_11978, n13973);
  not g25570 (n_11979, n13974);
  and g25571 (n13976, n_11978, n_11979);
  not g25572 (n_11980, n13975);
  not g25573 (n_11981, n13976);
  and g25574 (n13977, n_11980, n_11981);
  and g25575 (n13978, \b[19] , n7446);
  and g25576 (n13979, \b[17] , n7787);
  and g25577 (n13980, \b[18] , n7441);
  and g25583 (n13983, n1708, n7449);
  not g25586 (n_11986, n13984);
  and g25587 (n13985, \a[47] , n_11986);
  not g25588 (n_11987, n13985);
  and g25589 (n13986, \a[47] , n_11987);
  and g25590 (n13987, n_11986, n_11987);
  not g25591 (n_11988, n13986);
  not g25592 (n_11989, n13987);
  and g25593 (n13988, n_11988, n_11989);
  not g25594 (n_11990, n13977);
  and g25595 (n13989, n_11990, n13988);
  not g25596 (n_11991, n13988);
  and g25597 (n13990, n13977, n_11991);
  not g25598 (n_11992, n13989);
  not g25599 (n_11993, n13990);
  and g25600 (n13991, n_11992, n_11993);
  and g25601 (n13992, n_11631, n_11634);
  not g25602 (n_11994, n13992);
  and g25603 (n13993, n13991, n_11994);
  not g25604 (n_11995, n13991);
  and g25605 (n13994, n_11995, n13992);
  not g25606 (n_11996, n13993);
  not g25607 (n_11997, n13994);
  and g25608 (n13995, n_11996, n_11997);
  not g25609 (n_11998, n13879);
  and g25610 (n13996, n_11998, n13995);
  not g25611 (n_11999, n13996);
  and g25612 (n13997, n13995, n_11999);
  and g25613 (n13998, n_11998, n_11999);
  not g25614 (n_12000, n13997);
  not g25615 (n_12001, n13998);
  and g25616 (n13999, n_12000, n_12001);
  and g25617 (n14000, n_11638, n_11642);
  and g25618 (n14001, n13999, n14000);
  not g25619 (n_12002, n13999);
  not g25620 (n_12003, n14000);
  and g25621 (n14002, n_12002, n_12003);
  not g25622 (n_12004, n14001);
  not g25623 (n_12005, n14002);
  and g25624 (n14003, n_12004, n_12005);
  and g25625 (n14004, \b[25] , n5777);
  and g25626 (n14005, \b[23] , n6059);
  and g25627 (n14006, \b[24] , n5772);
  and g25633 (n14009, n2485, n5780);
  not g25636 (n_12010, n14010);
  and g25637 (n14011, \a[41] , n_12010);
  not g25638 (n_12011, n14011);
  and g25639 (n14012, \a[41] , n_12011);
  and g25640 (n14013, n_12010, n_12011);
  not g25641 (n_12012, n14012);
  not g25642 (n_12013, n14013);
  and g25643 (n14014, n_12012, n_12013);
  not g25644 (n_12014, n14014);
  and g25645 (n14015, n14003, n_12014);
  not g25646 (n_12015, n14015);
  and g25647 (n14016, n14003, n_12015);
  and g25648 (n14017, n_12014, n_12015);
  not g25649 (n_12016, n14016);
  not g25650 (n_12017, n14017);
  and g25651 (n14018, n_12016, n_12017);
  and g25652 (n14019, n_11653, n_11659);
  and g25653 (n14020, n14018, n14019);
  not g25654 (n_12018, n14018);
  not g25655 (n_12019, n14019);
  and g25656 (n14021, n_12018, n_12019);
  not g25657 (n_12020, n14020);
  not g25658 (n_12021, n14021);
  and g25659 (n14022, n_12020, n_12021);
  and g25660 (n14023, \b[28] , n5035);
  and g25661 (n14024, \b[26] , n5277);
  and g25662 (n14025, \b[27] , n5030);
  and g25668 (n14028, n3189, n5038);
  not g25671 (n_12026, n14029);
  and g25672 (n14030, \a[38] , n_12026);
  not g25673 (n_12027, n14030);
  and g25674 (n14031, \a[38] , n_12027);
  and g25675 (n14032, n_12026, n_12027);
  not g25676 (n_12028, n14031);
  not g25677 (n_12029, n14032);
  and g25678 (n14033, n_12028, n_12029);
  not g25679 (n_12030, n14033);
  and g25680 (n14034, n14022, n_12030);
  not g25681 (n_12031, n14034);
  and g25682 (n14035, n14022, n_12031);
  and g25683 (n14036, n_12030, n_12031);
  not g25684 (n_12032, n14035);
  not g25685 (n_12033, n14036);
  and g25686 (n14037, n_12032, n_12033);
  and g25687 (n14038, n_11669, n_11675);
  and g25688 (n14039, n14037, n14038);
  not g25689 (n_12034, n14037);
  not g25690 (n_12035, n14038);
  and g25691 (n14040, n_12034, n_12035);
  not g25692 (n_12036, n14039);
  not g25693 (n_12037, n14040);
  and g25694 (n14041, n_12036, n_12037);
  and g25695 (n14042, \b[31] , n4287);
  and g25696 (n14043, \b[29] , n4532);
  and g25697 (n14044, \b[30] , n4282);
  and g25703 (n14047, n3796, n4290);
  not g25706 (n_12042, n14048);
  and g25707 (n14049, \a[35] , n_12042);
  not g25708 (n_12043, n14049);
  and g25709 (n14050, \a[35] , n_12043);
  and g25710 (n14051, n_12042, n_12043);
  not g25711 (n_12044, n14050);
  not g25712 (n_12045, n14051);
  and g25713 (n14052, n_12044, n_12045);
  not g25714 (n_12046, n14041);
  and g25715 (n14053, n_12046, n14052);
  not g25716 (n_12047, n14052);
  and g25717 (n14054, n14041, n_12047);
  not g25718 (n_12048, n14053);
  not g25719 (n_12049, n14054);
  and g25720 (n14055, n_12048, n_12049);
  and g25721 (n14056, n_11687, n_11690);
  not g25722 (n_12050, n14056);
  and g25723 (n14057, n14055, n_12050);
  not g25724 (n_12051, n14055);
  and g25725 (n14058, n_12051, n14056);
  not g25726 (n_12052, n14057);
  not g25727 (n_12053, n14058);
  and g25728 (n14059, n_12052, n_12053);
  not g25729 (n_12054, n13868);
  and g25730 (n14060, n_12054, n14059);
  not g25731 (n_12055, n14060);
  and g25732 (n14061, n14059, n_12055);
  and g25733 (n14062, n_12054, n_12055);
  not g25734 (n_12056, n14061);
  not g25735 (n_12057, n14062);
  and g25736 (n14063, n_12056, n_12057);
  and g25737 (n14064, n_11696, n_11697);
  not g25738 (n_12058, n14064);
  and g25739 (n14065, n_11693, n_12058);
  and g25740 (n14066, n14063, n14065);
  not g25741 (n_12059, n14063);
  not g25742 (n_12060, n14065);
  and g25743 (n14067, n_12059, n_12060);
  not g25744 (n_12061, n14066);
  not g25745 (n_12062, n14067);
  and g25746 (n14068, n_12061, n_12062);
  and g25747 (n14069, \b[37] , n3050);
  and g25748 (n14070, \b[35] , n3243);
  and g25749 (n14071, \b[36] , n3045);
  and g25755 (n14074, n3053, n5181);
  not g25758 (n_12067, n14075);
  and g25759 (n14076, \a[29] , n_12067);
  not g25760 (n_12068, n14076);
  and g25761 (n14077, \a[29] , n_12068);
  and g25762 (n14078, n_12067, n_12068);
  not g25763 (n_12069, n14077);
  not g25764 (n_12070, n14078);
  and g25765 (n14079, n_12069, n_12070);
  not g25766 (n_12071, n14079);
  and g25767 (n14080, n14068, n_12071);
  not g25768 (n_12072, n14080);
  and g25769 (n14081, n14068, n_12072);
  and g25770 (n14082, n_12071, n_12072);
  not g25771 (n_12073, n14081);
  not g25772 (n_12074, n14082);
  and g25773 (n14083, n_12073, n_12074);
  and g25774 (n14084, n_11710, n_11715);
  and g25775 (n14085, n14083, n14084);
  not g25776 (n_12075, n14083);
  not g25777 (n_12076, n14084);
  and g25778 (n14086, n_12075, n_12076);
  not g25779 (n_12077, n14085);
  not g25780 (n_12078, n14086);
  and g25781 (n14087, n_12077, n_12078);
  and g25782 (n14088, \b[40] , n2539);
  and g25783 (n14089, \b[38] , n2685);
  and g25784 (n14090, \b[39] , n2534);
  and g25790 (n14093, n2542, n5955);
  not g25793 (n_12083, n14094);
  and g25794 (n14095, \a[26] , n_12083);
  not g25795 (n_12084, n14095);
  and g25796 (n14096, \a[26] , n_12084);
  and g25797 (n14097, n_12083, n_12084);
  not g25798 (n_12085, n14096);
  not g25799 (n_12086, n14097);
  and g25800 (n14098, n_12085, n_12086);
  not g25801 (n_12087, n14098);
  and g25802 (n14099, n14087, n_12087);
  not g25803 (n_12088, n14099);
  and g25804 (n14100, n14087, n_12088);
  and g25805 (n14101, n_12087, n_12088);
  not g25806 (n_12089, n14100);
  not g25807 (n_12090, n14101);
  and g25808 (n14102, n_12089, n_12090);
  and g25809 (n14103, n_11727, n_11730);
  not g25810 (n_12091, n14102);
  not g25811 (n_12092, n14103);
  and g25812 (n14104, n_12091, n_12092);
  not g25813 (n_12093, n14104);
  and g25814 (n14105, n_12091, n_12093);
  and g25815 (n14106, n_12092, n_12093);
  not g25816 (n_12094, n14105);
  not g25817 (n_12095, n14106);
  and g25818 (n14107, n_12094, n_12095);
  and g25819 (n14108, \b[43] , n2048);
  and g25820 (n14109, \b[41] , n2198);
  and g25821 (n14110, \b[42] , n2043);
  and g25827 (n14113, n2051, n6515);
  not g25830 (n_12100, n14114);
  and g25831 (n14115, \a[23] , n_12100);
  not g25832 (n_12101, n14115);
  and g25833 (n14116, \a[23] , n_12101);
  and g25834 (n14117, n_12100, n_12101);
  not g25835 (n_12102, n14116);
  not g25836 (n_12103, n14117);
  and g25837 (n14118, n_12102, n_12103);
  not g25838 (n_12104, n14107);
  and g25839 (n14119, n_12104, n14118);
  not g25840 (n_12105, n14118);
  and g25841 (n14120, n14107, n_12105);
  not g25842 (n_12106, n14119);
  not g25843 (n_12107, n14120);
  and g25844 (n14121, n_12106, n_12107);
  not g25845 (n_12108, n13857);
  not g25846 (n_12109, n14121);
  and g25847 (n14122, n_12108, n_12109);
  and g25848 (n14123, n13857, n14121);
  not g25849 (n_12110, n14122);
  not g25850 (n_12111, n14123);
  and g25851 (n14124, n_12110, n_12111);
  not g25852 (n_12112, n13856);
  and g25853 (n14125, n_12112, n14124);
  not g25854 (n_12113, n14125);
  and g25855 (n14126, n_12112, n_12113);
  and g25856 (n14127, n14124, n_12113);
  not g25857 (n_12114, n14126);
  not g25858 (n_12115, n14127);
  and g25859 (n14128, n_12114, n_12115);
  not g25860 (n_12116, n13845);
  not g25861 (n_12117, n14128);
  and g25862 (n14129, n_12116, n_12117);
  and g25863 (n14130, n13845, n_12115);
  and g25864 (n14131, n_12114, n14130);
  not g25865 (n_12118, n14129);
  not g25866 (n_12119, n14131);
  and g25867 (n14132, n_12118, n_12119);
  not g25868 (n_12120, n13844);
  and g25869 (n14133, n_12120, n14132);
  not g25870 (n_12121, n14133);
  and g25871 (n14134, n_12120, n_12121);
  and g25872 (n14135, n14132, n_12121);
  not g25873 (n_12122, n14134);
  not g25874 (n_12123, n14135);
  and g25875 (n14136, n_12122, n_12123);
  not g25876 (n_12124, n13833);
  not g25877 (n_12125, n14136);
  and g25878 (n14137, n_12124, n_12125);
  and g25879 (n14138, n13833, n_12123);
  and g25880 (n14139, n_12122, n14138);
  not g25881 (n_12126, n14137);
  not g25882 (n_12127, n14139);
  and g25883 (n14140, n_12126, n_12127);
  not g25884 (n_12128, n13832);
  and g25885 (n14141, n_12128, n14140);
  not g25886 (n_12129, n14140);
  and g25887 (n14142, n13832, n_12129);
  not g25888 (n_12130, n14141);
  not g25889 (n_12131, n14142);
  and g25890 (n14143, n_12130, n_12131);
  not g25891 (n_12132, n13821);
  and g25892 (n14144, n_12132, n14143);
  not g25893 (n_12133, n14143);
  and g25894 (n14145, n13821, n_12133);
  not g25895 (n_12134, n14144);
  not g25896 (n_12135, n14145);
  and g25897 (n14146, n_12134, n_12135);
  not g25898 (n_12136, n13820);
  and g25899 (n14147, n_12136, n14146);
  not g25900 (n_12137, n14146);
  and g25901 (n14148, n13820, n_12137);
  not g25902 (n_12138, n14147);
  not g25903 (n_12139, n14148);
  and g25904 (n14149, n_12138, n_12139);
  not g25905 (n_12140, n13809);
  and g25906 (n14150, n_12140, n14149);
  not g25907 (n_12141, n14149);
  and g25908 (n14151, n13809, n_12141);
  not g25909 (n_12142, n14150);
  not g25910 (n_12143, n14151);
  and g25911 (n14152, n_12142, n_12143);
  and g25912 (n14153, \b[58] , n511);
  and g25913 (n14154, \b[56] , n541);
  and g25914 (n14155, \b[57] , n506);
  and g25920 (n14158, n514, n11436);
  not g25923 (n_12148, n14159);
  and g25924 (n14160, \a[8] , n_12148);
  not g25925 (n_12149, n14160);
  and g25926 (n14161, \a[8] , n_12149);
  and g25927 (n14162, n_12148, n_12149);
  not g25928 (n_12150, n14161);
  not g25929 (n_12151, n14162);
  and g25930 (n14163, n_12150, n_12151);
  not g25931 (n_12152, n14163);
  and g25932 (n14164, n14152, n_12152);
  not g25933 (n_12153, n14164);
  and g25934 (n14165, n14152, n_12153);
  and g25935 (n14166, n_12152, n_12153);
  not g25936 (n_12154, n14165);
  not g25937 (n_12155, n14166);
  and g25938 (n14167, n_12154, n_12155);
  and g25939 (n14168, \b[61] , n362);
  and g25940 (n14169, \b[59] , n403);
  and g25941 (n14170, \b[60] , n357);
  and g25947 (n14173, n365, n12969);
  not g25950 (n_12160, n14174);
  and g25951 (n14175, \a[5] , n_12160);
  not g25952 (n_12161, n14175);
  and g25953 (n14176, \a[5] , n_12161);
  and g25954 (n14177, n_12160, n_12161);
  not g25955 (n_12162, n14176);
  not g25956 (n_12163, n14177);
  and g25957 (n14178, n_12162, n_12163);
  not g25958 (n_12164, n14167);
  and g25959 (n14179, n_12164, n14178);
  not g25960 (n_12165, n14178);
  and g25961 (n14180, n14167, n_12165);
  not g25962 (n_12166, n14179);
  not g25963 (n_12167, n14180);
  and g25964 (n14181, n_12166, n_12167);
  not g25965 (n_12168, n13808);
  not g25966 (n_12169, n14181);
  and g25967 (n14182, n_12168, n_12169);
  and g25968 (n14183, n13808, n14181);
  not g25969 (n_12170, n14182);
  not g25970 (n_12171, n14183);
  and g25971 (n14184, n_12170, n_12171);
  not g25972 (n_12172, n13806);
  and g25973 (n14185, n_12172, n14184);
  not g25974 (n_12173, n14184);
  and g25975 (n14186, n13806, n_12173);
  not g25976 (n_12174, n14185);
  not g25977 (n_12175, n14186);
  and g25978 (n14187, n_12174, n_12175);
  not g25979 (n_12176, n13792);
  and g25980 (n14188, n_12176, n14187);
  not g25981 (n_12177, n14187);
  and g25982 (n14189, n13792, n_12177);
  not g25983 (n_12178, n14188);
  not g25984 (n_12179, n14189);
  and g25985 (n14190, n_12178, n_12179);
  not g25986 (n_12180, n13791);
  and g25987 (n14191, n_12180, n14190);
  not g25988 (n_12181, n14190);
  and g25989 (n14192, n13791, n_12181);
  not g25990 (n_12182, n14191);
  not g25991 (n_12183, n14192);
  and g25992 (\f[64] , n_12182, n_12183);
  and g25993 (n14194, \b[53] , n951);
  and g25994 (n14195, \b[51] , n1056);
  and g25995 (n14196, \b[52] , n946);
  and g26001 (n14199, n954, n9972);
  not g26004 (n_12188, n14200);
  and g26005 (n14201, \a[14] , n_12188);
  not g26006 (n_12189, n14201);
  and g26007 (n14202, \a[14] , n_12189);
  and g26008 (n14203, n_12188, n_12189);
  not g26009 (n_12190, n14202);
  not g26010 (n_12191, n14203);
  and g26011 (n14204, n_12190, n_12191);
  and g26012 (n14205, n_12121, n_12126);
  and g26013 (n14206, n_12113, n_12118);
  and g26014 (n14207, \b[47] , n1627);
  and g26015 (n14208, \b[45] , n1763);
  and g26016 (n14209, \b[46] , n1622);
  and g26022 (n14212, n1630, n7703);
  not g26025 (n_12196, n14213);
  and g26026 (n14214, \a[20] , n_12196);
  not g26027 (n_12197, n14214);
  and g26028 (n14215, \a[20] , n_12197);
  and g26029 (n14216, n_12196, n_12197);
  not g26030 (n_12198, n14215);
  not g26031 (n_12199, n14216);
  and g26032 (n14217, n_12198, n_12199);
  and g26033 (n14218, n_12088, n_12093);
  and g26034 (n14219, n_12049, n_12052);
  and g26035 (n14220, n_11999, n_12005);
  and g26036 (n14221, n_11993, n_11996);
  and g26037 (n14222, n_11975, n_11981);
  and g26038 (n14223, n_11969, n_11972);
  and g26039 (n14224, \b[14] , n9339);
  and g26040 (n14225, \b[12] , n9732);
  and g26041 (n14226, \b[13] , n9334);
  and g26047 (n14229, n1034, n9342);
  not g26050 (n_12204, n14230);
  and g26051 (n14231, \a[53] , n_12204);
  not g26052 (n_12205, n14231);
  and g26053 (n14232, \a[53] , n_12205);
  and g26054 (n14233, n_12204, n_12205);
  not g26055 (n_12206, n14232);
  not g26056 (n_12207, n14233);
  and g26057 (n14234, n_12206, n_12207);
  and g26058 (n14235, n_11950, n_11957);
  and g26059 (n14236, n_11944, n_11947);
  and g26060 (n14237, \b[1] , n13903);
  and g26061 (n14238, \b[2] , n_11555);
  not g26062 (n_12208, n14237);
  not g26063 (n_12209, n14238);
  and g26064 (n14239, n_12208, n_12209);
  and g26065 (n14240, \b[5] , n12668);
  and g26066 (n14241, \b[3] , n13047);
  and g26067 (n14242, \b[4] , n12663);
  and g26073 (n14245, n394, n12671);
  not g26076 (n_12214, n14246);
  and g26077 (n14247, \a[62] , n_12214);
  not g26078 (n_12215, n14247);
  and g26079 (n14248, \a[62] , n_12215);
  and g26080 (n14249, n_12214, n_12215);
  not g26081 (n_12216, n14248);
  not g26082 (n_12217, n14249);
  and g26083 (n14250, n_12216, n_12217);
  not g26084 (n_12218, n14239);
  not g26085 (n_12219, n14250);
  and g26086 (n14251, n_12218, n_12219);
  not g26087 (n_12220, n14251);
  and g26088 (n14252, n_12218, n_12220);
  and g26089 (n14253, n_12219, n_12220);
  not g26090 (n_12221, n14252);
  not g26091 (n_12222, n14253);
  and g26092 (n14254, n_12221, n_12222);
  and g26093 (n14255, n_11926, n_11932);
  and g26094 (n14256, n14254, n14255);
  not g26095 (n_12223, n14254);
  not g26096 (n_12224, n14255);
  and g26097 (n14257, n_12223, n_12224);
  not g26098 (n_12225, n14256);
  not g26099 (n_12226, n14257);
  and g26100 (n14258, n_12225, n_12226);
  and g26101 (n14259, \b[8] , n11531);
  and g26102 (n14260, \b[6] , n11896);
  and g26103 (n14261, \b[7] , n11526);
  and g26109 (n14264, n585, n11534);
  not g26112 (n_12231, n14265);
  and g26113 (n14266, \a[59] , n_12231);
  not g26114 (n_12232, n14266);
  and g26115 (n14267, \a[59] , n_12232);
  and g26116 (n14268, n_12231, n_12232);
  not g26117 (n_12233, n14267);
  not g26118 (n_12234, n14268);
  and g26119 (n14269, n_12233, n_12234);
  not g26120 (n_12235, n14269);
  and g26121 (n14270, n14258, n_12235);
  not g26122 (n_12236, n14258);
  and g26123 (n14271, n_12236, n14269);
  not g26124 (n_12237, n14236);
  not g26125 (n_12238, n14271);
  and g26126 (n14272, n_12237, n_12238);
  not g26127 (n_12239, n14270);
  and g26128 (n14273, n_12239, n14272);
  not g26129 (n_12240, n14273);
  and g26130 (n14274, n_12237, n_12240);
  and g26131 (n14275, n_12239, n_12240);
  and g26132 (n14276, n_12238, n14275);
  not g26133 (n_12241, n14274);
  not g26134 (n_12242, n14276);
  and g26135 (n14277, n_12241, n_12242);
  and g26136 (n14278, \b[11] , n10426);
  and g26137 (n14279, \b[9] , n10796);
  and g26138 (n14280, \b[10] , n10421);
  and g26144 (n14283, n818, n10429);
  not g26147 (n_12247, n14284);
  and g26148 (n14285, \a[56] , n_12247);
  not g26149 (n_12248, n14285);
  and g26150 (n14286, \a[56] , n_12248);
  and g26151 (n14287, n_12247, n_12248);
  not g26152 (n_12249, n14286);
  not g26153 (n_12250, n14287);
  and g26154 (n14288, n_12249, n_12250);
  and g26155 (n14289, n14277, n14288);
  not g26156 (n_12251, n14277);
  not g26157 (n_12252, n14288);
  and g26158 (n14290, n_12251, n_12252);
  not g26159 (n_12253, n14289);
  not g26160 (n_12254, n14290);
  and g26161 (n14291, n_12253, n_12254);
  not g26162 (n_12255, n14235);
  and g26163 (n14292, n_12255, n14291);
  not g26164 (n_12256, n14291);
  and g26165 (n14293, n14235, n_12256);
  not g26166 (n_12257, n14292);
  not g26167 (n_12258, n14293);
  and g26168 (n14294, n_12257, n_12258);
  not g26169 (n_12259, n14234);
  and g26170 (n14295, n_12259, n14294);
  not g26171 (n_12260, n14295);
  and g26172 (n14296, n14294, n_12260);
  and g26173 (n14297, n_12259, n_12260);
  not g26174 (n_12261, n14296);
  not g26175 (n_12262, n14297);
  and g26176 (n14298, n_12261, n_12262);
  not g26177 (n_12263, n14223);
  and g26178 (n14299, n_12263, n14298);
  not g26179 (n_12264, n14298);
  and g26180 (n14300, n14223, n_12264);
  not g26181 (n_12265, n14299);
  not g26182 (n_12266, n14300);
  and g26183 (n14301, n_12265, n_12266);
  and g26184 (n14302, \b[17] , n8362);
  and g26185 (n14303, \b[15] , n8715);
  and g26186 (n14304, \b[16] , n8357);
  and g26192 (n14307, n1356, n8365);
  not g26195 (n_12271, n14308);
  and g26196 (n14309, \a[50] , n_12271);
  not g26197 (n_12272, n14309);
  and g26198 (n14310, \a[50] , n_12272);
  and g26199 (n14311, n_12271, n_12272);
  not g26200 (n_12273, n14310);
  not g26201 (n_12274, n14311);
  and g26202 (n14312, n_12273, n_12274);
  not g26203 (n_12275, n14301);
  not g26204 (n_12276, n14312);
  and g26205 (n14313, n_12275, n_12276);
  and g26206 (n14314, n14301, n14312);
  not g26207 (n_12277, n14313);
  not g26208 (n_12278, n14314);
  and g26209 (n14315, n_12277, n_12278);
  not g26210 (n_12279, n14315);
  and g26211 (n14316, n14222, n_12279);
  not g26212 (n_12280, n14222);
  and g26213 (n14317, n_12280, n14315);
  not g26214 (n_12281, n14316);
  not g26215 (n_12282, n14317);
  and g26216 (n14318, n_12281, n_12282);
  and g26217 (n14319, \b[20] , n7446);
  and g26218 (n14320, \b[18] , n7787);
  and g26219 (n14321, \b[19] , n7441);
  and g26225 (n14324, n1846, n7449);
  not g26228 (n_12287, n14325);
  and g26229 (n14326, \a[47] , n_12287);
  not g26230 (n_12288, n14326);
  and g26231 (n14327, \a[47] , n_12288);
  and g26232 (n14328, n_12287, n_12288);
  not g26233 (n_12289, n14327);
  not g26234 (n_12290, n14328);
  and g26235 (n14329, n_12289, n_12290);
  not g26236 (n_12291, n14329);
  and g26237 (n14330, n14318, n_12291);
  not g26238 (n_12292, n14330);
  and g26239 (n14331, n14318, n_12292);
  and g26240 (n14332, n_12291, n_12292);
  not g26241 (n_12293, n14331);
  not g26242 (n_12294, n14332);
  and g26243 (n14333, n_12293, n_12294);
  not g26244 (n_12295, n14221);
  and g26245 (n14334, n_12295, n14333);
  not g26246 (n_12296, n14333);
  and g26247 (n14335, n14221, n_12296);
  not g26248 (n_12297, n14334);
  not g26249 (n_12298, n14335);
  and g26250 (n14336, n_12297, n_12298);
  and g26251 (n14337, \b[23] , n6595);
  and g26252 (n14338, \b[21] , n6902);
  and g26253 (n14339, \b[22] , n6590);
  and g26259 (n14342, n2300, n6598);
  not g26262 (n_12303, n14343);
  and g26263 (n14344, \a[44] , n_12303);
  not g26264 (n_12304, n14344);
  and g26265 (n14345, \a[44] , n_12304);
  and g26266 (n14346, n_12303, n_12304);
  not g26267 (n_12305, n14345);
  not g26268 (n_12306, n14346);
  and g26269 (n14347, n_12305, n_12306);
  not g26270 (n_12307, n14336);
  not g26271 (n_12308, n14347);
  and g26272 (n14348, n_12307, n_12308);
  and g26273 (n14349, n14336, n14347);
  not g26274 (n_12309, n14348);
  not g26275 (n_12310, n14349);
  and g26276 (n14350, n_12309, n_12310);
  not g26277 (n_12311, n14350);
  and g26278 (n14351, n14220, n_12311);
  not g26279 (n_12312, n14220);
  and g26280 (n14352, n_12312, n14350);
  not g26281 (n_12313, n14351);
  not g26282 (n_12314, n14352);
  and g26283 (n14353, n_12313, n_12314);
  and g26284 (n14354, \b[26] , n5777);
  and g26285 (n14355, \b[24] , n6059);
  and g26286 (n14356, \b[25] , n5772);
  and g26292 (n14359, n2813, n5780);
  not g26295 (n_12319, n14360);
  and g26296 (n14361, \a[41] , n_12319);
  not g26297 (n_12320, n14361);
  and g26298 (n14362, \a[41] , n_12320);
  and g26299 (n14363, n_12319, n_12320);
  not g26300 (n_12321, n14362);
  not g26301 (n_12322, n14363);
  and g26302 (n14364, n_12321, n_12322);
  not g26303 (n_12323, n14364);
  and g26304 (n14365, n14353, n_12323);
  not g26305 (n_12324, n14365);
  and g26306 (n14366, n14353, n_12324);
  and g26307 (n14367, n_12323, n_12324);
  not g26308 (n_12325, n14366);
  not g26309 (n_12326, n14367);
  and g26310 (n14368, n_12325, n_12326);
  and g26311 (n14369, n_12015, n_12021);
  and g26312 (n14370, n14368, n14369);
  not g26313 (n_12327, n14368);
  not g26314 (n_12328, n14369);
  and g26315 (n14371, n_12327, n_12328);
  not g26316 (n_12329, n14370);
  not g26317 (n_12330, n14371);
  and g26318 (n14372, n_12329, n_12330);
  and g26319 (n14373, \b[29] , n5035);
  and g26320 (n14374, \b[27] , n5277);
  and g26321 (n14375, \b[28] , n5030);
  and g26327 (n14378, n3383, n5038);
  not g26330 (n_12335, n14379);
  and g26331 (n14380, \a[38] , n_12335);
  not g26332 (n_12336, n14380);
  and g26333 (n14381, \a[38] , n_12336);
  and g26334 (n14382, n_12335, n_12336);
  not g26335 (n_12337, n14381);
  not g26336 (n_12338, n14382);
  and g26337 (n14383, n_12337, n_12338);
  not g26338 (n_12339, n14383);
  and g26339 (n14384, n14372, n_12339);
  not g26340 (n_12340, n14384);
  and g26341 (n14385, n14372, n_12340);
  and g26342 (n14386, n_12339, n_12340);
  not g26343 (n_12341, n14385);
  not g26344 (n_12342, n14386);
  and g26345 (n14387, n_12341, n_12342);
  and g26346 (n14388, n_12031, n_12037);
  and g26347 (n14389, n14387, n14388);
  not g26348 (n_12343, n14387);
  not g26349 (n_12344, n14388);
  and g26350 (n14390, n_12343, n_12344);
  not g26351 (n_12345, n14389);
  not g26352 (n_12346, n14390);
  and g26353 (n14391, n_12345, n_12346);
  and g26354 (n14392, \b[32] , n4287);
  and g26355 (n14393, \b[30] , n4532);
  and g26356 (n14394, \b[31] , n4282);
  and g26362 (n14397, n4013, n4290);
  not g26365 (n_12351, n14398);
  and g26366 (n14399, \a[35] , n_12351);
  not g26367 (n_12352, n14399);
  and g26368 (n14400, \a[35] , n_12352);
  and g26369 (n14401, n_12351, n_12352);
  not g26370 (n_12353, n14400);
  not g26371 (n_12354, n14401);
  and g26372 (n14402, n_12353, n_12354);
  not g26373 (n_12355, n14402);
  and g26374 (n14403, n14391, n_12355);
  not g26375 (n_12356, n14391);
  and g26376 (n14404, n_12356, n14402);
  not g26377 (n_12357, n14219);
  not g26378 (n_12358, n14404);
  and g26379 (n14405, n_12357, n_12358);
  not g26380 (n_12359, n14403);
  and g26381 (n14406, n_12359, n14405);
  not g26382 (n_12360, n14406);
  and g26383 (n14407, n_12357, n_12360);
  and g26384 (n14408, n_12359, n_12360);
  and g26385 (n14409, n_12358, n14408);
  not g26386 (n_12361, n14407);
  not g26387 (n_12362, n14409);
  and g26388 (n14410, n_12361, n_12362);
  and g26389 (n14411, \b[35] , n3638);
  and g26390 (n14412, \b[33] , n3843);
  and g26391 (n14413, \b[34] , n3633);
  and g26397 (n14416, n3641, n4696);
  not g26400 (n_12367, n14417);
  and g26401 (n14418, \a[32] , n_12367);
  not g26402 (n_12368, n14418);
  and g26403 (n14419, \a[32] , n_12368);
  and g26404 (n14420, n_12367, n_12368);
  not g26405 (n_12369, n14419);
  not g26406 (n_12370, n14420);
  and g26407 (n14421, n_12369, n_12370);
  not g26408 (n_12371, n14410);
  not g26409 (n_12372, n14421);
  and g26410 (n14422, n_12371, n_12372);
  not g26411 (n_12373, n14422);
  and g26412 (n14423, n_12371, n_12373);
  and g26413 (n14424, n_12372, n_12373);
  not g26414 (n_12374, n14423);
  not g26415 (n_12375, n14424);
  and g26416 (n14425, n_12374, n_12375);
  and g26417 (n14426, n_12055, n_12062);
  and g26418 (n14427, n14425, n14426);
  not g26419 (n_12376, n14425);
  not g26420 (n_12377, n14426);
  and g26421 (n14428, n_12376, n_12377);
  not g26422 (n_12378, n14427);
  not g26423 (n_12379, n14428);
  and g26424 (n14429, n_12378, n_12379);
  and g26425 (n14430, \b[38] , n3050);
  and g26426 (n14431, \b[36] , n3243);
  and g26427 (n14432, \b[37] , n3045);
  and g26433 (n14435, n3053, n5205);
  not g26436 (n_12384, n14436);
  and g26437 (n14437, \a[29] , n_12384);
  not g26438 (n_12385, n14437);
  and g26439 (n14438, \a[29] , n_12385);
  and g26440 (n14439, n_12384, n_12385);
  not g26441 (n_12386, n14438);
  not g26442 (n_12387, n14439);
  and g26443 (n14440, n_12386, n_12387);
  not g26444 (n_12388, n14440);
  and g26445 (n14441, n14429, n_12388);
  not g26446 (n_12389, n14441);
  and g26447 (n14442, n14429, n_12389);
  and g26448 (n14443, n_12388, n_12389);
  not g26449 (n_12390, n14442);
  not g26450 (n_12391, n14443);
  and g26451 (n14444, n_12390, n_12391);
  and g26452 (n14445, n_12072, n_12078);
  and g26453 (n14446, n14444, n14445);
  not g26454 (n_12392, n14444);
  not g26455 (n_12393, n14445);
  and g26456 (n14447, n_12392, n_12393);
  not g26457 (n_12394, n14446);
  not g26458 (n_12395, n14447);
  and g26459 (n14448, n_12394, n_12395);
  and g26460 (n14449, \b[41] , n2539);
  and g26461 (n14450, \b[39] , n2685);
  and g26462 (n14451, \b[40] , n2534);
  and g26468 (n14454, n2542, n6219);
  not g26471 (n_12400, n14455);
  and g26472 (n14456, \a[26] , n_12400);
  not g26473 (n_12401, n14456);
  and g26474 (n14457, \a[26] , n_12401);
  and g26475 (n14458, n_12400, n_12401);
  not g26476 (n_12402, n14457);
  not g26477 (n_12403, n14458);
  and g26478 (n14459, n_12402, n_12403);
  not g26479 (n_12404, n14459);
  and g26480 (n14460, n14448, n_12404);
  not g26481 (n_12405, n14448);
  and g26482 (n14461, n_12405, n14459);
  not g26483 (n_12406, n14218);
  not g26484 (n_12407, n14461);
  and g26485 (n14462, n_12406, n_12407);
  not g26486 (n_12408, n14460);
  and g26487 (n14463, n_12408, n14462);
  not g26488 (n_12409, n14463);
  and g26489 (n14464, n_12406, n_12409);
  and g26490 (n14465, n_12408, n_12409);
  and g26491 (n14466, n_12407, n14465);
  not g26492 (n_12410, n14464);
  not g26493 (n_12411, n14466);
  and g26494 (n14467, n_12410, n_12411);
  and g26495 (n14468, \b[44] , n2048);
  and g26496 (n14469, \b[42] , n2198);
  and g26497 (n14470, \b[43] , n2043);
  and g26503 (n14473, n2051, n7072);
  not g26506 (n_12416, n14474);
  and g26507 (n14475, \a[23] , n_12416);
  not g26508 (n_12417, n14475);
  and g26509 (n14476, \a[23] , n_12417);
  and g26510 (n14477, n_12416, n_12417);
  not g26511 (n_12418, n14476);
  not g26512 (n_12419, n14477);
  and g26513 (n14478, n_12418, n_12419);
  not g26514 (n_12420, n14467);
  not g26515 (n_12421, n14478);
  and g26516 (n14479, n_12420, n_12421);
  not g26517 (n_12422, n14479);
  and g26518 (n14480, n_12420, n_12422);
  and g26519 (n14481, n_12421, n_12422);
  not g26520 (n_12423, n14480);
  not g26521 (n_12424, n14481);
  and g26522 (n14482, n_12423, n_12424);
  and g26523 (n14483, n_12104, n_12105);
  not g26524 (n_12425, n14483);
  and g26525 (n14484, n_12110, n_12425);
  not g26526 (n_12426, n14482);
  not g26527 (n_12427, n14484);
  and g26528 (n14485, n_12426, n_12427);
  and g26529 (n14486, n14482, n14484);
  not g26530 (n_12428, n14485);
  not g26531 (n_12429, n14486);
  and g26532 (n14487, n_12428, n_12429);
  not g26533 (n_12430, n14217);
  and g26534 (n14488, n_12430, n14487);
  not g26535 (n_12431, n14488);
  and g26536 (n14489, n_12430, n_12431);
  and g26537 (n14490, n14487, n_12431);
  not g26538 (n_12432, n14489);
  not g26539 (n_12433, n14490);
  and g26540 (n14491, n_12432, n_12433);
  not g26541 (n_12434, n14206);
  not g26542 (n_12435, n14491);
  and g26543 (n14492, n_12434, n_12435);
  not g26544 (n_12436, n14492);
  and g26545 (n14493, n_12434, n_12436);
  and g26546 (n14494, n_12435, n_12436);
  not g26547 (n_12437, n14493);
  not g26548 (n_12438, n14494);
  and g26549 (n14495, n_12437, n_12438);
  and g26550 (n14496, \b[50] , n1302);
  and g26551 (n14497, \b[48] , n1391);
  and g26552 (n14498, \b[49] , n1297);
  and g26558 (n14501, n1305, n8949);
  not g26561 (n_12443, n14502);
  and g26562 (n14503, \a[17] , n_12443);
  not g26563 (n_12444, n14503);
  and g26564 (n14504, \a[17] , n_12444);
  and g26565 (n14505, n_12443, n_12444);
  not g26566 (n_12445, n14504);
  not g26567 (n_12446, n14505);
  and g26568 (n14506, n_12445, n_12446);
  and g26569 (n14507, n14495, n14506);
  not g26570 (n_12447, n14495);
  not g26571 (n_12448, n14506);
  and g26572 (n14508, n_12447, n_12448);
  not g26573 (n_12449, n14507);
  not g26574 (n_12450, n14508);
  and g26575 (n14509, n_12449, n_12450);
  not g26576 (n_12451, n14205);
  and g26577 (n14510, n_12451, n14509);
  not g26578 (n_12452, n14509);
  and g26579 (n14511, n14205, n_12452);
  not g26580 (n_12453, n14510);
  not g26581 (n_12454, n14511);
  and g26582 (n14512, n_12453, n_12454);
  not g26583 (n_12455, n14204);
  and g26584 (n14513, n_12455, n14512);
  not g26585 (n_12456, n14513);
  and g26586 (n14514, n14512, n_12456);
  and g26587 (n14515, n_12455, n_12456);
  not g26588 (n_12457, n14514);
  not g26589 (n_12458, n14515);
  and g26590 (n14516, n_12457, n_12458);
  and g26591 (n14517, n_12130, n_12134);
  and g26592 (n14518, n14516, n14517);
  not g26593 (n_12459, n14516);
  not g26594 (n_12460, n14517);
  and g26595 (n14519, n_12459, n_12460);
  not g26596 (n_12461, n14518);
  not g26597 (n_12462, n14519);
  and g26598 (n14520, n_12461, n_12462);
  and g26599 (n14521, \b[56] , n700);
  and g26600 (n14522, \b[54] , n767);
  and g26601 (n14523, \b[55] , n695);
  and g26607 (n14526, n703, n10708);
  not g26610 (n_12467, n14527);
  and g26611 (n14528, \a[11] , n_12467);
  not g26612 (n_12468, n14528);
  and g26613 (n14529, \a[11] , n_12468);
  and g26614 (n14530, n_12467, n_12468);
  not g26615 (n_12469, n14529);
  not g26616 (n_12470, n14530);
  and g26617 (n14531, n_12469, n_12470);
  not g26618 (n_12471, n14520);
  and g26619 (n14532, n_12471, n14531);
  not g26620 (n_12472, n14531);
  and g26621 (n14533, n14520, n_12472);
  not g26622 (n_12473, n14532);
  not g26623 (n_12474, n14533);
  and g26624 (n14534, n_12473, n_12474);
  and g26625 (n14535, \b[59] , n511);
  and g26626 (n14536, \b[57] , n541);
  and g26627 (n14537, \b[58] , n506);
  and g26633 (n14540, n514, n12179);
  not g26636 (n_12479, n14541);
  and g26637 (n14542, \a[8] , n_12479);
  not g26638 (n_12480, n14542);
  and g26639 (n14543, \a[8] , n_12480);
  and g26640 (n14544, n_12479, n_12480);
  not g26641 (n_12481, n14543);
  not g26642 (n_12482, n14544);
  and g26643 (n14545, n_12481, n_12482);
  not g26644 (n_12483, n14545);
  and g26645 (n14546, n14534, n_12483);
  not g26646 (n_12484, n14546);
  and g26647 (n14547, n14534, n_12484);
  and g26648 (n14548, n_12483, n_12484);
  not g26649 (n_12485, n14547);
  not g26650 (n_12486, n14548);
  and g26651 (n14549, n_12485, n_12486);
  and g26652 (n14550, n_12138, n_12142);
  and g26653 (n14551, n14549, n14550);
  not g26654 (n_12487, n14549);
  not g26655 (n_12488, n14550);
  and g26656 (n14552, n_12487, n_12488);
  not g26657 (n_12489, n14551);
  not g26658 (n_12490, n14552);
  and g26659 (n14553, n_12489, n_12490);
  and g26660 (n14554, \b[62] , n362);
  and g26661 (n14555, \b[60] , n403);
  and g26662 (n14556, \b[61] , n357);
  and g26668 (n14559, n365, n13370);
  not g26671 (n_12495, n14560);
  and g26672 (n14561, \a[5] , n_12495);
  not g26673 (n_12496, n14561);
  and g26674 (n14562, \a[5] , n_12496);
  and g26675 (n14563, n_12495, n_12496);
  not g26676 (n_12497, n14562);
  not g26677 (n_12498, n14563);
  and g26678 (n14564, n_12497, n_12498);
  not g26679 (n_12499, n14564);
  and g26680 (n14565, n14553, n_12499);
  not g26681 (n_12500, n14565);
  and g26682 (n14566, n14553, n_12500);
  and g26683 (n14567, n_12499, n_12500);
  not g26684 (n_12501, n14566);
  not g26685 (n_12502, n14567);
  and g26686 (n14568, n_12501, n_12502);
  and g26687 (n14569, n_12164, n_12165);
  not g26688 (n_12503, n14569);
  and g26689 (n14570, n_12153, n_12503);
  and g26690 (n14571, n269, n13797);
  not g26691 (n_12504, n14571);
  and g26692 (n14572, n_5, n_12504);
  and g26693 (n14573, \b[63] , n284);
  not g26694 (n_12505, n14573);
  and g26695 (n14574, n_12504, n_12505);
  not g26696 (n_12506, n14574);
  and g26697 (n14575, \a[2] , n_12506);
  not g26698 (n_12507, n14572);
  not g26699 (n_12508, n14575);
  and g26700 (n14576, n_12507, n_12508);
  not g26701 (n_12509, n14570);
  and g26702 (n14577, n_12509, n14576);
  not g26703 (n_12510, n14576);
  and g26704 (n14578, n14570, n_12510);
  not g26705 (n_12511, n14577);
  not g26706 (n_12512, n14578);
  and g26707 (n14579, n_12511, n_12512);
  not g26708 (n_12513, n14568);
  and g26709 (n14580, n_12513, n14579);
  not g26710 (n_12514, n14580);
  and g26711 (n14581, n_12513, n_12514);
  and g26712 (n14582, n14579, n_12514);
  not g26713 (n_12515, n14581);
  not g26714 (n_12516, n14582);
  and g26715 (n14583, n_12515, n_12516);
  and g26716 (n14584, n_12170, n_12174);
  and g26717 (n14585, n14583, n14584);
  not g26718 (n_12517, n14583);
  not g26719 (n_12518, n14584);
  and g26720 (n14586, n_12517, n_12518);
  not g26721 (n_12519, n14585);
  not g26722 (n_12520, n14586);
  and g26723 (n14587, n_12519, n_12520);
  and g26724 (n14588, n_12178, n_12182);
  not g26725 (n_12521, n14588);
  and g26726 (n14589, n14587, n_12521);
  not g26727 (n_12522, n14587);
  and g26728 (n14590, n_12522, n14588);
  not g26729 (n_12523, n14589);
  not g26730 (n_12524, n14590);
  and g26731 (\f[65] , n_12523, n_12524);
  and g26732 (n14592, n_12490, n_12500);
  and g26733 (n14593, \b[63] , n362);
  and g26734 (n14594, \b[61] , n403);
  and g26735 (n14595, \b[62] , n357);
  and g26741 (n14598, n365, n13771);
  not g26744 (n_12529, n14599);
  and g26745 (n14600, \a[5] , n_12529);
  not g26746 (n_12530, n14600);
  and g26747 (n14601, \a[5] , n_12530);
  and g26748 (n14602, n_12529, n_12530);
  not g26749 (n_12531, n14601);
  not g26750 (n_12532, n14602);
  and g26751 (n14603, n_12531, n_12532);
  not g26752 (n_12533, n14592);
  not g26753 (n_12534, n14603);
  and g26754 (n14604, n_12533, n_12534);
  not g26755 (n_12535, n14604);
  and g26756 (n14605, n_12533, n_12535);
  and g26757 (n14606, n_12534, n_12535);
  not g26758 (n_12536, n14605);
  not g26759 (n_12537, n14606);
  and g26760 (n14607, n_12536, n_12537);
  and g26761 (n14608, \b[57] , n700);
  and g26762 (n14609, \b[55] , n767);
  and g26763 (n14610, \b[56] , n695);
  and g26769 (n14613, n703, n11410);
  not g26772 (n_12542, n14614);
  and g26773 (n14615, \a[11] , n_12542);
  not g26774 (n_12543, n14615);
  and g26775 (n14616, \a[11] , n_12543);
  and g26776 (n14617, n_12542, n_12543);
  not g26777 (n_12544, n14616);
  not g26778 (n_12545, n14617);
  and g26779 (n14618, n_12544, n_12545);
  and g26780 (n14619, n_12456, n_12462);
  and g26781 (n14620, n14618, n14619);
  not g26782 (n_12546, n14618);
  not g26783 (n_12547, n14619);
  and g26784 (n14621, n_12546, n_12547);
  not g26785 (n_12548, n14620);
  not g26786 (n_12549, n14621);
  and g26787 (n14622, n_12548, n_12549);
  and g26788 (n14623, \b[51] , n1302);
  and g26789 (n14624, \b[49] , n1391);
  and g26790 (n14625, \b[50] , n1297);
  and g26796 (n14628, n1305, n8976);
  not g26799 (n_12554, n14629);
  and g26800 (n14630, \a[17] , n_12554);
  not g26801 (n_12555, n14630);
  and g26802 (n14631, \a[17] , n_12555);
  and g26803 (n14632, n_12554, n_12555);
  not g26804 (n_12556, n14631);
  not g26805 (n_12557, n14632);
  and g26806 (n14633, n_12556, n_12557);
  and g26807 (n14634, n_12431, n_12436);
  and g26808 (n14635, n14633, n14634);
  not g26809 (n_12558, n14633);
  not g26810 (n_12559, n14634);
  and g26811 (n14636, n_12558, n_12559);
  not g26812 (n_12560, n14635);
  not g26813 (n_12561, n14636);
  and g26814 (n14637, n_12560, n_12561);
  and g26815 (n14638, \b[48] , n1627);
  and g26816 (n14639, \b[46] , n1763);
  and g26817 (n14640, \b[47] , n1622);
  and g26823 (n14643, n1630, n8009);
  not g26826 (n_12566, n14644);
  and g26827 (n14645, \a[20] , n_12566);
  not g26828 (n_12567, n14645);
  and g26829 (n14646, \a[20] , n_12567);
  and g26830 (n14647, n_12566, n_12567);
  not g26831 (n_12568, n14646);
  not g26832 (n_12569, n14647);
  and g26833 (n14648, n_12568, n_12569);
  and g26834 (n14649, n_12422, n_12428);
  and g26835 (n14650, n14648, n14649);
  not g26836 (n_12570, n14648);
  not g26837 (n_12571, n14649);
  and g26838 (n14651, n_12570, n_12571);
  not g26839 (n_12572, n14650);
  not g26840 (n_12573, n14651);
  and g26841 (n14652, n_12572, n_12573);
  and g26842 (n14653, \b[45] , n2048);
  and g26843 (n14654, \b[43] , n2198);
  and g26844 (n14655, \b[44] , n2043);
  and g26850 (n14658, n2051, n7361);
  not g26853 (n_12578, n14659);
  and g26854 (n14660, \a[23] , n_12578);
  not g26855 (n_12579, n14660);
  and g26856 (n14661, \a[23] , n_12579);
  and g26857 (n14662, n_12578, n_12579);
  not g26858 (n_12580, n14661);
  not g26859 (n_12581, n14662);
  and g26860 (n14663, n_12580, n_12581);
  not g26861 (n_12582, n14465);
  and g26862 (n14664, n_12582, n14663);
  not g26863 (n_12583, n14663);
  and g26864 (n14665, n14465, n_12583);
  not g26865 (n_12584, n14664);
  not g26866 (n_12585, n14665);
  and g26867 (n14666, n_12584, n_12585);
  and g26868 (n14667, \b[42] , n2539);
  and g26869 (n14668, \b[40] , n2685);
  and g26870 (n14669, \b[41] , n2534);
  and g26876 (n14672, n2542, n6489);
  not g26879 (n_12590, n14673);
  and g26880 (n14674, \a[26] , n_12590);
  not g26881 (n_12591, n14674);
  and g26882 (n14675, \a[26] , n_12591);
  and g26883 (n14676, n_12590, n_12591);
  not g26884 (n_12592, n14675);
  not g26885 (n_12593, n14676);
  and g26886 (n14677, n_12592, n_12593);
  and g26887 (n14678, n_12389, n_12395);
  and g26888 (n14679, n14677, n14678);
  not g26889 (n_12594, n14677);
  not g26890 (n_12595, n14678);
  and g26891 (n14680, n_12594, n_12595);
  not g26892 (n_12596, n14679);
  not g26893 (n_12597, n14680);
  and g26894 (n14681, n_12596, n_12597);
  and g26895 (n14682, n_12373, n_12379);
  and g26896 (n14683, \b[39] , n3050);
  and g26897 (n14684, \b[37] , n3243);
  and g26898 (n14685, \b[38] , n3045);
  not g26899 (n_12598, n14684);
  not g26900 (n_12599, n14685);
  and g26901 (n14686, n_12598, n_12599);
  not g26902 (n_12600, n14683);
  and g26903 (n14687, n_12600, n14686);
  not g26904 (n_12601, n3053);
  and g26905 (n14688, n_12601, n14687);
  not g26906 (n_12602, n5451);
  and g26907 (n14689, n_12602, n14687);
  not g26908 (n_12603, n14688);
  not g26909 (n_12604, n14689);
  and g26910 (n14690, n_12603, n_12604);
  not g26911 (n_12605, n14690);
  and g26912 (n14691, \a[29] , n_12605);
  and g26913 (n14692, n_2476, n14690);
  not g26914 (n_12606, n14691);
  not g26915 (n_12607, n14692);
  and g26916 (n14693, n_12606, n_12607);
  not g26917 (n_12608, n14682);
  not g26918 (n_12609, n14693);
  and g26919 (n14694, n_12608, n_12609);
  and g26920 (n14695, n14682, n14693);
  not g26921 (n_12610, n14694);
  not g26922 (n_12611, n14695);
  and g26923 (n14696, n_12610, n_12611);
  and g26924 (n14697, \b[33] , n4287);
  and g26925 (n14698, \b[31] , n4532);
  and g26926 (n14699, \b[32] , n4282);
  and g26932 (n14702, n4223, n4290);
  not g26935 (n_12616, n14703);
  and g26936 (n14704, \a[35] , n_12616);
  not g26937 (n_12617, n14704);
  and g26938 (n14705, \a[35] , n_12617);
  and g26939 (n14706, n_12616, n_12617);
  not g26940 (n_12618, n14705);
  not g26941 (n_12619, n14706);
  and g26942 (n14707, n_12618, n_12619);
  and g26943 (n14708, \b[24] , n6595);
  and g26944 (n14709, \b[22] , n6902);
  and g26945 (n14710, \b[23] , n6590);
  and g26951 (n14713, n2458, n6598);
  not g26954 (n_12624, n14714);
  and g26955 (n14715, \a[44] , n_12624);
  not g26956 (n_12625, n14715);
  and g26957 (n14716, \a[44] , n_12625);
  and g26958 (n14717, n_12624, n_12625);
  not g26959 (n_12626, n14716);
  not g26960 (n_12627, n14717);
  and g26961 (n14718, n_12626, n_12627);
  and g26962 (n14719, \b[15] , n9339);
  and g26963 (n14720, \b[13] , n9732);
  and g26964 (n14721, \b[14] , n9334);
  and g26970 (n14724, n1131, n9342);
  not g26973 (n_12632, n14725);
  and g26974 (n14726, \a[53] , n_12632);
  not g26975 (n_12633, n14726);
  and g26976 (n14727, \a[53] , n_12633);
  and g26977 (n14728, n_12632, n_12633);
  not g26978 (n_12634, n14727);
  not g26979 (n_12635, n14728);
  and g26980 (n14729, n_12634, n_12635);
  and g26981 (n14730, n_12254, n_12257);
  and g26982 (n14731, n_12220, n_12226);
  and g26983 (n14732, \b[2] , n13903);
  and g26984 (n14733, \b[3] , n_11555);
  not g26985 (n_12636, n14732);
  not g26986 (n_12637, n14733);
  and g26987 (n14734, n_12636, n_12637);
  not g26988 (n_12638, n14734);
  and g26989 (n14735, \a[2] , n_12638);
  and g26990 (n14736, n_5, n14734);
  not g26991 (n_12639, n14735);
  not g26992 (n_12640, n14736);
  and g26993 (n14737, n_12639, n_12640);
  and g26994 (n14738, \b[6] , n12668);
  and g26995 (n14739, \b[4] , n13047);
  and g26996 (n14740, \b[5] , n12663);
  not g26997 (n_12641, n14739);
  not g26998 (n_12642, n14740);
  and g26999 (n14741, n_12641, n_12642);
  not g27000 (n_12643, n14738);
  and g27001 (n14742, n_12643, n14741);
  not g27002 (n_12644, n12671);
  and g27003 (n14743, n_12644, n14742);
  not g27004 (n_12645, n459);
  and g27005 (n14744, n_12645, n14742);
  not g27006 (n_12646, n14743);
  not g27007 (n_12647, n14744);
  and g27008 (n14745, n_12646, n_12647);
  not g27009 (n_12648, n14745);
  and g27010 (n14746, \a[62] , n_12648);
  and g27011 (n14747, n_10843, n14745);
  not g27012 (n_12649, n14746);
  not g27013 (n_12650, n14747);
  and g27014 (n14748, n_12649, n_12650);
  not g27015 (n_12651, n14748);
  and g27016 (n14749, n14737, n_12651);
  not g27017 (n_12652, n14737);
  and g27018 (n14750, n_12652, n14748);
  not g27019 (n_12653, n14749);
  not g27020 (n_12654, n14750);
  and g27021 (n14751, n_12653, n_12654);
  not g27022 (n_12655, n14731);
  and g27023 (n14752, n_12655, n14751);
  not g27024 (n_12656, n14751);
  and g27025 (n14753, n14731, n_12656);
  not g27026 (n_12657, n14752);
  not g27027 (n_12658, n14753);
  and g27028 (n14754, n_12657, n_12658);
  and g27029 (n14755, \b[9] , n11531);
  and g27030 (n14756, \b[7] , n11896);
  and g27031 (n14757, \b[8] , n11526);
  and g27037 (n14760, n651, n11534);
  not g27040 (n_12663, n14761);
  and g27041 (n14762, \a[59] , n_12663);
  not g27042 (n_12664, n14762);
  and g27043 (n14763, \a[59] , n_12664);
  and g27044 (n14764, n_12663, n_12664);
  not g27045 (n_12665, n14763);
  not g27046 (n_12666, n14764);
  and g27047 (n14765, n_12665, n_12666);
  not g27048 (n_12667, n14765);
  and g27049 (n14766, n14754, n_12667);
  not g27050 (n_12668, n14766);
  and g27051 (n14767, n14754, n_12668);
  and g27052 (n14768, n_12667, n_12668);
  not g27053 (n_12669, n14767);
  not g27054 (n_12670, n14768);
  and g27055 (n14769, n_12669, n_12670);
  not g27056 (n_12671, n14275);
  and g27057 (n14770, n_12671, n14769);
  not g27058 (n_12672, n14769);
  and g27059 (n14771, n14275, n_12672);
  not g27060 (n_12673, n14770);
  not g27061 (n_12674, n14771);
  and g27062 (n14772, n_12673, n_12674);
  and g27063 (n14773, \b[12] , n10426);
  and g27064 (n14774, \b[10] , n10796);
  and g27065 (n14775, \b[11] , n10421);
  and g27071 (n14778, n842, n10429);
  not g27074 (n_12679, n14779);
  and g27075 (n14780, \a[56] , n_12679);
  not g27076 (n_12680, n14780);
  and g27077 (n14781, \a[56] , n_12680);
  and g27078 (n14782, n_12679, n_12680);
  not g27079 (n_12681, n14781);
  not g27080 (n_12682, n14782);
  and g27081 (n14783, n_12681, n_12682);
  and g27082 (n14784, n14772, n14783);
  not g27083 (n_12683, n14772);
  not g27084 (n_12684, n14783);
  and g27085 (n14785, n_12683, n_12684);
  not g27086 (n_12685, n14784);
  not g27087 (n_12686, n14785);
  and g27088 (n14786, n_12685, n_12686);
  not g27089 (n_12687, n14730);
  and g27090 (n14787, n_12687, n14786);
  not g27091 (n_12688, n14786);
  and g27092 (n14788, n14730, n_12688);
  not g27093 (n_12689, n14787);
  not g27094 (n_12690, n14788);
  and g27095 (n14789, n_12689, n_12690);
  not g27096 (n_12691, n14729);
  and g27097 (n14790, n_12691, n14789);
  not g27098 (n_12692, n14790);
  and g27099 (n14791, n14789, n_12692);
  and g27100 (n14792, n_12691, n_12692);
  not g27101 (n_12693, n14791);
  not g27102 (n_12694, n14792);
  and g27103 (n14793, n_12693, n_12694);
  and g27104 (n14794, n_12263, n_12264);
  not g27105 (n_12695, n14794);
  and g27106 (n14795, n_12260, n_12695);
  and g27107 (n14796, n14793, n14795);
  not g27108 (n_12696, n14793);
  not g27109 (n_12697, n14795);
  and g27110 (n14797, n_12696, n_12697);
  not g27111 (n_12698, n14796);
  not g27112 (n_12699, n14797);
  and g27113 (n14798, n_12698, n_12699);
  and g27114 (n14799, \b[18] , n8362);
  and g27115 (n14800, \b[16] , n8715);
  and g27116 (n14801, \b[17] , n8357);
  and g27122 (n14804, n1566, n8365);
  not g27125 (n_12704, n14805);
  and g27126 (n14806, \a[50] , n_12704);
  not g27127 (n_12705, n14806);
  and g27128 (n14807, \a[50] , n_12705);
  and g27129 (n14808, n_12704, n_12705);
  not g27130 (n_12706, n14807);
  not g27131 (n_12707, n14808);
  and g27132 (n14809, n_12706, n_12707);
  not g27133 (n_12708, n14809);
  and g27134 (n14810, n14798, n_12708);
  not g27135 (n_12709, n14810);
  and g27136 (n14811, n14798, n_12709);
  and g27137 (n14812, n_12708, n_12709);
  not g27138 (n_12710, n14811);
  not g27139 (n_12711, n14812);
  and g27140 (n14813, n_12710, n_12711);
  and g27141 (n14814, n_12277, n_12282);
  and g27142 (n14815, n14813, n14814);
  not g27143 (n_12712, n14813);
  not g27144 (n_12713, n14814);
  and g27145 (n14816, n_12712, n_12713);
  not g27146 (n_12714, n14815);
  not g27147 (n_12715, n14816);
  and g27148 (n14817, n_12714, n_12715);
  and g27149 (n14818, \b[21] , n7446);
  and g27150 (n14819, \b[19] , n7787);
  and g27151 (n14820, \b[20] , n7441);
  and g27157 (n14823, n1984, n7449);
  not g27160 (n_12720, n14824);
  and g27161 (n14825, \a[47] , n_12720);
  not g27162 (n_12721, n14825);
  and g27163 (n14826, \a[47] , n_12721);
  and g27164 (n14827, n_12720, n_12721);
  not g27165 (n_12722, n14826);
  not g27166 (n_12723, n14827);
  and g27167 (n14828, n_12722, n_12723);
  not g27168 (n_12724, n14817);
  and g27169 (n14829, n_12724, n14828);
  not g27170 (n_12725, n14828);
  and g27171 (n14830, n14817, n_12725);
  not g27172 (n_12726, n14829);
  not g27173 (n_12727, n14830);
  and g27174 (n14831, n_12726, n_12727);
  and g27175 (n14832, n_12295, n_12296);
  not g27176 (n_12728, n14832);
  and g27177 (n14833, n_12292, n_12728);
  not g27178 (n_12729, n14833);
  and g27179 (n14834, n14831, n_12729);
  not g27180 (n_12730, n14831);
  and g27181 (n14835, n_12730, n14833);
  not g27182 (n_12731, n14834);
  not g27183 (n_12732, n14835);
  and g27184 (n14836, n_12731, n_12732);
  not g27185 (n_12733, n14718);
  and g27186 (n14837, n_12733, n14836);
  not g27187 (n_12734, n14837);
  and g27188 (n14838, n14836, n_12734);
  and g27189 (n14839, n_12733, n_12734);
  not g27190 (n_12735, n14838);
  not g27191 (n_12736, n14839);
  and g27192 (n14840, n_12735, n_12736);
  and g27193 (n14841, n_12309, n_12314);
  and g27194 (n14842, n14840, n14841);
  not g27195 (n_12737, n14840);
  not g27196 (n_12738, n14841);
  and g27197 (n14843, n_12737, n_12738);
  not g27198 (n_12739, n14842);
  not g27199 (n_12740, n14843);
  and g27200 (n14844, n_12739, n_12740);
  and g27201 (n14845, \b[27] , n5777);
  and g27202 (n14846, \b[25] , n6059);
  and g27203 (n14847, \b[26] , n5772);
  and g27209 (n14850, n2990, n5780);
  not g27212 (n_12745, n14851);
  and g27213 (n14852, \a[41] , n_12745);
  not g27214 (n_12746, n14852);
  and g27215 (n14853, \a[41] , n_12746);
  and g27216 (n14854, n_12745, n_12746);
  not g27217 (n_12747, n14853);
  not g27218 (n_12748, n14854);
  and g27219 (n14855, n_12747, n_12748);
  not g27220 (n_12749, n14855);
  and g27221 (n14856, n14844, n_12749);
  not g27222 (n_12750, n14856);
  and g27223 (n14857, n14844, n_12750);
  and g27224 (n14858, n_12749, n_12750);
  not g27225 (n_12751, n14857);
  not g27226 (n_12752, n14858);
  and g27227 (n14859, n_12751, n_12752);
  and g27228 (n14860, n_12324, n_12330);
  and g27229 (n14861, n14859, n14860);
  not g27230 (n_12753, n14859);
  not g27231 (n_12754, n14860);
  and g27232 (n14862, n_12753, n_12754);
  not g27233 (n_12755, n14861);
  not g27234 (n_12756, n14862);
  and g27235 (n14863, n_12755, n_12756);
  and g27236 (n14864, \b[30] , n5035);
  and g27237 (n14865, \b[28] , n5277);
  and g27238 (n14866, \b[29] , n5030);
  and g27244 (n14869, n3577, n5038);
  not g27247 (n_12761, n14870);
  and g27248 (n14871, \a[38] , n_12761);
  not g27249 (n_12762, n14871);
  and g27250 (n14872, \a[38] , n_12762);
  and g27251 (n14873, n_12761, n_12762);
  not g27252 (n_12763, n14872);
  not g27253 (n_12764, n14873);
  and g27254 (n14874, n_12763, n_12764);
  not g27255 (n_12765, n14863);
  and g27256 (n14875, n_12765, n14874);
  not g27257 (n_12766, n14874);
  and g27258 (n14876, n14863, n_12766);
  not g27259 (n_12767, n14875);
  not g27260 (n_12768, n14876);
  and g27261 (n14877, n_12767, n_12768);
  and g27262 (n14878, n_12340, n_12346);
  not g27263 (n_12769, n14878);
  and g27264 (n14879, n14877, n_12769);
  not g27265 (n_12770, n14877);
  and g27266 (n14880, n_12770, n14878);
  not g27267 (n_12771, n14879);
  not g27268 (n_12772, n14880);
  and g27269 (n14881, n_12771, n_12772);
  not g27270 (n_12773, n14707);
  and g27271 (n14882, n_12773, n14881);
  not g27272 (n_12774, n14882);
  and g27273 (n14883, n14881, n_12774);
  and g27274 (n14884, n_12773, n_12774);
  not g27275 (n_12775, n14883);
  not g27276 (n_12776, n14884);
  and g27277 (n14885, n_12775, n_12776);
  and g27278 (n14886, \b[36] , n3638);
  and g27279 (n14887, \b[34] , n3843);
  and g27280 (n14888, \b[35] , n3633);
  not g27281 (n_12777, n14887);
  not g27282 (n_12778, n14888);
  and g27283 (n14889, n_12777, n_12778);
  not g27284 (n_12779, n14886);
  and g27285 (n14890, n_12779, n14889);
  not g27286 (n_12780, n3641);
  and g27287 (n14891, n_12780, n14890);
  not g27288 (n_12781, n4922);
  and g27289 (n14892, n_12781, n14890);
  not g27290 (n_12782, n14891);
  not g27291 (n_12783, n14892);
  and g27292 (n14893, n_12782, n_12783);
  not g27293 (n_12784, n14893);
  and g27294 (n14894, \a[32] , n_12784);
  and g27295 (n14895, n_2992, n14893);
  not g27296 (n_12785, n14894);
  not g27297 (n_12786, n14895);
  and g27298 (n14896, n_12785, n_12786);
  not g27299 (n_12787, n14408);
  not g27300 (n_12788, n14896);
  and g27301 (n14897, n_12787, n_12788);
  not g27302 (n_12789, n14897);
  and g27303 (n14898, n_12787, n_12789);
  and g27304 (n14899, n_12788, n_12789);
  not g27305 (n_12790, n14898);
  not g27306 (n_12791, n14899);
  and g27307 (n14900, n_12790, n_12791);
  not g27308 (n_12792, n14885);
  not g27309 (n_12793, n14900);
  and g27310 (n14901, n_12792, n_12793);
  not g27311 (n_12794, n14901);
  and g27312 (n14902, n_12792, n_12794);
  and g27313 (n14903, n_12793, n_12794);
  not g27314 (n_12795, n14902);
  not g27315 (n_12796, n14903);
  and g27316 (n14904, n_12795, n_12796);
  not g27317 (n_12797, n14904);
  and g27318 (n14905, n14696, n_12797);
  not g27319 (n_12798, n14905);
  and g27320 (n14906, n14696, n_12798);
  and g27321 (n14907, n_12797, n_12798);
  not g27322 (n_12799, n14906);
  not g27323 (n_12800, n14907);
  and g27324 (n14908, n_12799, n_12800);
  not g27325 (n_12801, n14908);
  and g27326 (n14909, n14681, n_12801);
  not g27327 (n_12802, n14681);
  and g27328 (n14910, n_12802, n14908);
  not g27329 (n_12803, n14666);
  not g27330 (n_12804, n14910);
  and g27331 (n14911, n_12803, n_12804);
  not g27332 (n_12805, n14909);
  and g27333 (n14912, n_12805, n14911);
  not g27334 (n_12806, n14912);
  and g27335 (n14913, n_12803, n_12806);
  and g27336 (n14914, n_12804, n_12806);
  and g27337 (n14915, n_12805, n14914);
  not g27338 (n_12807, n14913);
  not g27339 (n_12808, n14915);
  and g27340 (n14916, n_12807, n_12808);
  not g27341 (n_12809, n14916);
  and g27342 (n14917, n14652, n_12809);
  not g27343 (n_12810, n14652);
  and g27344 (n14918, n_12810, n14916);
  not g27345 (n_12811, n14918);
  and g27346 (n14919, n14637, n_12811);
  not g27347 (n_12812, n14917);
  and g27348 (n14920, n_12812, n14919);
  not g27349 (n_12813, n14920);
  and g27350 (n14921, n14637, n_12813);
  and g27351 (n14922, n_12811, n_12813);
  and g27352 (n14923, n_12812, n14922);
  not g27353 (n_12814, n14921);
  not g27354 (n_12815, n14923);
  and g27355 (n14924, n_12814, n_12815);
  and g27356 (n14925, n_12450, n_12453);
  and g27357 (n14926, \b[54] , n951);
  and g27358 (n14927, \b[52] , n1056);
  and g27359 (n14928, \b[53] , n946);
  not g27360 (n_12816, n14927);
  not g27361 (n_12817, n14928);
  and g27362 (n14929, n_12816, n_12817);
  not g27363 (n_12818, n14926);
  and g27364 (n14930, n_12818, n14929);
  not g27365 (n_12819, n954);
  and g27366 (n14931, n_12819, n14930);
  not g27367 (n_12820, n9998);
  and g27368 (n14932, n_12820, n14930);
  not g27369 (n_12821, n14931);
  not g27370 (n_12822, n14932);
  and g27371 (n14933, n_12821, n_12822);
  not g27372 (n_12823, n14933);
  and g27373 (n14934, \a[14] , n_12823);
  and g27374 (n14935, n_623, n14933);
  not g27375 (n_12824, n14934);
  not g27376 (n_12825, n14935);
  and g27377 (n14936, n_12824, n_12825);
  not g27378 (n_12826, n14925);
  not g27379 (n_12827, n14936);
  and g27380 (n14937, n_12826, n_12827);
  not g27381 (n_12828, n14937);
  and g27382 (n14938, n_12826, n_12828);
  and g27383 (n14939, n_12827, n_12828);
  not g27384 (n_12829, n14938);
  not g27385 (n_12830, n14939);
  and g27386 (n14940, n_12829, n_12830);
  not g27387 (n_12831, n14924);
  not g27388 (n_12832, n14940);
  and g27389 (n14941, n_12831, n_12832);
  not g27390 (n_12833, n14941);
  and g27391 (n14942, n_12831, n_12833);
  and g27392 (n14943, n_12832, n_12833);
  not g27393 (n_12834, n14942);
  not g27394 (n_12835, n14943);
  and g27395 (n14944, n_12834, n_12835);
  not g27396 (n_12836, n14944);
  and g27397 (n14945, n14622, n_12836);
  not g27398 (n_12837, n14945);
  and g27399 (n14946, n14622, n_12837);
  and g27400 (n14947, n_12836, n_12837);
  not g27401 (n_12838, n14946);
  not g27402 (n_12839, n14947);
  and g27403 (n14948, n_12838, n_12839);
  and g27404 (n14949, \b[60] , n511);
  and g27405 (n14950, \b[58] , n541);
  and g27406 (n14951, \b[59] , n506);
  and g27412 (n14954, n514, n12211);
  not g27415 (n_12844, n14955);
  and g27416 (n14956, \a[8] , n_12844);
  not g27417 (n_12845, n14956);
  and g27418 (n14957, \a[8] , n_12845);
  and g27419 (n14958, n_12844, n_12845);
  not g27420 (n_12846, n14957);
  not g27421 (n_12847, n14958);
  and g27422 (n14959, n_12846, n_12847);
  and g27423 (n14960, n_12474, n_12484);
  not g27424 (n_12848, n14959);
  not g27425 (n_12849, n14960);
  and g27426 (n14961, n_12848, n_12849);
  not g27427 (n_12850, n14961);
  and g27428 (n14962, n_12848, n_12850);
  and g27429 (n14963, n_12849, n_12850);
  not g27430 (n_12851, n14962);
  not g27431 (n_12852, n14963);
  and g27432 (n14964, n_12851, n_12852);
  not g27433 (n_12853, n14948);
  not g27434 (n_12854, n14964);
  and g27435 (n14965, n_12853, n_12854);
  not g27436 (n_12855, n14965);
  and g27437 (n14966, n_12853, n_12855);
  and g27438 (n14967, n_12854, n_12855);
  not g27439 (n_12856, n14966);
  not g27440 (n_12857, n14967);
  and g27441 (n14968, n_12856, n_12857);
  not g27442 (n_12858, n14607);
  not g27443 (n_12859, n14968);
  and g27444 (n14969, n_12858, n_12859);
  not g27445 (n_12860, n14969);
  and g27446 (n14970, n_12858, n_12860);
  and g27447 (n14971, n_12859, n_12860);
  not g27448 (n_12861, n14970);
  not g27449 (n_12862, n14971);
  and g27450 (n14972, n_12861, n_12862);
  and g27451 (n14973, n_12511, n_12514);
  and g27452 (n14974, n14972, n14973);
  not g27453 (n_12863, n14972);
  not g27454 (n_12864, n14973);
  and g27455 (n14975, n_12863, n_12864);
  not g27456 (n_12865, n14974);
  not g27457 (n_12866, n14975);
  and g27458 (n14976, n_12865, n_12866);
  and g27459 (n14977, n_12520, n_12523);
  not g27460 (n_12867, n14977);
  and g27461 (n14978, n14976, n_12867);
  not g27462 (n_12868, n14976);
  and g27463 (n14979, n_12868, n14977);
  not g27464 (n_12869, n14978);
  not g27465 (n_12870, n14979);
  and g27466 (\f[66] , n_12869, n_12870);
  and g27467 (n14981, n_12866, n_12869);
  and g27468 (n14982, n_12535, n_12860);
  and g27469 (n14983, \b[55] , n951);
  and g27470 (n14984, \b[53] , n1056);
  and g27471 (n14985, \b[54] , n946);
  and g27477 (n14988, n954, n10684);
  not g27480 (n_12875, n14989);
  and g27481 (n14990, \a[14] , n_12875);
  not g27482 (n_12876, n14990);
  and g27483 (n14991, \a[14] , n_12876);
  and g27484 (n14992, n_12875, n_12876);
  not g27485 (n_12877, n14991);
  not g27486 (n_12878, n14992);
  and g27487 (n14993, n_12877, n_12878);
  and g27488 (n14994, n_12561, n_12813);
  and g27489 (n14995, n14993, n14994);
  not g27490 (n_12879, n14993);
  not g27491 (n_12880, n14994);
  and g27492 (n14996, n_12879, n_12880);
  not g27493 (n_12881, n14995);
  not g27494 (n_12882, n14996);
  and g27495 (n14997, n_12881, n_12882);
  and g27496 (n14998, \b[49] , n1627);
  and g27497 (n14999, \b[47] , n1763);
  and g27498 (n15000, \b[48] , n1622);
  and g27504 (n15003, n1630, n8625);
  not g27507 (n_12887, n15004);
  and g27508 (n15005, \a[20] , n_12887);
  not g27509 (n_12888, n15005);
  and g27510 (n15006, \a[20] , n_12888);
  and g27511 (n15007, n_12887, n_12888);
  not g27512 (n_12889, n15006);
  not g27513 (n_12890, n15007);
  and g27514 (n15008, n_12889, n_12890);
  and g27515 (n15009, n_12582, n_12583);
  not g27516 (n_12891, n15009);
  and g27517 (n15010, n_12806, n_12891);
  and g27518 (n15011, n15008, n15010);
  not g27519 (n_12892, n15008);
  not g27520 (n_12893, n15010);
  and g27521 (n15012, n_12892, n_12893);
  not g27522 (n_12894, n15011);
  not g27523 (n_12895, n15012);
  and g27524 (n15013, n_12894, n_12895);
  and g27525 (n15014, \b[43] , n2539);
  and g27526 (n15015, \b[41] , n2685);
  and g27527 (n15016, \b[42] , n2534);
  and g27533 (n15019, n2542, n6515);
  not g27536 (n_12900, n15020);
  and g27537 (n15021, \a[26] , n_12900);
  not g27538 (n_12901, n15021);
  and g27539 (n15022, \a[26] , n_12901);
  and g27540 (n15023, n_12900, n_12901);
  not g27541 (n_12902, n15022);
  not g27542 (n_12903, n15023);
  and g27543 (n15024, n_12902, n_12903);
  and g27544 (n15025, n_12610, n_12798);
  and g27545 (n15026, n15024, n15025);
  not g27546 (n_12904, n15024);
  not g27547 (n_12905, n15025);
  and g27548 (n15027, n_12904, n_12905);
  not g27549 (n_12906, n15026);
  not g27550 (n_12907, n15027);
  and g27551 (n15028, n_12906, n_12907);
  and g27552 (n15029, n_12771, n_12774);
  and g27553 (n15030, \b[37] , n3638);
  and g27554 (n15031, \b[35] , n3843);
  and g27555 (n15032, \b[36] , n3633);
  not g27556 (n_12908, n15031);
  not g27557 (n_12909, n15032);
  and g27558 (n15033, n_12908, n_12909);
  not g27559 (n_12910, n15030);
  and g27560 (n15034, n_12910, n15033);
  and g27561 (n15035, n_12780, n15034);
  not g27562 (n_12911, n5181);
  and g27563 (n15036, n_12911, n15034);
  not g27564 (n_12912, n15035);
  not g27565 (n_12913, n15036);
  and g27566 (n15037, n_12912, n_12913);
  not g27567 (n_12914, n15037);
  and g27568 (n15038, \a[32] , n_12914);
  and g27569 (n15039, n_2992, n15037);
  not g27570 (n_12915, n15038);
  not g27571 (n_12916, n15039);
  and g27572 (n15040, n_12915, n_12916);
  not g27573 (n_12917, n15029);
  not g27574 (n_12918, n15040);
  and g27575 (n15041, n_12917, n_12918);
  and g27576 (n15042, n15029, n15040);
  not g27577 (n_12919, n15041);
  not g27578 (n_12920, n15042);
  and g27579 (n15043, n_12919, n_12920);
  and g27580 (n15044, \b[34] , n4287);
  and g27581 (n15045, \b[32] , n4532);
  and g27582 (n15046, \b[33] , n4282);
  and g27588 (n15049, n4290, n4466);
  not g27591 (n_12925, n15050);
  and g27592 (n15051, \a[35] , n_12925);
  not g27593 (n_12926, n15051);
  and g27594 (n15052, \a[35] , n_12926);
  and g27595 (n15053, n_12925, n_12926);
  not g27596 (n_12927, n15052);
  not g27597 (n_12928, n15053);
  and g27598 (n15054, n_12927, n_12928);
  and g27599 (n15055, n_12756, n_12768);
  and g27600 (n15056, \b[16] , n9339);
  and g27601 (n15057, \b[14] , n9732);
  and g27602 (n15058, \b[15] , n9334);
  and g27608 (n15061, n1237, n9342);
  not g27611 (n_12933, n15062);
  and g27612 (n15063, \a[53] , n_12933);
  not g27613 (n_12934, n15063);
  and g27614 (n15064, \a[53] , n_12934);
  and g27615 (n15065, n_12933, n_12934);
  not g27616 (n_12935, n15064);
  not g27617 (n_12936, n15065);
  and g27618 (n15066, n_12935, n_12936);
  and g27619 (n15067, \b[7] , n12668);
  and g27620 (n15068, \b[5] , n13047);
  and g27621 (n15069, \b[6] , n12663);
  and g27627 (n15072, n484, n12671);
  not g27630 (n_12941, n15073);
  and g27631 (n15074, \a[62] , n_12941);
  not g27632 (n_12942, n15074);
  and g27633 (n15075, \a[62] , n_12942);
  and g27634 (n15076, n_12941, n_12942);
  not g27635 (n_12943, n15075);
  not g27636 (n_12944, n15076);
  and g27637 (n15077, n_12943, n_12944);
  and g27638 (n15078, \b[3] , n13903);
  and g27639 (n15079, \b[4] , n_11555);
  not g27640 (n_12945, n15078);
  not g27641 (n_12946, n15079);
  and g27642 (n15080, n_12945, n_12946);
  not g27643 (n_12947, n15080);
  and g27644 (n15081, \a[2] , n_12947);
  not g27645 (n_12948, n15081);
  and g27646 (n15082, \a[2] , n_12948);
  and g27647 (n15083, n_12947, n_12948);
  not g27648 (n_12949, n15082);
  not g27649 (n_12950, n15083);
  and g27650 (n15084, n_12949, n_12950);
  not g27651 (n_12951, n15077);
  not g27652 (n_12952, n15084);
  and g27653 (n15085, n_12951, n_12952);
  not g27654 (n_12953, n15085);
  and g27655 (n15086, n_12951, n_12953);
  and g27656 (n15087, n_12952, n_12953);
  not g27657 (n_12954, n15086);
  not g27658 (n_12955, n15087);
  and g27659 (n15088, n_12954, n_12955);
  and g27660 (n15089, n_12639, n_12653);
  and g27661 (n15090, n15088, n15089);
  not g27662 (n_12956, n15088);
  not g27663 (n_12957, n15089);
  and g27664 (n15091, n_12956, n_12957);
  not g27665 (n_12958, n15090);
  not g27666 (n_12959, n15091);
  and g27667 (n15092, n_12958, n_12959);
  and g27668 (n15093, \b[10] , n11531);
  and g27669 (n15094, \b[8] , n11896);
  and g27670 (n15095, \b[9] , n11526);
  and g27676 (n15098, n738, n11534);
  not g27679 (n_12964, n15099);
  and g27680 (n15100, \a[59] , n_12964);
  not g27681 (n_12965, n15100);
  and g27682 (n15101, \a[59] , n_12965);
  and g27683 (n15102, n_12964, n_12965);
  not g27684 (n_12966, n15101);
  not g27685 (n_12967, n15102);
  and g27686 (n15103, n_12966, n_12967);
  not g27687 (n_12968, n15103);
  and g27688 (n15104, n15092, n_12968);
  not g27689 (n_12969, n15104);
  and g27690 (n15105, n15092, n_12969);
  and g27691 (n15106, n_12968, n_12969);
  not g27692 (n_12970, n15105);
  not g27693 (n_12971, n15106);
  and g27694 (n15107, n_12970, n_12971);
  and g27695 (n15108, n_12657, n_12668);
  and g27696 (n15109, n15107, n15108);
  not g27697 (n_12972, n15107);
  not g27698 (n_12973, n15108);
  and g27699 (n15110, n_12972, n_12973);
  not g27700 (n_12974, n15109);
  not g27701 (n_12975, n15110);
  and g27702 (n15111, n_12974, n_12975);
  and g27703 (n15112, \b[13] , n10426);
  and g27704 (n15113, \b[11] , n10796);
  and g27705 (n15114, \b[12] , n10421);
  and g27711 (n15117, n1008, n10429);
  not g27714 (n_12980, n15118);
  and g27715 (n15119, \a[56] , n_12980);
  not g27716 (n_12981, n15119);
  and g27717 (n15120, \a[56] , n_12981);
  and g27718 (n15121, n_12980, n_12981);
  not g27719 (n_12982, n15120);
  not g27720 (n_12983, n15121);
  and g27721 (n15122, n_12982, n_12983);
  not g27722 (n_12984, n15111);
  and g27723 (n15123, n_12984, n15122);
  not g27724 (n_12985, n15122);
  and g27725 (n15124, n15111, n_12985);
  not g27726 (n_12986, n15123);
  not g27727 (n_12987, n15124);
  and g27728 (n15125, n_12986, n_12987);
  and g27729 (n15126, n_12671, n_12672);
  not g27730 (n_12988, n15126);
  and g27731 (n15127, n_12686, n_12988);
  not g27732 (n_12989, n15127);
  and g27733 (n15128, n15125, n_12989);
  not g27734 (n_12990, n15125);
  and g27735 (n15129, n_12990, n15127);
  not g27736 (n_12991, n15128);
  not g27737 (n_12992, n15129);
  and g27738 (n15130, n_12991, n_12992);
  not g27739 (n_12993, n15066);
  and g27740 (n15131, n_12993, n15130);
  not g27741 (n_12994, n15131);
  and g27742 (n15132, n15130, n_12994);
  and g27743 (n15133, n_12993, n_12994);
  not g27744 (n_12995, n15132);
  not g27745 (n_12996, n15133);
  and g27746 (n15134, n_12995, n_12996);
  and g27747 (n15135, n_12689, n_12692);
  and g27748 (n15136, n15134, n15135);
  not g27749 (n_12997, n15134);
  not g27750 (n_12998, n15135);
  and g27751 (n15137, n_12997, n_12998);
  not g27752 (n_12999, n15136);
  not g27753 (n_13000, n15137);
  and g27754 (n15138, n_12999, n_13000);
  and g27755 (n15139, \b[19] , n8362);
  and g27756 (n15140, \b[17] , n8715);
  and g27757 (n15141, \b[18] , n8357);
  and g27763 (n15144, n1708, n8365);
  not g27766 (n_13005, n15145);
  and g27767 (n15146, \a[50] , n_13005);
  not g27768 (n_13006, n15146);
  and g27769 (n15147, \a[50] , n_13006);
  and g27770 (n15148, n_13005, n_13006);
  not g27771 (n_13007, n15147);
  not g27772 (n_13008, n15148);
  and g27773 (n15149, n_13007, n_13008);
  not g27774 (n_13009, n15149);
  and g27775 (n15150, n15138, n_13009);
  not g27776 (n_13010, n15150);
  and g27777 (n15151, n15138, n_13010);
  and g27778 (n15152, n_13009, n_13010);
  not g27779 (n_13011, n15151);
  not g27780 (n_13012, n15152);
  and g27781 (n15153, n_13011, n_13012);
  and g27782 (n15154, n_12699, n_12709);
  and g27783 (n15155, n15153, n15154);
  not g27784 (n_13013, n15153);
  not g27785 (n_13014, n15154);
  and g27786 (n15156, n_13013, n_13014);
  not g27787 (n_13015, n15155);
  not g27788 (n_13016, n15156);
  and g27789 (n15157, n_13015, n_13016);
  and g27790 (n15158, \b[22] , n7446);
  and g27791 (n15159, \b[20] , n7787);
  and g27792 (n15160, \b[21] , n7441);
  and g27798 (n15163, n2145, n7449);
  not g27801 (n_13021, n15164);
  and g27802 (n15165, \a[47] , n_13021);
  not g27803 (n_13022, n15165);
  and g27804 (n15166, \a[47] , n_13022);
  and g27805 (n15167, n_13021, n_13022);
  not g27806 (n_13023, n15166);
  not g27807 (n_13024, n15167);
  and g27808 (n15168, n_13023, n_13024);
  not g27809 (n_13025, n15168);
  and g27810 (n15169, n15157, n_13025);
  not g27811 (n_13026, n15169);
  and g27812 (n15170, n15157, n_13026);
  and g27813 (n15171, n_13025, n_13026);
  not g27814 (n_13027, n15170);
  not g27815 (n_13028, n15171);
  and g27816 (n15172, n_13027, n_13028);
  and g27817 (n15173, n_12715, n_12727);
  not g27818 (n_13029, n15172);
  not g27819 (n_13030, n15173);
  and g27820 (n15174, n_13029, n_13030);
  not g27821 (n_13031, n15174);
  and g27822 (n15175, n_13029, n_13031);
  and g27823 (n15176, n_13030, n_13031);
  not g27824 (n_13032, n15175);
  not g27825 (n_13033, n15176);
  and g27826 (n15177, n_13032, n_13033);
  and g27827 (n15178, \b[25] , n6595);
  and g27828 (n15179, \b[23] , n6902);
  and g27829 (n15180, \b[24] , n6590);
  and g27835 (n15183, n2485, n6598);
  not g27838 (n_13038, n15184);
  and g27839 (n15185, \a[44] , n_13038);
  not g27840 (n_13039, n15185);
  and g27841 (n15186, \a[44] , n_13039);
  and g27842 (n15187, n_13038, n_13039);
  not g27843 (n_13040, n15186);
  not g27844 (n_13041, n15187);
  and g27845 (n15188, n_13040, n_13041);
  not g27846 (n_13042, n15177);
  not g27847 (n_13043, n15188);
  and g27848 (n15189, n_13042, n_13043);
  not g27849 (n_13044, n15189);
  and g27850 (n15190, n_13042, n_13044);
  and g27851 (n15191, n_13043, n_13044);
  not g27852 (n_13045, n15190);
  not g27853 (n_13046, n15191);
  and g27854 (n15192, n_13045, n_13046);
  and g27855 (n15193, n_12731, n_12734);
  and g27856 (n15194, n15192, n15193);
  not g27857 (n_13047, n15192);
  not g27858 (n_13048, n15193);
  and g27859 (n15195, n_13047, n_13048);
  not g27860 (n_13049, n15194);
  not g27861 (n_13050, n15195);
  and g27862 (n15196, n_13049, n_13050);
  and g27863 (n15197, \b[28] , n5777);
  and g27864 (n15198, \b[26] , n6059);
  and g27865 (n15199, \b[27] , n5772);
  and g27871 (n15202, n3189, n5780);
  not g27874 (n_13055, n15203);
  and g27875 (n15204, \a[41] , n_13055);
  not g27876 (n_13056, n15204);
  and g27877 (n15205, \a[41] , n_13056);
  and g27878 (n15206, n_13055, n_13056);
  not g27879 (n_13057, n15205);
  not g27880 (n_13058, n15206);
  and g27881 (n15207, n_13057, n_13058);
  not g27882 (n_13059, n15207);
  and g27883 (n15208, n15196, n_13059);
  not g27884 (n_13060, n15208);
  and g27885 (n15209, n15196, n_13060);
  and g27886 (n15210, n_13059, n_13060);
  not g27887 (n_13061, n15209);
  not g27888 (n_13062, n15210);
  and g27889 (n15211, n_13061, n_13062);
  and g27890 (n15212, n_12740, n_12750);
  and g27891 (n15213, n15211, n15212);
  not g27892 (n_13063, n15211);
  not g27893 (n_13064, n15212);
  and g27894 (n15214, n_13063, n_13064);
  not g27895 (n_13065, n15213);
  not g27896 (n_13066, n15214);
  and g27897 (n15215, n_13065, n_13066);
  and g27898 (n15216, \b[31] , n5035);
  and g27899 (n15217, \b[29] , n5277);
  and g27900 (n15218, \b[30] , n5030);
  and g27906 (n15221, n3796, n5038);
  not g27909 (n_13071, n15222);
  and g27910 (n15223, \a[38] , n_13071);
  not g27911 (n_13072, n15223);
  and g27912 (n15224, \a[38] , n_13072);
  and g27913 (n15225, n_13071, n_13072);
  not g27914 (n_13073, n15224);
  not g27915 (n_13074, n15225);
  and g27916 (n15226, n_13073, n_13074);
  not g27917 (n_13075, n15215);
  and g27918 (n15227, n_13075, n15226);
  not g27919 (n_13076, n15226);
  and g27920 (n15228, n15215, n_13076);
  not g27921 (n_13077, n15227);
  not g27922 (n_13078, n15228);
  and g27923 (n15229, n_13077, n_13078);
  not g27924 (n_13079, n15055);
  and g27925 (n15230, n_13079, n15229);
  not g27926 (n_13080, n15230);
  and g27927 (n15231, n_13079, n_13080);
  and g27928 (n15232, n15229, n_13080);
  not g27929 (n_13081, n15231);
  not g27930 (n_13082, n15232);
  and g27931 (n15233, n_13081, n_13082);
  not g27932 (n_13083, n15054);
  not g27933 (n_13084, n15233);
  and g27934 (n15234, n_13083, n_13084);
  not g27935 (n_13085, n15234);
  and g27936 (n15235, n_13083, n_13085);
  and g27937 (n15236, n_13084, n_13085);
  not g27938 (n_13086, n15235);
  not g27939 (n_13087, n15236);
  and g27940 (n15237, n_13086, n_13087);
  not g27941 (n_13088, n15043);
  and g27942 (n15238, n_13088, n15237);
  not g27943 (n_13089, n15237);
  and g27944 (n15239, n15043, n_13089);
  not g27945 (n_13090, n15238);
  not g27946 (n_13091, n15239);
  and g27947 (n15240, n_13090, n_13091);
  and g27948 (n15241, n_12789, n_12794);
  and g27949 (n15242, \b[40] , n3050);
  and g27950 (n15243, \b[38] , n3243);
  and g27951 (n15244, \b[39] , n3045);
  not g27952 (n_13092, n15243);
  not g27953 (n_13093, n15244);
  and g27954 (n15245, n_13092, n_13093);
  not g27955 (n_13094, n15242);
  and g27956 (n15246, n_13094, n15245);
  and g27957 (n15247, n_12601, n15246);
  not g27958 (n_13095, n5955);
  and g27959 (n15248, n_13095, n15246);
  not g27960 (n_13096, n15247);
  not g27961 (n_13097, n15248);
  and g27962 (n15249, n_13096, n_13097);
  not g27963 (n_13098, n15249);
  and g27964 (n15250, \a[29] , n_13098);
  and g27965 (n15251, n_2476, n15249);
  not g27966 (n_13099, n15250);
  not g27967 (n_13100, n15251);
  and g27968 (n15252, n_13099, n_13100);
  not g27969 (n_13101, n15241);
  not g27970 (n_13102, n15252);
  and g27971 (n15253, n_13101, n_13102);
  not g27972 (n_13103, n15253);
  and g27973 (n15254, n_13101, n_13103);
  and g27974 (n15255, n_13102, n_13103);
  not g27975 (n_13104, n15254);
  not g27976 (n_13105, n15255);
  and g27977 (n15256, n_13104, n_13105);
  not g27978 (n_13106, n15256);
  and g27979 (n15257, n15240, n_13106);
  not g27980 (n_13107, n15257);
  and g27981 (n15258, n15240, n_13107);
  and g27982 (n15259, n_13106, n_13107);
  not g27983 (n_13108, n15258);
  not g27984 (n_13109, n15259);
  and g27985 (n15260, n_13108, n_13109);
  not g27986 (n_13110, n15260);
  and g27987 (n15261, n15028, n_13110);
  not g27988 (n_13111, n15261);
  and g27989 (n15262, n15028, n_13111);
  and g27990 (n15263, n_13110, n_13111);
  not g27991 (n_13112, n15262);
  not g27992 (n_13113, n15263);
  and g27993 (n15264, n_13112, n_13113);
  and g27994 (n15265, \b[46] , n2048);
  and g27995 (n15266, \b[44] , n2198);
  and g27996 (n15267, \b[45] , n2043);
  and g28002 (n15270, n2051, n7677);
  not g28005 (n_13118, n15271);
  and g28006 (n15272, \a[23] , n_13118);
  not g28007 (n_13119, n15272);
  and g28008 (n15273, \a[23] , n_13119);
  and g28009 (n15274, n_13118, n_13119);
  not g28010 (n_13120, n15273);
  not g28011 (n_13121, n15274);
  and g28012 (n15275, n_13120, n_13121);
  and g28013 (n15276, n_12597, n_12805);
  not g28014 (n_13122, n15275);
  not g28015 (n_13123, n15276);
  and g28016 (n15277, n_13122, n_13123);
  not g28017 (n_13124, n15277);
  and g28018 (n15278, n_13122, n_13124);
  and g28019 (n15279, n_13123, n_13124);
  not g28020 (n_13125, n15278);
  not g28021 (n_13126, n15279);
  and g28022 (n15280, n_13125, n_13126);
  not g28023 (n_13127, n15264);
  and g28024 (n15281, n_13127, n15280);
  not g28025 (n_13128, n15280);
  and g28026 (n15282, n15264, n_13128);
  not g28027 (n_13129, n15281);
  not g28028 (n_13130, n15282);
  and g28029 (n15283, n_13129, n_13130);
  not g28030 (n_13131, n15283);
  and g28031 (n15284, n15013, n_13131);
  not g28032 (n_13132, n15284);
  and g28033 (n15285, n15013, n_13132);
  and g28034 (n15286, n_13131, n_13132);
  not g28035 (n_13133, n15285);
  not g28036 (n_13134, n15286);
  and g28037 (n15287, n_13133, n_13134);
  and g28038 (n15288, \b[52] , n1302);
  and g28039 (n15289, \b[50] , n1391);
  and g28040 (n15290, \b[51] , n1297);
  and g28046 (n15293, n1305, n9628);
  not g28049 (n_13139, n15294);
  and g28050 (n15295, \a[17] , n_13139);
  not g28051 (n_13140, n15295);
  and g28052 (n15296, \a[17] , n_13140);
  and g28053 (n15297, n_13139, n_13140);
  not g28054 (n_13141, n15296);
  not g28055 (n_13142, n15297);
  and g28056 (n15298, n_13141, n_13142);
  and g28057 (n15299, n_12573, n_12812);
  not g28058 (n_13143, n15298);
  not g28059 (n_13144, n15299);
  and g28060 (n15300, n_13143, n_13144);
  not g28061 (n_13145, n15300);
  and g28062 (n15301, n_13143, n_13145);
  and g28063 (n15302, n_13144, n_13145);
  not g28064 (n_13146, n15301);
  not g28065 (n_13147, n15302);
  and g28066 (n15303, n_13146, n_13147);
  not g28067 (n_13148, n15287);
  and g28068 (n15304, n_13148, n15303);
  not g28069 (n_13149, n15303);
  and g28070 (n15305, n15287, n_13149);
  not g28071 (n_13150, n15304);
  not g28072 (n_13151, n15305);
  and g28073 (n15306, n_13150, n_13151);
  not g28074 (n_13152, n15306);
  and g28075 (n15307, n14997, n_13152);
  not g28076 (n_13153, n15307);
  and g28077 (n15308, n14997, n_13153);
  and g28078 (n15309, n_13152, n_13153);
  not g28079 (n_13154, n15308);
  not g28080 (n_13155, n15309);
  and g28081 (n15310, n_13154, n_13155);
  and g28082 (n15311, n_12828, n_12833);
  and g28083 (n15312, \b[58] , n700);
  and g28084 (n15313, \b[56] , n767);
  and g28085 (n15314, \b[57] , n695);
  not g28086 (n_13156, n15313);
  not g28087 (n_13157, n15314);
  and g28088 (n15315, n_13156, n_13157);
  not g28089 (n_13158, n15312);
  and g28090 (n15316, n_13158, n15315);
  not g28091 (n_13159, n703);
  and g28092 (n15317, n_13159, n15316);
  not g28093 (n_13160, n11436);
  and g28094 (n15318, n_13160, n15316);
  not g28095 (n_13161, n15317);
  not g28096 (n_13162, n15318);
  and g28097 (n15319, n_13161, n_13162);
  not g28098 (n_13163, n15319);
  and g28099 (n15320, \a[11] , n_13163);
  and g28100 (n15321, n_400, n15319);
  not g28101 (n_13164, n15320);
  not g28102 (n_13165, n15321);
  and g28103 (n15322, n_13164, n_13165);
  not g28104 (n_13166, n15311);
  not g28105 (n_13167, n15322);
  and g28106 (n15323, n_13166, n_13167);
  not g28107 (n_13168, n15323);
  and g28108 (n15324, n_13166, n_13168);
  and g28109 (n15325, n_13167, n_13168);
  not g28110 (n_13169, n15324);
  not g28111 (n_13170, n15325);
  and g28112 (n15326, n_13169, n_13170);
  not g28113 (n_13171, n15310);
  not g28114 (n_13172, n15326);
  and g28115 (n15327, n_13171, n_13172);
  not g28116 (n_13173, n15327);
  and g28117 (n15328, n_13171, n_13173);
  and g28118 (n15329, n_13172, n_13173);
  not g28119 (n_13174, n15328);
  not g28120 (n_13175, n15329);
  and g28121 (n15330, n_13174, n_13175);
  and g28122 (n15331, n_12549, n_12837);
  and g28123 (n15332, \b[61] , n511);
  and g28124 (n15333, \b[59] , n541);
  and g28125 (n15334, \b[60] , n506);
  not g28126 (n_13176, n15333);
  not g28127 (n_13177, n15334);
  and g28128 (n15335, n_13176, n_13177);
  not g28129 (n_13178, n15332);
  and g28130 (n15336, n_13178, n15335);
  not g28131 (n_13179, n514);
  and g28132 (n15337, n_13179, n15336);
  not g28133 (n_13180, n12969);
  and g28134 (n15338, n_13180, n15336);
  not g28135 (n_13181, n15337);
  not g28136 (n_13182, n15338);
  and g28137 (n15339, n_13181, n_13182);
  not g28138 (n_13183, n15339);
  and g28139 (n15340, \a[8] , n_13183);
  and g28140 (n15341, n_234, n15339);
  not g28141 (n_13184, n15340);
  not g28142 (n_13185, n15341);
  and g28143 (n15342, n_13184, n_13185);
  not g28144 (n_13186, n15331);
  not g28145 (n_13187, n15342);
  and g28146 (n15343, n_13186, n_13187);
  not g28147 (n_13188, n15343);
  and g28148 (n15344, n_13186, n_13188);
  and g28149 (n15345, n_13187, n_13188);
  not g28150 (n_13189, n15344);
  not g28151 (n_13190, n15345);
  and g28152 (n15346, n_13189, n_13190);
  not g28153 (n_13191, n15330);
  not g28154 (n_13192, n15346);
  and g28155 (n15347, n_13191, n_13192);
  not g28156 (n_13193, n15347);
  and g28157 (n15348, n_13191, n_13193);
  and g28158 (n15349, n_13192, n_13193);
  not g28159 (n_13194, n15348);
  not g28160 (n_13195, n15349);
  and g28161 (n15350, n_13194, n_13195);
  and g28162 (n15351, n_12850, n_12855);
  and g28163 (n15352, \b[62] , n403);
  and g28164 (n15353, \b[63] , n357);
  not g28165 (n_13196, n15352);
  not g28166 (n_13197, n15353);
  and g28167 (n15354, n_13196, n_13197);
  and g28168 (n15355, n_141, n15354);
  and g28169 (n15356, n13800, n15354);
  not g28170 (n_13198, n15355);
  not g28171 (n_13199, n15356);
  and g28172 (n15357, n_13198, n_13199);
  not g28173 (n_13200, n15357);
  and g28174 (n15358, \a[5] , n_13200);
  and g28175 (n15359, n_99, n15357);
  not g28176 (n_13201, n15358);
  not g28177 (n_13202, n15359);
  and g28178 (n15360, n_13201, n_13202);
  not g28179 (n_13203, n15351);
  not g28180 (n_13204, n15360);
  and g28181 (n15361, n_13203, n_13204);
  not g28182 (n_13205, n15361);
  and g28183 (n15362, n_13203, n_13205);
  and g28184 (n15363, n_13204, n_13205);
  not g28185 (n_13206, n15362);
  not g28186 (n_13207, n15363);
  and g28187 (n15364, n_13206, n_13207);
  not g28188 (n_13208, n15350);
  not g28189 (n_13209, n15364);
  and g28190 (n15365, n_13208, n_13209);
  and g28191 (n15366, n15350, n_13207);
  and g28192 (n15367, n_13206, n15366);
  not g28193 (n_13210, n15365);
  not g28194 (n_13211, n15367);
  and g28195 (n15368, n_13210, n_13211);
  not g28196 (n_13212, n14982);
  and g28197 (n15369, n_13212, n15368);
  not g28198 (n_13213, n15369);
  and g28199 (n15370, n_13212, n_13213);
  and g28200 (n15371, n15368, n_13213);
  not g28201 (n_13214, n15370);
  not g28202 (n_13215, n15371);
  and g28203 (n15372, n_13214, n_13215);
  not g28204 (n_13216, n14981);
  not g28205 (n_13217, n15372);
  and g28206 (n15373, n_13216, n_13217);
  and g28207 (n15374, n14981, n_13215);
  and g28208 (n15375, n_13214, n15374);
  not g28209 (n_13218, n15373);
  not g28210 (n_13219, n15375);
  and g28211 (\f[67] , n_13218, n_13219);
  and g28212 (n15377, n_13213, n_13218);
  and g28213 (n15378, n_13205, n_13210);
  and g28214 (n15379, n_13188, n_13193);
  and g28215 (n15380, \b[63] , n403);
  and g28216 (n15381, n365, n13797);
  not g28217 (n_13220, n15380);
  not g28218 (n_13221, n15381);
  and g28219 (n15382, n_13220, n_13221);
  not g28220 (n_13222, n15382);
  and g28221 (n15383, \a[5] , n_13222);
  not g28222 (n_13223, n15383);
  and g28223 (n15384, \a[5] , n_13223);
  and g28224 (n15385, n_13222, n_13223);
  not g28225 (n_13224, n15384);
  not g28226 (n_13225, n15385);
  and g28227 (n15386, n_13224, n_13225);
  not g28228 (n_13226, n15379);
  not g28229 (n_13227, n15386);
  and g28230 (n15387, n_13226, n_13227);
  not g28231 (n_13228, n15387);
  and g28232 (n15388, n_13226, n_13228);
  and g28233 (n15389, n_13227, n_13228);
  not g28234 (n_13229, n15388);
  not g28235 (n_13230, n15389);
  and g28236 (n15390, n_13229, n_13230);
  and g28237 (n15391, \b[59] , n700);
  and g28238 (n15392, \b[57] , n767);
  and g28239 (n15393, \b[58] , n695);
  and g28245 (n15396, n703, n12179);
  not g28248 (n_13235, n15397);
  and g28249 (n15398, \a[11] , n_13235);
  not g28250 (n_13236, n15398);
  and g28251 (n15399, \a[11] , n_13236);
  and g28252 (n15400, n_13235, n_13236);
  not g28253 (n_13237, n15399);
  not g28254 (n_13238, n15400);
  and g28255 (n15401, n_13237, n_13238);
  and g28256 (n15402, n_12882, n_13153);
  and g28257 (n15403, n15401, n15402);
  not g28258 (n_13239, n15401);
  not g28259 (n_13240, n15402);
  and g28260 (n15404, n_13239, n_13240);
  not g28261 (n_13241, n15403);
  not g28262 (n_13242, n15404);
  and g28263 (n15405, n_13241, n_13242);
  and g28264 (n15406, \b[56] , n951);
  and g28265 (n15407, \b[54] , n1056);
  and g28266 (n15408, \b[55] , n946);
  and g28272 (n15411, n954, n10708);
  not g28275 (n_13247, n15412);
  and g28276 (n15413, \a[14] , n_13247);
  not g28277 (n_13248, n15413);
  and g28278 (n15414, \a[14] , n_13248);
  and g28279 (n15415, n_13247, n_13248);
  not g28280 (n_13249, n15414);
  not g28281 (n_13250, n15415);
  and g28282 (n15416, n_13249, n_13250);
  and g28283 (n15417, n_13148, n_13149);
  not g28284 (n_13251, n15417);
  and g28285 (n15418, n_13145, n_13251);
  not g28286 (n_13252, n15416);
  not g28287 (n_13253, n15418);
  and g28288 (n15419, n_13252, n_13253);
  not g28289 (n_13254, n15419);
  and g28290 (n15420, n_13252, n_13254);
  and g28291 (n15421, n_13253, n_13254);
  not g28292 (n_13255, n15420);
  not g28293 (n_13256, n15421);
  and g28294 (n15422, n_13255, n_13256);
  and g28295 (n15423, n_12895, n_13132);
  and g28296 (n15424, \b[53] , n1302);
  and g28297 (n15425, \b[51] , n1391);
  and g28298 (n15426, \b[52] , n1297);
  not g28299 (n_13257, n15425);
  not g28300 (n_13258, n15426);
  and g28301 (n15427, n_13257, n_13258);
  not g28302 (n_13259, n15424);
  and g28303 (n15428, n_13259, n15427);
  not g28304 (n_13260, n1305);
  and g28305 (n15429, n_13260, n15428);
  not g28306 (n_13261, n9972);
  and g28307 (n15430, n_13261, n15428);
  not g28308 (n_13262, n15429);
  not g28309 (n_13263, n15430);
  and g28310 (n15431, n_13262, n_13263);
  not g28311 (n_13264, n15431);
  and g28312 (n15432, \a[17] , n_13264);
  and g28313 (n15433, n_926, n15431);
  not g28314 (n_13265, n15432);
  not g28315 (n_13266, n15433);
  and g28316 (n15434, n_13265, n_13266);
  not g28317 (n_13267, n15423);
  not g28318 (n_13268, n15434);
  and g28319 (n15435, n_13267, n_13268);
  and g28320 (n15436, n15423, n15434);
  not g28321 (n_13269, n15435);
  not g28322 (n_13270, n15436);
  and g28323 (n15437, n_13269, n_13270);
  and g28324 (n15438, \b[50] , n1627);
  and g28325 (n15439, \b[48] , n1763);
  and g28326 (n15440, \b[49] , n1622);
  and g28332 (n15443, n1630, n8949);
  not g28335 (n_13275, n15444);
  and g28336 (n15445, \a[20] , n_13275);
  not g28337 (n_13276, n15445);
  and g28338 (n15446, \a[20] , n_13276);
  and g28339 (n15447, n_13275, n_13276);
  not g28340 (n_13277, n15446);
  not g28341 (n_13278, n15447);
  and g28342 (n15448, n_13277, n_13278);
  and g28343 (n15449, n_13127, n_13128);
  not g28344 (n_13279, n15449);
  and g28345 (n15450, n_13124, n_13279);
  not g28346 (n_13280, n15448);
  not g28347 (n_13281, n15450);
  and g28348 (n15451, n_13280, n_13281);
  not g28349 (n_13282, n15451);
  and g28350 (n15452, n_13280, n_13282);
  and g28351 (n15453, n_13281, n_13282);
  not g28352 (n_13283, n15452);
  not g28353 (n_13284, n15453);
  and g28354 (n15454, n_13283, n_13284);
  and g28355 (n15455, \b[47] , n2048);
  and g28356 (n15456, \b[45] , n2198);
  and g28357 (n15457, \b[46] , n2043);
  and g28363 (n15460, n2051, n7703);
  not g28366 (n_13289, n15461);
  and g28367 (n15462, \a[23] , n_13289);
  not g28368 (n_13290, n15462);
  and g28369 (n15463, \a[23] , n_13290);
  and g28370 (n15464, n_13289, n_13290);
  not g28371 (n_13291, n15463);
  not g28372 (n_13292, n15464);
  and g28373 (n15465, n_13291, n_13292);
  and g28374 (n15466, n_12907, n_13111);
  and g28375 (n15467, n15465, n15466);
  not g28376 (n_13293, n15465);
  not g28377 (n_13294, n15466);
  and g28378 (n15468, n_13293, n_13294);
  not g28379 (n_13295, n15467);
  not g28380 (n_13296, n15468);
  and g28381 (n15469, n_13295, n_13296);
  and g28382 (n15470, \b[41] , n3050);
  and g28383 (n15471, \b[39] , n3243);
  and g28384 (n15472, \b[40] , n3045);
  and g28390 (n15475, n3053, n6219);
  not g28393 (n_13301, n15476);
  and g28394 (n15477, \a[29] , n_13301);
  not g28395 (n_13302, n15477);
  and g28396 (n15478, \a[29] , n_13302);
  and g28397 (n15479, n_13301, n_13302);
  not g28398 (n_13303, n15478);
  not g28399 (n_13304, n15479);
  and g28400 (n15480, n_13303, n_13304);
  and g28401 (n15481, n_12919, n_13091);
  and g28402 (n15482, n15480, n15481);
  not g28403 (n_13305, n15480);
  not g28404 (n_13306, n15481);
  and g28405 (n15483, n_13305, n_13306);
  not g28406 (n_13307, n15482);
  not g28407 (n_13308, n15483);
  and g28408 (n15484, n_13307, n_13308);
  and g28409 (n15485, \b[35] , n4287);
  and g28410 (n15486, \b[33] , n4532);
  and g28411 (n15487, \b[34] , n4282);
  and g28417 (n15490, n4290, n4696);
  not g28420 (n_13313, n15491);
  and g28421 (n15492, \a[35] , n_13313);
  not g28422 (n_13314, n15492);
  and g28423 (n15493, \a[35] , n_13314);
  and g28424 (n15494, n_13313, n_13314);
  not g28425 (n_13315, n15493);
  not g28426 (n_13316, n15494);
  and g28427 (n15495, n_13315, n_13316);
  and g28428 (n15496, \b[23] , n7446);
  and g28429 (n15497, \b[21] , n7787);
  and g28430 (n15498, \b[22] , n7441);
  and g28436 (n15501, n2300, n7449);
  not g28439 (n_13321, n15502);
  and g28440 (n15503, \a[47] , n_13321);
  not g28441 (n_13322, n15503);
  and g28442 (n15504, \a[47] , n_13322);
  and g28443 (n15505, n_13321, n_13322);
  not g28444 (n_13323, n15504);
  not g28445 (n_13324, n15505);
  and g28446 (n15506, n_13323, n_13324);
  and g28447 (n15507, \b[14] , n10426);
  and g28448 (n15508, \b[12] , n10796);
  and g28449 (n15509, \b[13] , n10421);
  and g28455 (n15512, n1034, n10429);
  not g28458 (n_13329, n15513);
  and g28459 (n15514, \a[56] , n_13329);
  not g28460 (n_13330, n15514);
  and g28461 (n15515, \a[56] , n_13330);
  and g28462 (n15516, n_13329, n_13330);
  not g28463 (n_13331, n15515);
  not g28464 (n_13332, n15516);
  and g28465 (n15517, n_13331, n_13332);
  and g28466 (n15518, \b[8] , n12668);
  and g28467 (n15519, \b[6] , n13047);
  and g28468 (n15520, \b[7] , n12663);
  and g28474 (n15523, n585, n12671);
  not g28477 (n_13337, n15524);
  and g28478 (n15525, \a[62] , n_13337);
  not g28479 (n_13338, n15525);
  and g28480 (n15526, \a[62] , n_13338);
  and g28481 (n15527, n_13337, n_13338);
  not g28482 (n_13339, n15526);
  not g28483 (n_13340, n15527);
  and g28484 (n15528, n_13339, n_13340);
  and g28485 (n15529, \b[4] , n13903);
  and g28486 (n15530, \b[5] , n_11555);
  not g28487 (n_13341, n15529);
  not g28488 (n_13342, n15530);
  and g28489 (n15531, n_13341, n_13342);
  not g28490 (n_13343, n15531);
  and g28491 (n15532, \a[2] , n_13343);
  not g28492 (n_13344, n15532);
  and g28493 (n15533, \a[2] , n_13344);
  and g28494 (n15534, n_13343, n_13344);
  not g28495 (n_13345, n15533);
  not g28496 (n_13346, n15534);
  and g28497 (n15535, n_13345, n_13346);
  not g28498 (n_13347, n15528);
  not g28499 (n_13348, n15535);
  and g28500 (n15536, n_13347, n_13348);
  not g28501 (n_13349, n15536);
  and g28502 (n15537, n_13347, n_13349);
  and g28503 (n15538, n_13348, n_13349);
  not g28504 (n_13350, n15537);
  not g28505 (n_13351, n15538);
  and g28506 (n15539, n_13350, n_13351);
  and g28507 (n15540, n_12948, n_12953);
  and g28508 (n15541, n15539, n15540);
  not g28509 (n_13352, n15539);
  not g28510 (n_13353, n15540);
  and g28511 (n15542, n_13352, n_13353);
  not g28512 (n_13354, n15541);
  not g28513 (n_13355, n15542);
  and g28514 (n15543, n_13354, n_13355);
  and g28515 (n15544, \b[11] , n11531);
  and g28516 (n15545, \b[9] , n11896);
  and g28517 (n15546, \b[10] , n11526);
  and g28523 (n15549, n818, n11534);
  not g28526 (n_13360, n15550);
  and g28527 (n15551, \a[59] , n_13360);
  not g28528 (n_13361, n15551);
  and g28529 (n15552, \a[59] , n_13361);
  and g28530 (n15553, n_13360, n_13361);
  not g28531 (n_13362, n15552);
  not g28532 (n_13363, n15553);
  and g28533 (n15554, n_13362, n_13363);
  not g28534 (n_13364, n15543);
  and g28535 (n15555, n_13364, n15554);
  not g28536 (n_13365, n15554);
  and g28537 (n15556, n15543, n_13365);
  not g28538 (n_13366, n15555);
  not g28539 (n_13367, n15556);
  and g28540 (n15557, n_13366, n_13367);
  and g28541 (n15558, n_12959, n_12969);
  not g28542 (n_13368, n15558);
  and g28543 (n15559, n15557, n_13368);
  not g28544 (n_13369, n15557);
  and g28545 (n15560, n_13369, n15558);
  not g28546 (n_13370, n15559);
  not g28547 (n_13371, n15560);
  and g28548 (n15561, n_13370, n_13371);
  not g28549 (n_13372, n15517);
  and g28550 (n15562, n_13372, n15561);
  not g28551 (n_13373, n15562);
  and g28552 (n15563, n15561, n_13373);
  and g28553 (n15564, n_13372, n_13373);
  not g28554 (n_13374, n15563);
  not g28555 (n_13375, n15564);
  and g28556 (n15565, n_13374, n_13375);
  and g28557 (n15566, n_12975, n_12987);
  not g28558 (n_13376, n15565);
  not g28559 (n_13377, n15566);
  and g28560 (n15567, n_13376, n_13377);
  not g28561 (n_13378, n15567);
  and g28562 (n15568, n_13376, n_13378);
  and g28563 (n15569, n_13377, n_13378);
  not g28564 (n_13379, n15568);
  not g28565 (n_13380, n15569);
  and g28566 (n15570, n_13379, n_13380);
  and g28567 (n15571, \b[17] , n9339);
  and g28568 (n15572, \b[15] , n9732);
  and g28569 (n15573, \b[16] , n9334);
  and g28575 (n15576, n1356, n9342);
  not g28578 (n_13385, n15577);
  and g28579 (n15578, \a[53] , n_13385);
  not g28580 (n_13386, n15578);
  and g28581 (n15579, \a[53] , n_13386);
  and g28582 (n15580, n_13385, n_13386);
  not g28583 (n_13387, n15579);
  not g28584 (n_13388, n15580);
  and g28585 (n15581, n_13387, n_13388);
  not g28586 (n_13389, n15570);
  not g28587 (n_13390, n15581);
  and g28588 (n15582, n_13389, n_13390);
  not g28589 (n_13391, n15582);
  and g28590 (n15583, n_13389, n_13391);
  and g28591 (n15584, n_13390, n_13391);
  not g28592 (n_13392, n15583);
  not g28593 (n_13393, n15584);
  and g28594 (n15585, n_13392, n_13393);
  and g28595 (n15586, n_12991, n_12994);
  and g28596 (n15587, n15585, n15586);
  not g28597 (n_13394, n15585);
  not g28598 (n_13395, n15586);
  and g28599 (n15588, n_13394, n_13395);
  not g28600 (n_13396, n15587);
  not g28601 (n_13397, n15588);
  and g28602 (n15589, n_13396, n_13397);
  and g28603 (n15590, \b[20] , n8362);
  and g28604 (n15591, \b[18] , n8715);
  and g28605 (n15592, \b[19] , n8357);
  and g28611 (n15595, n1846, n8365);
  not g28614 (n_13402, n15596);
  and g28615 (n15597, \a[50] , n_13402);
  not g28616 (n_13403, n15597);
  and g28617 (n15598, \a[50] , n_13403);
  and g28618 (n15599, n_13402, n_13403);
  not g28619 (n_13404, n15598);
  not g28620 (n_13405, n15599);
  and g28621 (n15600, n_13404, n_13405);
  not g28622 (n_13406, n15589);
  and g28623 (n15601, n_13406, n15600);
  not g28624 (n_13407, n15600);
  and g28625 (n15602, n15589, n_13407);
  not g28626 (n_13408, n15601);
  not g28627 (n_13409, n15602);
  and g28628 (n15603, n_13408, n_13409);
  and g28629 (n15604, n_13000, n_13010);
  not g28630 (n_13410, n15604);
  and g28631 (n15605, n15603, n_13410);
  not g28632 (n_13411, n15603);
  and g28633 (n15606, n_13411, n15604);
  not g28634 (n_13412, n15605);
  not g28635 (n_13413, n15606);
  and g28636 (n15607, n_13412, n_13413);
  not g28637 (n_13414, n15506);
  and g28638 (n15608, n_13414, n15607);
  not g28639 (n_13415, n15608);
  and g28640 (n15609, n15607, n_13415);
  and g28641 (n15610, n_13414, n_13415);
  not g28642 (n_13416, n15609);
  not g28643 (n_13417, n15610);
  and g28644 (n15611, n_13416, n_13417);
  and g28645 (n15612, n_13016, n_13026);
  and g28646 (n15613, n15611, n15612);
  not g28647 (n_13418, n15611);
  not g28648 (n_13419, n15612);
  and g28649 (n15614, n_13418, n_13419);
  not g28650 (n_13420, n15613);
  not g28651 (n_13421, n15614);
  and g28652 (n15615, n_13420, n_13421);
  and g28653 (n15616, \b[26] , n6595);
  and g28654 (n15617, \b[24] , n6902);
  and g28655 (n15618, \b[25] , n6590);
  and g28661 (n15621, n2813, n6598);
  not g28664 (n_13426, n15622);
  and g28665 (n15623, \a[44] , n_13426);
  not g28666 (n_13427, n15623);
  and g28667 (n15624, \a[44] , n_13427);
  and g28668 (n15625, n_13426, n_13427);
  not g28669 (n_13428, n15624);
  not g28670 (n_13429, n15625);
  and g28671 (n15626, n_13428, n_13429);
  not g28672 (n_13430, n15626);
  and g28673 (n15627, n15615, n_13430);
  not g28674 (n_13431, n15627);
  and g28675 (n15628, n15615, n_13431);
  and g28676 (n15629, n_13430, n_13431);
  not g28677 (n_13432, n15628);
  not g28678 (n_13433, n15629);
  and g28679 (n15630, n_13432, n_13433);
  and g28680 (n15631, n_13031, n_13044);
  and g28681 (n15632, n15630, n15631);
  not g28682 (n_13434, n15630);
  not g28683 (n_13435, n15631);
  and g28684 (n15633, n_13434, n_13435);
  not g28685 (n_13436, n15632);
  not g28686 (n_13437, n15633);
  and g28687 (n15634, n_13436, n_13437);
  and g28688 (n15635, \b[29] , n5777);
  and g28689 (n15636, \b[27] , n6059);
  and g28690 (n15637, \b[28] , n5772);
  and g28696 (n15640, n3383, n5780);
  not g28699 (n_13442, n15641);
  and g28700 (n15642, \a[41] , n_13442);
  not g28701 (n_13443, n15642);
  and g28702 (n15643, \a[41] , n_13443);
  and g28703 (n15644, n_13442, n_13443);
  not g28704 (n_13444, n15643);
  not g28705 (n_13445, n15644);
  and g28706 (n15645, n_13444, n_13445);
  not g28707 (n_13446, n15645);
  and g28708 (n15646, n15634, n_13446);
  not g28709 (n_13447, n15646);
  and g28710 (n15647, n15634, n_13447);
  and g28711 (n15648, n_13446, n_13447);
  not g28712 (n_13448, n15647);
  not g28713 (n_13449, n15648);
  and g28714 (n15649, n_13448, n_13449);
  and g28715 (n15650, n_13050, n_13060);
  and g28716 (n15651, n15649, n15650);
  not g28717 (n_13450, n15649);
  not g28718 (n_13451, n15650);
  and g28719 (n15652, n_13450, n_13451);
  not g28720 (n_13452, n15651);
  not g28721 (n_13453, n15652);
  and g28722 (n15653, n_13452, n_13453);
  and g28723 (n15654, \b[32] , n5035);
  and g28724 (n15655, \b[30] , n5277);
  and g28725 (n15656, \b[31] , n5030);
  and g28731 (n15659, n4013, n5038);
  not g28734 (n_13458, n15660);
  and g28735 (n15661, \a[38] , n_13458);
  not g28736 (n_13459, n15661);
  and g28737 (n15662, \a[38] , n_13459);
  and g28738 (n15663, n_13458, n_13459);
  not g28739 (n_13460, n15662);
  not g28740 (n_13461, n15663);
  and g28741 (n15664, n_13460, n_13461);
  not g28742 (n_13462, n15653);
  and g28743 (n15665, n_13462, n15664);
  not g28744 (n_13463, n15664);
  and g28745 (n15666, n15653, n_13463);
  not g28746 (n_13464, n15665);
  not g28747 (n_13465, n15666);
  and g28748 (n15667, n_13464, n_13465);
  and g28749 (n15668, n_13066, n_13078);
  not g28750 (n_13466, n15668);
  and g28751 (n15669, n15667, n_13466);
  not g28752 (n_13467, n15667);
  and g28753 (n15670, n_13467, n15668);
  not g28754 (n_13468, n15669);
  not g28755 (n_13469, n15670);
  and g28756 (n15671, n_13468, n_13469);
  not g28757 (n_13470, n15495);
  and g28758 (n15672, n_13470, n15671);
  not g28759 (n_13471, n15672);
  and g28760 (n15673, n15671, n_13471);
  and g28761 (n15674, n_13470, n_13471);
  not g28762 (n_13472, n15673);
  not g28763 (n_13473, n15674);
  and g28764 (n15675, n_13472, n_13473);
  and g28765 (n15676, n_13080, n_13085);
  and g28766 (n15677, \b[38] , n3638);
  and g28767 (n15678, \b[36] , n3843);
  and g28768 (n15679, \b[37] , n3633);
  not g28769 (n_13474, n15678);
  not g28770 (n_13475, n15679);
  and g28771 (n15680, n_13474, n_13475);
  not g28772 (n_13476, n15677);
  and g28773 (n15681, n_13476, n15680);
  and g28774 (n15682, n_12780, n15681);
  not g28775 (n_13477, n5205);
  and g28776 (n15683, n_13477, n15681);
  not g28777 (n_13478, n15682);
  not g28778 (n_13479, n15683);
  and g28779 (n15684, n_13478, n_13479);
  not g28780 (n_13480, n15684);
  and g28781 (n15685, \a[32] , n_13480);
  and g28782 (n15686, n_2992, n15684);
  not g28783 (n_13481, n15685);
  not g28784 (n_13482, n15686);
  and g28785 (n15687, n_13481, n_13482);
  not g28786 (n_13483, n15676);
  not g28787 (n_13484, n15687);
  and g28788 (n15688, n_13483, n_13484);
  and g28789 (n15689, n15676, n15687);
  not g28790 (n_13485, n15688);
  not g28791 (n_13486, n15689);
  and g28792 (n15690, n_13485, n_13486);
  not g28793 (n_13487, n15675);
  and g28794 (n15691, n_13487, n15690);
  not g28795 (n_13488, n15691);
  and g28796 (n15692, n_13487, n_13488);
  and g28797 (n15693, n15690, n_13488);
  not g28798 (n_13489, n15692);
  not g28799 (n_13490, n15693);
  and g28800 (n15694, n_13489, n_13490);
  not g28801 (n_13491, n15694);
  and g28802 (n15695, n15484, n_13491);
  not g28803 (n_13492, n15695);
  and g28804 (n15696, n15484, n_13492);
  and g28805 (n15697, n_13491, n_13492);
  not g28806 (n_13493, n15696);
  not g28807 (n_13494, n15697);
  and g28808 (n15698, n_13493, n_13494);
  and g28809 (n15699, n_13103, n_13107);
  and g28810 (n15700, \b[44] , n2539);
  and g28811 (n15701, \b[42] , n2685);
  and g28812 (n15702, \b[43] , n2534);
  not g28813 (n_13495, n15701);
  not g28814 (n_13496, n15702);
  and g28815 (n15703, n_13495, n_13496);
  not g28816 (n_13497, n15700);
  and g28817 (n15704, n_13497, n15703);
  not g28818 (n_13498, n2542);
  and g28819 (n15705, n_13498, n15704);
  not g28820 (n_13499, n7072);
  and g28821 (n15706, n_13499, n15704);
  not g28822 (n_13500, n15705);
  not g28823 (n_13501, n15706);
  and g28824 (n15707, n_13500, n_13501);
  not g28825 (n_13502, n15707);
  and g28826 (n15708, \a[26] , n_13502);
  and g28827 (n15709, n_2025, n15707);
  not g28828 (n_13503, n15708);
  not g28829 (n_13504, n15709);
  and g28830 (n15710, n_13503, n_13504);
  not g28831 (n_13505, n15699);
  not g28832 (n_13506, n15710);
  and g28833 (n15711, n_13505, n_13506);
  not g28834 (n_13507, n15711);
  and g28835 (n15712, n_13505, n_13507);
  and g28836 (n15713, n_13506, n_13507);
  not g28837 (n_13508, n15712);
  not g28838 (n_13509, n15713);
  and g28839 (n15714, n_13508, n_13509);
  not g28840 (n_13510, n15698);
  not g28841 (n_13511, n15714);
  and g28842 (n15715, n_13510, n_13511);
  not g28843 (n_13512, n15715);
  and g28844 (n15716, n_13510, n_13512);
  and g28845 (n15717, n_13511, n_13512);
  not g28846 (n_13513, n15716);
  not g28847 (n_13514, n15717);
  and g28848 (n15718, n_13513, n_13514);
  not g28849 (n_13515, n15718);
  and g28850 (n15719, n15469, n_13515);
  not g28851 (n_13516, n15719);
  and g28852 (n15720, n15469, n_13516);
  and g28853 (n15721, n_13515, n_13516);
  not g28854 (n_13517, n15720);
  not g28855 (n_13518, n15721);
  and g28856 (n15722, n_13517, n_13518);
  not g28857 (n_13519, n15454);
  and g28858 (n15723, n_13519, n15722);
  not g28859 (n_13520, n15722);
  and g28860 (n15724, n15454, n_13520);
  not g28861 (n_13521, n15723);
  not g28862 (n_13522, n15724);
  and g28863 (n15725, n_13521, n_13522);
  not g28864 (n_13523, n15725);
  and g28865 (n15726, n15437, n_13523);
  not g28866 (n_13524, n15726);
  and g28867 (n15727, n15437, n_13524);
  and g28868 (n15728, n_13523, n_13524);
  not g28869 (n_13525, n15727);
  not g28870 (n_13526, n15728);
  and g28871 (n15729, n_13525, n_13526);
  not g28872 (n_13527, n15422);
  and g28873 (n15730, n_13527, n15729);
  not g28874 (n_13528, n15729);
  and g28875 (n15731, n15422, n_13528);
  not g28876 (n_13529, n15730);
  not g28877 (n_13530, n15731);
  and g28878 (n15732, n_13529, n_13530);
  not g28879 (n_13531, n15732);
  and g28880 (n15733, n15405, n_13531);
  not g28881 (n_13532, n15733);
  and g28882 (n15734, n15405, n_13532);
  and g28883 (n15735, n_13531, n_13532);
  not g28884 (n_13533, n15734);
  not g28885 (n_13534, n15735);
  and g28886 (n15736, n_13533, n_13534);
  and g28887 (n15737, n_13168, n_13173);
  and g28888 (n15738, \b[62] , n511);
  and g28889 (n15739, \b[60] , n541);
  and g28890 (n15740, \b[61] , n506);
  not g28891 (n_13535, n15739);
  not g28892 (n_13536, n15740);
  and g28893 (n15741, n_13535, n_13536);
  not g28894 (n_13537, n15738);
  and g28895 (n15742, n_13537, n15741);
  and g28896 (n15743, n_13179, n15742);
  not g28897 (n_13538, n13370);
  and g28898 (n15744, n_13538, n15742);
  not g28899 (n_13539, n15743);
  not g28900 (n_13540, n15744);
  and g28901 (n15745, n_13539, n_13540);
  not g28902 (n_13541, n15745);
  and g28903 (n15746, \a[8] , n_13541);
  and g28904 (n15747, n_234, n15745);
  not g28905 (n_13542, n15746);
  not g28906 (n_13543, n15747);
  and g28907 (n15748, n_13542, n_13543);
  not g28908 (n_13544, n15737);
  not g28909 (n_13545, n15748);
  and g28910 (n15749, n_13544, n_13545);
  not g28911 (n_13546, n15749);
  and g28912 (n15750, n_13544, n_13546);
  and g28913 (n15751, n_13545, n_13546);
  not g28914 (n_13547, n15750);
  not g28915 (n_13548, n15751);
  and g28916 (n15752, n_13547, n_13548);
  not g28917 (n_13549, n15736);
  not g28918 (n_13550, n15752);
  and g28919 (n15753, n_13549, n_13550);
  and g28920 (n15754, n15736, n_13548);
  and g28921 (n15755, n_13547, n15754);
  not g28922 (n_13551, n15753);
  not g28923 (n_13552, n15755);
  and g28924 (n15756, n_13551, n_13552);
  not g28925 (n_13553, n15390);
  and g28926 (n15757, n_13553, n15756);
  not g28927 (n_13554, n15756);
  and g28928 (n15758, n15390, n_13554);
  not g28929 (n_13555, n15757);
  not g28930 (n_13556, n15758);
  and g28931 (n15759, n_13555, n_13556);
  not g28932 (n_13557, n15378);
  and g28933 (n15760, n_13557, n15759);
  not g28934 (n_13558, n15760);
  and g28935 (n15761, n_13557, n_13558);
  and g28936 (n15762, n15759, n_13558);
  not g28937 (n_13559, n15761);
  not g28938 (n_13560, n15762);
  and g28939 (n15763, n_13559, n_13560);
  not g28940 (n_13561, n15377);
  not g28941 (n_13562, n15763);
  and g28942 (n15764, n_13561, n_13562);
  and g28943 (n15765, n15377, n_13560);
  and g28944 (n15766, n_13559, n15765);
  not g28945 (n_13563, n15764);
  not g28946 (n_13564, n15766);
  and g28947 (\f[68] , n_13563, n_13564);
  and g28948 (n15768, n_13558, n_13563);
  and g28949 (n15769, n_13228, n_13555);
  and g28950 (n15770, n_13546, n_13551);
  and g28951 (n15771, \b[63] , n511);
  and g28952 (n15772, \b[61] , n541);
  and g28953 (n15773, \b[62] , n506);
  and g28959 (n15776, n514, n13771);
  not g28962 (n_13569, n15777);
  and g28963 (n15778, \a[8] , n_13569);
  not g28964 (n_13570, n15778);
  and g28965 (n15779, \a[8] , n_13570);
  and g28966 (n15780, n_13569, n_13570);
  not g28967 (n_13571, n15779);
  not g28968 (n_13572, n15780);
  and g28969 (n15781, n_13571, n_13572);
  not g28970 (n_13573, n15770);
  not g28971 (n_13574, n15781);
  and g28972 (n15782, n_13573, n_13574);
  not g28973 (n_13575, n15782);
  and g28974 (n15783, n_13573, n_13575);
  and g28975 (n15784, n_13574, n_13575);
  not g28976 (n_13576, n15783);
  not g28977 (n_13577, n15784);
  and g28978 (n15785, n_13576, n_13577);
  and g28979 (n15786, \b[60] , n700);
  and g28980 (n15787, \b[58] , n767);
  and g28981 (n15788, \b[59] , n695);
  and g28987 (n15791, n703, n12211);
  not g28990 (n_13582, n15792);
  and g28991 (n15793, \a[11] , n_13582);
  not g28992 (n_13583, n15793);
  and g28993 (n15794, \a[11] , n_13583);
  and g28994 (n15795, n_13582, n_13583);
  not g28995 (n_13584, n15794);
  not g28996 (n_13585, n15795);
  and g28997 (n15796, n_13584, n_13585);
  and g28998 (n15797, n_13242, n_13532);
  and g28999 (n15798, n15796, n15797);
  not g29000 (n_13586, n15796);
  not g29001 (n_13587, n15797);
  and g29002 (n15799, n_13586, n_13587);
  not g29003 (n_13588, n15798);
  not g29004 (n_13589, n15799);
  and g29005 (n15800, n_13588, n_13589);
  and g29006 (n15801, n_13269, n_13524);
  and g29007 (n15802, \b[54] , n1302);
  and g29008 (n15803, \b[52] , n1391);
  and g29009 (n15804, \b[53] , n1297);
  and g29015 (n15807, n1305, n9998);
  not g29018 (n_13594, n15808);
  and g29019 (n15809, \a[17] , n_13594);
  not g29020 (n_13595, n15809);
  and g29021 (n15810, \a[17] , n_13595);
  and g29022 (n15811, n_13594, n_13595);
  not g29023 (n_13596, n15810);
  not g29024 (n_13597, n15811);
  and g29025 (n15812, n_13596, n_13597);
  not g29026 (n_13598, n15801);
  not g29027 (n_13599, n15812);
  and g29028 (n15813, n_13598, n_13599);
  not g29029 (n_13600, n15813);
  and g29030 (n15814, n_13598, n_13600);
  and g29031 (n15815, n_13599, n_13600);
  not g29032 (n_13601, n15814);
  not g29033 (n_13602, n15815);
  and g29034 (n15816, n_13601, n_13602);
  and g29035 (n15817, \b[48] , n2048);
  and g29036 (n15818, \b[46] , n2198);
  and g29037 (n15819, \b[47] , n2043);
  and g29043 (n15822, n2051, n8009);
  not g29046 (n_13607, n15823);
  and g29047 (n15824, \a[23] , n_13607);
  not g29048 (n_13608, n15824);
  and g29049 (n15825, \a[23] , n_13608);
  and g29050 (n15826, n_13607, n_13608);
  not g29051 (n_13609, n15825);
  not g29052 (n_13610, n15826);
  and g29053 (n15827, n_13609, n_13610);
  and g29054 (n15828, n_13296, n_13516);
  and g29055 (n15829, n15827, n15828);
  not g29056 (n_13611, n15827);
  not g29057 (n_13612, n15828);
  and g29058 (n15830, n_13611, n_13612);
  not g29059 (n_13613, n15829);
  not g29060 (n_13614, n15830);
  and g29061 (n15831, n_13613, n_13614);
  and g29062 (n15832, n_13507, n_13512);
  and g29063 (n15833, \b[45] , n2539);
  and g29064 (n15834, \b[43] , n2685);
  and g29065 (n15835, \b[44] , n2534);
  and g29071 (n15838, n2542, n7361);
  not g29074 (n_13619, n15839);
  and g29075 (n15840, \a[26] , n_13619);
  not g29076 (n_13620, n15840);
  and g29077 (n15841, \a[26] , n_13620);
  and g29078 (n15842, n_13619, n_13620);
  not g29079 (n_13621, n15841);
  not g29080 (n_13622, n15842);
  and g29081 (n15843, n_13621, n_13622);
  not g29082 (n_13623, n15832);
  not g29083 (n_13624, n15843);
  and g29084 (n15844, n_13623, n_13624);
  not g29085 (n_13625, n15844);
  and g29086 (n15845, n_13623, n_13625);
  and g29087 (n15846, n_13624, n_13625);
  not g29088 (n_13626, n15845);
  not g29089 (n_13627, n15846);
  and g29090 (n15847, n_13626, n_13627);
  and g29091 (n15848, \b[42] , n3050);
  and g29092 (n15849, \b[40] , n3243);
  and g29093 (n15850, \b[41] , n3045);
  and g29099 (n15853, n3053, n6489);
  not g29102 (n_13632, n15854);
  and g29103 (n15855, \a[29] , n_13632);
  not g29104 (n_13633, n15855);
  and g29105 (n15856, \a[29] , n_13633);
  and g29106 (n15857, n_13632, n_13633);
  not g29107 (n_13634, n15856);
  not g29108 (n_13635, n15857);
  and g29109 (n15858, n_13634, n_13635);
  and g29110 (n15859, n_13308, n_13492);
  and g29111 (n15860, n15858, n15859);
  not g29112 (n_13636, n15858);
  not g29113 (n_13637, n15859);
  and g29114 (n15861, n_13636, n_13637);
  not g29115 (n_13638, n15860);
  not g29116 (n_13639, n15861);
  and g29117 (n15862, n_13638, n_13639);
  and g29118 (n15863, n_13468, n_13471);
  and g29119 (n15864, n_13453, n_13465);
  and g29120 (n15865, n_13437, n_13447);
  and g29121 (n15866, n_13412, n_13415);
  and g29122 (n15867, n_13397, n_13409);
  and g29123 (n15868, n_13355, n_13367);
  and g29124 (n15869, \b[12] , n11531);
  and g29125 (n15870, \b[10] , n11896);
  and g29126 (n15871, \b[11] , n11526);
  and g29132 (n15874, n842, n11534);
  not g29135 (n_13644, n15875);
  and g29136 (n15876, \a[59] , n_13644);
  not g29137 (n_13645, n15876);
  and g29138 (n15877, \a[59] , n_13645);
  and g29139 (n15878, n_13644, n_13645);
  not g29140 (n_13646, n15877);
  not g29141 (n_13647, n15878);
  and g29142 (n15879, n_13646, n_13647);
  and g29143 (n15880, n_13344, n_13349);
  and g29144 (n15881, \b[5] , n13903);
  and g29145 (n15882, \b[6] , n_11555);
  not g29146 (n_13648, n15881);
  not g29147 (n_13649, n15882);
  and g29148 (n15883, n_13648, n_13649);
  and g29149 (n15884, \a[2] , n_99);
  and g29150 (n15885, n_5, \a[5] );
  not g29151 (n_13650, n15884);
  not g29152 (n_13651, n15885);
  and g29153 (n15886, n_13650, n_13651);
  not g29154 (n_13652, n15883);
  not g29155 (n_13653, n15886);
  and g29156 (n15887, n_13652, n_13653);
  and g29157 (n15888, n15883, n15886);
  not g29158 (n_13654, n15887);
  not g29159 (n_13655, n15888);
  and g29160 (n15889, n_13654, n_13655);
  not g29161 (n_13656, n15889);
  and g29162 (n15890, n15880, n_13656);
  not g29163 (n_13657, n15880);
  and g29164 (n15891, n_13657, n15889);
  not g29165 (n_13658, n15890);
  not g29166 (n_13659, n15891);
  and g29167 (n15892, n_13658, n_13659);
  and g29168 (n15893, \b[9] , n12668);
  and g29169 (n15894, \b[7] , n13047);
  and g29170 (n15895, \b[8] , n12663);
  and g29176 (n15898, n651, n12671);
  not g29179 (n_13664, n15899);
  and g29180 (n15900, \a[62] , n_13664);
  not g29181 (n_13665, n15900);
  and g29182 (n15901, \a[62] , n_13665);
  and g29183 (n15902, n_13664, n_13665);
  not g29184 (n_13666, n15901);
  not g29185 (n_13667, n15902);
  and g29186 (n15903, n_13666, n_13667);
  not g29187 (n_13668, n15892);
  and g29188 (n15904, n_13668, n15903);
  not g29189 (n_13669, n15903);
  and g29190 (n15905, n15892, n_13669);
  not g29191 (n_13670, n15904);
  not g29192 (n_13671, n15905);
  and g29193 (n15906, n_13670, n_13671);
  not g29194 (n_13672, n15879);
  and g29195 (n15907, n_13672, n15906);
  not g29196 (n_13673, n15907);
  and g29197 (n15908, n_13672, n_13673);
  and g29198 (n15909, n15906, n_13673);
  not g29199 (n_13674, n15908);
  not g29200 (n_13675, n15909);
  and g29201 (n15910, n_13674, n_13675);
  not g29202 (n_13676, n15868);
  not g29203 (n_13677, n15910);
  and g29204 (n15911, n_13676, n_13677);
  not g29205 (n_13678, n15911);
  and g29206 (n15912, n_13676, n_13678);
  and g29207 (n15913, n_13677, n_13678);
  not g29208 (n_13679, n15912);
  not g29209 (n_13680, n15913);
  and g29210 (n15914, n_13679, n_13680);
  and g29211 (n15915, \b[15] , n10426);
  and g29212 (n15916, \b[13] , n10796);
  and g29213 (n15917, \b[14] , n10421);
  and g29219 (n15920, n1131, n10429);
  not g29222 (n_13685, n15921);
  and g29223 (n15922, \a[56] , n_13685);
  not g29224 (n_13686, n15922);
  and g29225 (n15923, \a[56] , n_13686);
  and g29226 (n15924, n_13685, n_13686);
  not g29227 (n_13687, n15923);
  not g29228 (n_13688, n15924);
  and g29229 (n15925, n_13687, n_13688);
  not g29230 (n_13689, n15914);
  not g29231 (n_13690, n15925);
  and g29232 (n15926, n_13689, n_13690);
  not g29233 (n_13691, n15926);
  and g29234 (n15927, n_13689, n_13691);
  and g29235 (n15928, n_13690, n_13691);
  not g29236 (n_13692, n15927);
  not g29237 (n_13693, n15928);
  and g29238 (n15929, n_13692, n_13693);
  and g29239 (n15930, n_13370, n_13373);
  and g29240 (n15931, n15929, n15930);
  not g29241 (n_13694, n15929);
  not g29242 (n_13695, n15930);
  and g29243 (n15932, n_13694, n_13695);
  not g29244 (n_13696, n15931);
  not g29245 (n_13697, n15932);
  and g29246 (n15933, n_13696, n_13697);
  and g29247 (n15934, \b[18] , n9339);
  and g29248 (n15935, \b[16] , n9732);
  and g29249 (n15936, \b[17] , n9334);
  and g29255 (n15939, n1566, n9342);
  not g29258 (n_13702, n15940);
  and g29259 (n15941, \a[53] , n_13702);
  not g29260 (n_13703, n15941);
  and g29261 (n15942, \a[53] , n_13703);
  and g29262 (n15943, n_13702, n_13703);
  not g29263 (n_13704, n15942);
  not g29264 (n_13705, n15943);
  and g29265 (n15944, n_13704, n_13705);
  not g29266 (n_13706, n15944);
  and g29267 (n15945, n15933, n_13706);
  not g29268 (n_13707, n15945);
  and g29269 (n15946, n15933, n_13707);
  and g29270 (n15947, n_13706, n_13707);
  not g29271 (n_13708, n15946);
  not g29272 (n_13709, n15947);
  and g29273 (n15948, n_13708, n_13709);
  and g29274 (n15949, n_13378, n_13391);
  and g29275 (n15950, n15948, n15949);
  not g29276 (n_13710, n15948);
  not g29277 (n_13711, n15949);
  and g29278 (n15951, n_13710, n_13711);
  not g29279 (n_13712, n15950);
  not g29280 (n_13713, n15951);
  and g29281 (n15952, n_13712, n_13713);
  and g29282 (n15953, \b[21] , n8362);
  and g29283 (n15954, \b[19] , n8715);
  and g29284 (n15955, \b[20] , n8357);
  and g29290 (n15958, n1984, n8365);
  not g29293 (n_13718, n15959);
  and g29294 (n15960, \a[50] , n_13718);
  not g29295 (n_13719, n15960);
  and g29296 (n15961, \a[50] , n_13719);
  and g29297 (n15962, n_13718, n_13719);
  not g29298 (n_13720, n15961);
  not g29299 (n_13721, n15962);
  and g29300 (n15963, n_13720, n_13721);
  not g29301 (n_13722, n15963);
  and g29302 (n15964, n15952, n_13722);
  not g29303 (n_13723, n15964);
  and g29304 (n15965, n15952, n_13723);
  and g29305 (n15966, n_13722, n_13723);
  not g29306 (n_13724, n15965);
  not g29307 (n_13725, n15966);
  and g29308 (n15967, n_13724, n_13725);
  not g29309 (n_13726, n15867);
  and g29310 (n15968, n_13726, n15967);
  not g29311 (n_13727, n15967);
  and g29312 (n15969, n15867, n_13727);
  not g29313 (n_13728, n15968);
  not g29314 (n_13729, n15969);
  and g29315 (n15970, n_13728, n_13729);
  and g29316 (n15971, \b[24] , n7446);
  and g29317 (n15972, \b[22] , n7787);
  and g29318 (n15973, \b[23] , n7441);
  and g29324 (n15976, n2458, n7449);
  not g29327 (n_13734, n15977);
  and g29328 (n15978, \a[47] , n_13734);
  not g29329 (n_13735, n15978);
  and g29330 (n15979, \a[47] , n_13735);
  and g29331 (n15980, n_13734, n_13735);
  not g29332 (n_13736, n15979);
  not g29333 (n_13737, n15980);
  and g29334 (n15981, n_13736, n_13737);
  not g29335 (n_13738, n15970);
  not g29336 (n_13739, n15981);
  and g29337 (n15982, n_13738, n_13739);
  and g29338 (n15983, n15970, n15981);
  not g29339 (n_13740, n15982);
  not g29340 (n_13741, n15983);
  and g29341 (n15984, n_13740, n_13741);
  not g29342 (n_13742, n15984);
  and g29343 (n15985, n15866, n_13742);
  not g29344 (n_13743, n15866);
  and g29345 (n15986, n_13743, n15984);
  not g29346 (n_13744, n15985);
  not g29347 (n_13745, n15986);
  and g29348 (n15987, n_13744, n_13745);
  and g29349 (n15988, \b[27] , n6595);
  and g29350 (n15989, \b[25] , n6902);
  and g29351 (n15990, \b[26] , n6590);
  and g29357 (n15993, n2990, n6598);
  not g29360 (n_13750, n15994);
  and g29361 (n15995, \a[44] , n_13750);
  not g29362 (n_13751, n15995);
  and g29363 (n15996, \a[44] , n_13751);
  and g29364 (n15997, n_13750, n_13751);
  not g29365 (n_13752, n15996);
  not g29366 (n_13753, n15997);
  and g29367 (n15998, n_13752, n_13753);
  not g29368 (n_13754, n15998);
  and g29369 (n15999, n15987, n_13754);
  not g29370 (n_13755, n15999);
  and g29371 (n16000, n15987, n_13755);
  and g29372 (n16001, n_13754, n_13755);
  not g29373 (n_13756, n16000);
  not g29374 (n_13757, n16001);
  and g29375 (n16002, n_13756, n_13757);
  and g29376 (n16003, n_13421, n_13431);
  and g29377 (n16004, n16002, n16003);
  not g29378 (n_13758, n16002);
  not g29379 (n_13759, n16003);
  and g29380 (n16005, n_13758, n_13759);
  not g29381 (n_13760, n16004);
  not g29382 (n_13761, n16005);
  and g29383 (n16006, n_13760, n_13761);
  and g29384 (n16007, \b[30] , n5777);
  and g29385 (n16008, \b[28] , n6059);
  and g29386 (n16009, \b[29] , n5772);
  and g29392 (n16012, n3577, n5780);
  not g29395 (n_13766, n16013);
  and g29396 (n16014, \a[41] , n_13766);
  not g29397 (n_13767, n16014);
  and g29398 (n16015, \a[41] , n_13767);
  and g29399 (n16016, n_13766, n_13767);
  not g29400 (n_13768, n16015);
  not g29401 (n_13769, n16016);
  and g29402 (n16017, n_13768, n_13769);
  not g29403 (n_13770, n16017);
  and g29404 (n16018, n16006, n_13770);
  not g29405 (n_13771, n16006);
  and g29406 (n16019, n_13771, n16017);
  not g29407 (n_13772, n15865);
  not g29408 (n_13773, n16019);
  and g29409 (n16020, n_13772, n_13773);
  not g29410 (n_13774, n16018);
  and g29411 (n16021, n_13774, n16020);
  not g29412 (n_13775, n16021);
  and g29413 (n16022, n_13772, n_13775);
  and g29414 (n16023, n_13774, n_13775);
  and g29415 (n16024, n_13773, n16023);
  not g29416 (n_13776, n16022);
  not g29417 (n_13777, n16024);
  and g29418 (n16025, n_13776, n_13777);
  and g29419 (n16026, \b[33] , n5035);
  and g29420 (n16027, \b[31] , n5277);
  and g29421 (n16028, \b[32] , n5030);
  and g29427 (n16031, n4223, n5038);
  not g29430 (n_13782, n16032);
  and g29431 (n16033, \a[38] , n_13782);
  not g29432 (n_13783, n16033);
  and g29433 (n16034, \a[38] , n_13783);
  and g29434 (n16035, n_13782, n_13783);
  not g29435 (n_13784, n16034);
  not g29436 (n_13785, n16035);
  and g29437 (n16036, n_13784, n_13785);
  not g29438 (n_13786, n16025);
  not g29439 (n_13787, n16036);
  and g29440 (n16037, n_13786, n_13787);
  not g29441 (n_13788, n16037);
  and g29442 (n16038, n_13786, n_13788);
  and g29443 (n16039, n_13787, n_13788);
  not g29444 (n_13789, n16038);
  not g29445 (n_13790, n16039);
  and g29446 (n16040, n_13789, n_13790);
  not g29447 (n_13791, n15864);
  and g29448 (n16041, n_13791, n16040);
  not g29449 (n_13792, n16040);
  and g29450 (n16042, n15864, n_13792);
  not g29451 (n_13793, n16041);
  not g29452 (n_13794, n16042);
  and g29453 (n16043, n_13793, n_13794);
  and g29454 (n16044, \b[36] , n4287);
  and g29455 (n16045, \b[34] , n4532);
  and g29456 (n16046, \b[35] , n4282);
  and g29462 (n16049, n4290, n4922);
  not g29465 (n_13799, n16050);
  and g29466 (n16051, \a[35] , n_13799);
  not g29467 (n_13800, n16051);
  and g29468 (n16052, \a[35] , n_13800);
  and g29469 (n16053, n_13799, n_13800);
  not g29470 (n_13801, n16052);
  not g29471 (n_13802, n16053);
  and g29472 (n16054, n_13801, n_13802);
  not g29473 (n_13803, n16043);
  not g29474 (n_13804, n16054);
  and g29475 (n16055, n_13803, n_13804);
  and g29476 (n16056, n16043, n16054);
  not g29477 (n_13805, n16055);
  not g29478 (n_13806, n16056);
  and g29479 (n16057, n_13805, n_13806);
  not g29480 (n_13807, n16057);
  and g29481 (n16058, n15863, n_13807);
  not g29482 (n_13808, n15863);
  and g29483 (n16059, n_13808, n16057);
  not g29484 (n_13809, n16058);
  not g29485 (n_13810, n16059);
  and g29486 (n16060, n_13809, n_13810);
  and g29487 (n16061, \b[39] , n3638);
  and g29488 (n16062, \b[37] , n3843);
  and g29489 (n16063, \b[38] , n3633);
  and g29495 (n16066, n3641, n5451);
  not g29498 (n_13815, n16067);
  and g29499 (n16068, \a[32] , n_13815);
  not g29500 (n_13816, n16068);
  and g29501 (n16069, \a[32] , n_13816);
  and g29502 (n16070, n_13815, n_13816);
  not g29503 (n_13817, n16069);
  not g29504 (n_13818, n16070);
  and g29505 (n16071, n_13817, n_13818);
  and g29506 (n16072, n_13485, n_13488);
  and g29507 (n16073, n16071, n16072);
  not g29508 (n_13819, n16071);
  not g29509 (n_13820, n16072);
  and g29510 (n16074, n_13819, n_13820);
  not g29511 (n_13821, n16073);
  not g29512 (n_13822, n16074);
  and g29513 (n16075, n_13821, n_13822);
  and g29514 (n16076, n16060, n16075);
  not g29515 (n_13823, n16060);
  not g29516 (n_13824, n16075);
  and g29517 (n16077, n_13823, n_13824);
  not g29518 (n_13825, n16076);
  not g29519 (n_13826, n16077);
  and g29520 (n16078, n_13825, n_13826);
  and g29521 (n16079, n15862, n16078);
  not g29522 (n_13827, n15862);
  not g29523 (n_13828, n16078);
  and g29524 (n16080, n_13827, n_13828);
  not g29525 (n_13829, n16079);
  not g29526 (n_13830, n16080);
  and g29527 (n16081, n_13829, n_13830);
  not g29528 (n_13831, n15847);
  not g29529 (n_13832, n16081);
  and g29530 (n16082, n_13831, n_13832);
  and g29531 (n16083, n15847, n16081);
  not g29532 (n_13833, n16082);
  not g29533 (n_13834, n16083);
  and g29534 (n16084, n_13833, n_13834);
  not g29535 (n_13835, n16084);
  and g29536 (n16085, n15831, n_13835);
  not g29537 (n_13836, n16085);
  and g29538 (n16086, n15831, n_13836);
  and g29539 (n16087, n_13835, n_13836);
  not g29540 (n_13837, n16086);
  not g29541 (n_13838, n16087);
  and g29542 (n16088, n_13837, n_13838);
  and g29543 (n16089, \b[51] , n1627);
  and g29544 (n16090, \b[49] , n1763);
  and g29545 (n16091, \b[50] , n1622);
  and g29551 (n16094, n1630, n8976);
  not g29554 (n_13843, n16095);
  and g29555 (n16096, \a[20] , n_13843);
  not g29556 (n_13844, n16096);
  and g29557 (n16097, \a[20] , n_13844);
  and g29558 (n16098, n_13843, n_13844);
  not g29559 (n_13845, n16097);
  not g29560 (n_13846, n16098);
  and g29561 (n16099, n_13845, n_13846);
  and g29562 (n16100, n_13519, n_13520);
  not g29563 (n_13847, n16100);
  and g29564 (n16101, n_13282, n_13847);
  not g29565 (n_13848, n16099);
  not g29566 (n_13849, n16101);
  and g29567 (n16102, n_13848, n_13849);
  and g29568 (n16103, n16099, n16101);
  not g29569 (n_13850, n16102);
  not g29570 (n_13851, n16103);
  and g29571 (n16104, n_13850, n_13851);
  not g29572 (n_13852, n16088);
  and g29573 (n16105, n_13852, n16104);
  not g29574 (n_13853, n16105);
  and g29575 (n16106, n_13852, n_13853);
  and g29576 (n16107, n16104, n_13853);
  not g29577 (n_13854, n16106);
  not g29578 (n_13855, n16107);
  and g29579 (n16108, n_13854, n_13855);
  not g29580 (n_13856, n15816);
  not g29581 (n_13857, n16108);
  and g29582 (n16109, n_13856, n_13857);
  not g29583 (n_13858, n16109);
  and g29584 (n16110, n_13856, n_13858);
  and g29585 (n16111, n_13857, n_13858);
  not g29586 (n_13859, n16110);
  not g29587 (n_13860, n16111);
  and g29588 (n16112, n_13859, n_13860);
  and g29589 (n16113, \b[57] , n951);
  and g29590 (n16114, \b[55] , n1056);
  and g29591 (n16115, \b[56] , n946);
  and g29597 (n16118, n954, n11410);
  not g29600 (n_13865, n16119);
  and g29601 (n16120, \a[14] , n_13865);
  not g29602 (n_13866, n16120);
  and g29603 (n16121, \a[14] , n_13866);
  and g29604 (n16122, n_13865, n_13866);
  not g29605 (n_13867, n16121);
  not g29606 (n_13868, n16122);
  and g29607 (n16123, n_13867, n_13868);
  and g29608 (n16124, n_13527, n_13528);
  not g29609 (n_13869, n16124);
  and g29610 (n16125, n_13254, n_13869);
  not g29611 (n_13870, n16123);
  not g29612 (n_13871, n16125);
  and g29613 (n16126, n_13870, n_13871);
  and g29614 (n16127, n16123, n16125);
  not g29615 (n_13872, n16126);
  not g29616 (n_13873, n16127);
  and g29617 (n16128, n_13872, n_13873);
  not g29618 (n_13874, n16112);
  and g29619 (n16129, n_13874, n16128);
  not g29620 (n_13875, n16129);
  and g29621 (n16130, n_13874, n_13875);
  and g29622 (n16131, n16128, n_13875);
  not g29623 (n_13876, n16130);
  not g29624 (n_13877, n16131);
  and g29625 (n16132, n_13876, n_13877);
  not g29626 (n_13878, n16132);
  and g29627 (n16133, n15800, n_13878);
  not g29628 (n_13879, n16133);
  and g29629 (n16134, n15800, n_13879);
  and g29630 (n16135, n_13878, n_13879);
  not g29631 (n_13880, n16134);
  not g29632 (n_13881, n16135);
  and g29633 (n16136, n_13880, n_13881);
  not g29634 (n_13882, n15785);
  and g29635 (n16137, n_13882, n16136);
  not g29636 (n_13883, n16136);
  and g29637 (n16138, n15785, n_13883);
  not g29638 (n_13884, n16137);
  not g29639 (n_13885, n16138);
  and g29640 (n16139, n_13884, n_13885);
  not g29641 (n_13886, n15769);
  not g29642 (n_13887, n16139);
  and g29643 (n16140, n_13886, n_13887);
  and g29644 (n16141, n15769, n16139);
  not g29645 (n_13888, n16140);
  not g29646 (n_13889, n16141);
  and g29647 (n16142, n_13888, n_13889);
  not g29648 (n_13890, n15768);
  and g29649 (n16143, n_13890, n16142);
  not g29650 (n_13891, n16142);
  and g29651 (n16144, n15768, n_13891);
  not g29652 (n_13892, n16143);
  not g29653 (n_13893, n16144);
  and g29654 (\f[69] , n_13892, n_13893);
  and g29655 (n16146, n_13589, n_13879);
  and g29656 (n16147, \b[62] , n541);
  and g29657 (n16148, \b[63] , n506);
  not g29658 (n_13894, n16147);
  not g29659 (n_13895, n16148);
  and g29660 (n16149, n_13894, n_13895);
  and g29661 (n16150, n_13179, n16149);
  and g29662 (n16151, n13800, n16149);
  not g29663 (n_13896, n16150);
  not g29664 (n_13897, n16151);
  and g29665 (n16152, n_13896, n_13897);
  not g29666 (n_13898, n16152);
  and g29667 (n16153, \a[8] , n_13898);
  and g29668 (n16154, n_234, n16152);
  not g29669 (n_13899, n16153);
  not g29670 (n_13900, n16154);
  and g29671 (n16155, n_13899, n_13900);
  not g29672 (n_13901, n16146);
  not g29673 (n_13902, n16155);
  and g29674 (n16156, n_13901, n_13902);
  and g29675 (n16157, n16146, n16155);
  not g29676 (n_13903, n16156);
  not g29677 (n_13904, n16157);
  and g29678 (n16158, n_13903, n_13904);
  and g29679 (n16159, \b[61] , n700);
  and g29680 (n16160, \b[59] , n767);
  and g29681 (n16161, \b[60] , n695);
  and g29687 (n16164, n703, n12969);
  not g29690 (n_13909, n16165);
  and g29691 (n16166, \a[11] , n_13909);
  not g29692 (n_13910, n16166);
  and g29693 (n16167, \a[11] , n_13910);
  and g29694 (n16168, n_13909, n_13910);
  not g29695 (n_13911, n16167);
  not g29696 (n_13912, n16168);
  and g29697 (n16169, n_13911, n_13912);
  and g29698 (n16170, n_13872, n_13875);
  and g29699 (n16171, n16169, n16170);
  not g29700 (n_13913, n16169);
  not g29701 (n_13914, n16170);
  and g29702 (n16172, n_13913, n_13914);
  not g29703 (n_13915, n16171);
  not g29704 (n_13916, n16172);
  and g29705 (n16173, n_13915, n_13916);
  and g29706 (n16174, n_13600, n_13858);
  and g29707 (n16175, \b[58] , n951);
  and g29708 (n16176, \b[56] , n1056);
  and g29709 (n16177, \b[57] , n946);
  not g29710 (n_13917, n16176);
  not g29711 (n_13918, n16177);
  and g29712 (n16178, n_13917, n_13918);
  not g29713 (n_13919, n16175);
  and g29714 (n16179, n_13919, n16178);
  and g29715 (n16180, n_12819, n16179);
  and g29716 (n16181, n_13160, n16179);
  not g29717 (n_13920, n16180);
  not g29718 (n_13921, n16181);
  and g29719 (n16182, n_13920, n_13921);
  not g29720 (n_13922, n16182);
  and g29721 (n16183, \a[14] , n_13922);
  and g29722 (n16184, n_623, n16182);
  not g29723 (n_13923, n16183);
  not g29724 (n_13924, n16184);
  and g29725 (n16185, n_13923, n_13924);
  not g29726 (n_13925, n16174);
  not g29727 (n_13926, n16185);
  and g29728 (n16186, n_13925, n_13926);
  and g29729 (n16187, n16174, n16185);
  not g29730 (n_13927, n16186);
  not g29731 (n_13928, n16187);
  and g29732 (n16188, n_13927, n_13928);
  and g29733 (n16189, \b[55] , n1302);
  and g29734 (n16190, \b[53] , n1391);
  and g29735 (n16191, \b[54] , n1297);
  and g29741 (n16194, n1305, n10684);
  not g29744 (n_13933, n16195);
  and g29745 (n16196, \a[17] , n_13933);
  not g29746 (n_13934, n16196);
  and g29747 (n16197, \a[17] , n_13934);
  and g29748 (n16198, n_13933, n_13934);
  not g29749 (n_13935, n16197);
  not g29750 (n_13936, n16198);
  and g29751 (n16199, n_13935, n_13936);
  and g29752 (n16200, n_13850, n_13853);
  and g29753 (n16201, n16199, n16200);
  not g29754 (n_13937, n16199);
  not g29755 (n_13938, n16200);
  and g29756 (n16202, n_13937, n_13938);
  not g29757 (n_13939, n16201);
  not g29758 (n_13940, n16202);
  and g29759 (n16203, n_13939, n_13940);
  and g29760 (n16204, \b[52] , n1627);
  and g29761 (n16205, \b[50] , n1763);
  and g29762 (n16206, \b[51] , n1622);
  and g29768 (n16209, n1630, n9628);
  not g29771 (n_13945, n16210);
  and g29772 (n16211, \a[20] , n_13945);
  not g29773 (n_13946, n16211);
  and g29774 (n16212, \a[20] , n_13946);
  and g29775 (n16213, n_13945, n_13946);
  not g29776 (n_13947, n16212);
  not g29777 (n_13948, n16213);
  and g29778 (n16214, n_13947, n_13948);
  and g29779 (n16215, n_13614, n_13836);
  and g29780 (n16216, n16214, n16215);
  not g29781 (n_13949, n16214);
  not g29782 (n_13950, n16215);
  and g29783 (n16217, n_13949, n_13950);
  not g29784 (n_13951, n16216);
  not g29785 (n_13952, n16217);
  and g29786 (n16218, n_13951, n_13952);
  and g29787 (n16219, \b[49] , n2048);
  and g29788 (n16220, \b[47] , n2198);
  and g29789 (n16221, \b[48] , n2043);
  and g29795 (n16224, n2051, n8625);
  not g29798 (n_13957, n16225);
  and g29799 (n16226, \a[23] , n_13957);
  not g29800 (n_13958, n16226);
  and g29801 (n16227, \a[23] , n_13958);
  and g29802 (n16228, n_13957, n_13958);
  not g29803 (n_13959, n16227);
  not g29804 (n_13960, n16228);
  and g29805 (n16229, n_13959, n_13960);
  and g29806 (n16230, n_13831, n16081);
  not g29807 (n_13961, n16230);
  and g29808 (n16231, n_13625, n_13961);
  not g29809 (n_13962, n16229);
  not g29810 (n_13963, n16231);
  and g29811 (n16232, n_13962, n_13963);
  not g29812 (n_13964, n16232);
  and g29813 (n16233, n_13962, n_13964);
  and g29814 (n16234, n_13963, n_13964);
  not g29815 (n_13965, n16233);
  not g29816 (n_13966, n16234);
  and g29817 (n16235, n_13965, n_13966);
  and g29818 (n16236, n_13639, n_13829);
  and g29819 (n16237, \b[46] , n2539);
  and g29820 (n16238, \b[44] , n2685);
  and g29821 (n16239, \b[45] , n2534);
  not g29822 (n_13967, n16238);
  not g29823 (n_13968, n16239);
  and g29824 (n16240, n_13967, n_13968);
  not g29825 (n_13969, n16237);
  and g29826 (n16241, n_13969, n16240);
  and g29827 (n16242, n_13498, n16241);
  not g29828 (n_13970, n7677);
  and g29829 (n16243, n_13970, n16241);
  not g29830 (n_13971, n16242);
  not g29831 (n_13972, n16243);
  and g29832 (n16244, n_13971, n_13972);
  not g29833 (n_13973, n16244);
  and g29834 (n16245, \a[26] , n_13973);
  and g29835 (n16246, n_2025, n16244);
  not g29836 (n_13974, n16245);
  not g29837 (n_13975, n16246);
  and g29838 (n16247, n_13974, n_13975);
  not g29839 (n_13976, n16236);
  not g29840 (n_13977, n16247);
  and g29841 (n16248, n_13976, n_13977);
  and g29842 (n16249, n16236, n16247);
  not g29843 (n_13978, n16248);
  not g29844 (n_13979, n16249);
  and g29845 (n16250, n_13978, n_13979);
  and g29846 (n16251, \b[43] , n3050);
  and g29847 (n16252, \b[41] , n3243);
  and g29848 (n16253, \b[42] , n3045);
  and g29854 (n16256, n3053, n6515);
  not g29857 (n_13984, n16257);
  and g29858 (n16258, \a[29] , n_13984);
  not g29859 (n_13985, n16258);
  and g29860 (n16259, \a[29] , n_13985);
  and g29861 (n16260, n_13984, n_13985);
  not g29862 (n_13986, n16259);
  not g29863 (n_13987, n16260);
  and g29864 (n16261, n_13986, n_13987);
  and g29865 (n16262, n_13822, n_13825);
  not g29866 (n_13988, n16261);
  not g29867 (n_13989, n16262);
  and g29868 (n16263, n_13988, n_13989);
  not g29869 (n_13990, n16263);
  and g29870 (n16264, n_13988, n_13990);
  and g29871 (n16265, n_13989, n_13990);
  not g29872 (n_13991, n16264);
  not g29873 (n_13992, n16265);
  and g29874 (n16266, n_13991, n_13992);
  and g29875 (n16267, \b[40] , n3638);
  and g29876 (n16268, \b[38] , n3843);
  and g29877 (n16269, \b[39] , n3633);
  and g29883 (n16272, n3641, n5955);
  not g29886 (n_13997, n16273);
  and g29887 (n16274, \a[32] , n_13997);
  not g29888 (n_13998, n16274);
  and g29889 (n16275, \a[32] , n_13998);
  and g29890 (n16276, n_13997, n_13998);
  not g29891 (n_13999, n16275);
  not g29892 (n_14000, n16276);
  and g29893 (n16277, n_13999, n_14000);
  and g29894 (n16278, n_13805, n_13810);
  and g29895 (n16279, n16277, n16278);
  not g29896 (n_14001, n16277);
  not g29897 (n_14002, n16278);
  and g29898 (n16280, n_14001, n_14002);
  not g29899 (n_14003, n16279);
  not g29900 (n_14004, n16280);
  and g29901 (n16281, n_14003, n_14004);
  and g29902 (n16282, \b[37] , n4287);
  and g29903 (n16283, \b[35] , n4532);
  and g29904 (n16284, \b[36] , n4282);
  and g29910 (n16287, n4290, n5181);
  not g29913 (n_14009, n16288);
  and g29914 (n16289, \a[35] , n_14009);
  not g29915 (n_14010, n16289);
  and g29916 (n16290, \a[35] , n_14010);
  and g29917 (n16291, n_14009, n_14010);
  not g29918 (n_14011, n16290);
  not g29919 (n_14012, n16291);
  and g29920 (n16292, n_14011, n_14012);
  and g29921 (n16293, n_13791, n_13792);
  not g29922 (n_14013, n16293);
  and g29923 (n16294, n_13788, n_14013);
  and g29924 (n16295, \b[34] , n5035);
  and g29925 (n16296, \b[32] , n5277);
  and g29926 (n16297, \b[33] , n5030);
  and g29932 (n16300, n4466, n5038);
  not g29935 (n_14018, n16301);
  and g29936 (n16302, \a[38] , n_14018);
  not g29937 (n_14019, n16302);
  and g29938 (n16303, \a[38] , n_14019);
  and g29939 (n16304, n_14018, n_14019);
  not g29940 (n_14020, n16303);
  not g29941 (n_14021, n16304);
  and g29942 (n16305, n_14020, n_14021);
  and g29943 (n16306, n_13659, n_13671);
  and g29944 (n16307, n_5, n_99);
  not g29945 (n_14022, n16307);
  and g29946 (n16308, n_13654, n_14022);
  and g29947 (n16309, \b[6] , n13903);
  and g29948 (n16310, \b[7] , n_11555);
  not g29949 (n_14023, n16309);
  not g29950 (n_14024, n16310);
  and g29951 (n16311, n_14023, n_14024);
  not g29952 (n_14025, n16308);
  and g29953 (n16312, n_14025, n16311);
  not g29954 (n_14026, n16311);
  and g29955 (n16313, n16308, n_14026);
  not g29956 (n_14027, n16312);
  not g29957 (n_14028, n16313);
  and g29958 (n16314, n_14027, n_14028);
  and g29959 (n16315, \b[10] , n12668);
  and g29960 (n16316, \b[8] , n13047);
  and g29961 (n16317, \b[9] , n12663);
  not g29962 (n_14029, n16316);
  not g29963 (n_14030, n16317);
  and g29964 (n16318, n_14029, n_14030);
  not g29965 (n_14031, n16315);
  and g29966 (n16319, n_14031, n16318);
  and g29967 (n16320, n_12644, n16319);
  not g29968 (n_14032, n738);
  and g29969 (n16321, n_14032, n16319);
  not g29970 (n_14033, n16320);
  not g29971 (n_14034, n16321);
  and g29972 (n16322, n_14033, n_14034);
  not g29973 (n_14035, n16322);
  and g29974 (n16323, \a[62] , n_14035);
  and g29975 (n16324, n_10843, n16322);
  not g29976 (n_14036, n16323);
  not g29977 (n_14037, n16324);
  and g29978 (n16325, n_14036, n_14037);
  not g29979 (n_14038, n16325);
  and g29980 (n16326, n16314, n_14038);
  not g29981 (n_14039, n16314);
  and g29982 (n16327, n_14039, n16325);
  not g29983 (n_14040, n16326);
  not g29984 (n_14041, n16327);
  and g29985 (n16328, n_14040, n_14041);
  not g29986 (n_14042, n16306);
  and g29987 (n16329, n_14042, n16328);
  not g29988 (n_14043, n16328);
  and g29989 (n16330, n16306, n_14043);
  not g29990 (n_14044, n16329);
  not g29991 (n_14045, n16330);
  and g29992 (n16331, n_14044, n_14045);
  and g29993 (n16332, \b[13] , n11531);
  and g29994 (n16333, \b[11] , n11896);
  and g29995 (n16334, \b[12] , n11526);
  and g30001 (n16337, n1008, n11534);
  not g30004 (n_14050, n16338);
  and g30005 (n16339, \a[59] , n_14050);
  not g30006 (n_14051, n16339);
  and g30007 (n16340, \a[59] , n_14051);
  and g30008 (n16341, n_14050, n_14051);
  not g30009 (n_14052, n16340);
  not g30010 (n_14053, n16341);
  and g30011 (n16342, n_14052, n_14053);
  not g30012 (n_14054, n16342);
  and g30013 (n16343, n16331, n_14054);
  not g30014 (n_14055, n16343);
  and g30015 (n16344, n16331, n_14055);
  and g30016 (n16345, n_14054, n_14055);
  not g30017 (n_14056, n16344);
  not g30018 (n_14057, n16345);
  and g30019 (n16346, n_14056, n_14057);
  and g30020 (n16347, n_13673, n_13678);
  and g30021 (n16348, n16346, n16347);
  not g30022 (n_14058, n16346);
  not g30023 (n_14059, n16347);
  and g30024 (n16349, n_14058, n_14059);
  not g30025 (n_14060, n16348);
  not g30026 (n_14061, n16349);
  and g30027 (n16350, n_14060, n_14061);
  and g30028 (n16351, \b[16] , n10426);
  and g30029 (n16352, \b[14] , n10796);
  and g30030 (n16353, \b[15] , n10421);
  and g30036 (n16356, n1237, n10429);
  not g30039 (n_14066, n16357);
  and g30040 (n16358, \a[56] , n_14066);
  not g30041 (n_14067, n16358);
  and g30042 (n16359, \a[56] , n_14067);
  and g30043 (n16360, n_14066, n_14067);
  not g30044 (n_14068, n16359);
  not g30045 (n_14069, n16360);
  and g30046 (n16361, n_14068, n_14069);
  not g30047 (n_14070, n16361);
  and g30048 (n16362, n16350, n_14070);
  not g30049 (n_14071, n16362);
  and g30050 (n16363, n16350, n_14071);
  and g30051 (n16364, n_14070, n_14071);
  not g30052 (n_14072, n16363);
  not g30053 (n_14073, n16364);
  and g30054 (n16365, n_14072, n_14073);
  and g30055 (n16366, n_13691, n_13697);
  and g30056 (n16367, n16365, n16366);
  not g30057 (n_14074, n16365);
  not g30058 (n_14075, n16366);
  and g30059 (n16368, n_14074, n_14075);
  not g30060 (n_14076, n16367);
  not g30061 (n_14077, n16368);
  and g30062 (n16369, n_14076, n_14077);
  and g30063 (n16370, \b[19] , n9339);
  and g30064 (n16371, \b[17] , n9732);
  and g30065 (n16372, \b[18] , n9334);
  and g30071 (n16375, n1708, n9342);
  not g30074 (n_14082, n16376);
  and g30075 (n16377, \a[53] , n_14082);
  not g30076 (n_14083, n16377);
  and g30077 (n16378, \a[53] , n_14083);
  and g30078 (n16379, n_14082, n_14083);
  not g30079 (n_14084, n16378);
  not g30080 (n_14085, n16379);
  and g30081 (n16380, n_14084, n_14085);
  not g30082 (n_14086, n16380);
  and g30083 (n16381, n16369, n_14086);
  not g30084 (n_14087, n16381);
  and g30085 (n16382, n16369, n_14087);
  and g30086 (n16383, n_14086, n_14087);
  not g30087 (n_14088, n16382);
  not g30088 (n_14089, n16383);
  and g30089 (n16384, n_14088, n_14089);
  and g30090 (n16385, n_13707, n_13713);
  and g30091 (n16386, n16384, n16385);
  not g30092 (n_14090, n16384);
  not g30093 (n_14091, n16385);
  and g30094 (n16387, n_14090, n_14091);
  not g30095 (n_14092, n16386);
  not g30096 (n_14093, n16387);
  and g30097 (n16388, n_14092, n_14093);
  and g30098 (n16389, \b[22] , n8362);
  and g30099 (n16390, \b[20] , n8715);
  and g30100 (n16391, \b[21] , n8357);
  and g30106 (n16394, n2145, n8365);
  not g30109 (n_14098, n16395);
  and g30110 (n16396, \a[50] , n_14098);
  not g30111 (n_14099, n16396);
  and g30112 (n16397, \a[50] , n_14099);
  and g30113 (n16398, n_14098, n_14099);
  not g30114 (n_14100, n16397);
  not g30115 (n_14101, n16398);
  and g30116 (n16399, n_14100, n_14101);
  not g30117 (n_14102, n16399);
  and g30118 (n16400, n16388, n_14102);
  not g30119 (n_14103, n16400);
  and g30120 (n16401, n16388, n_14103);
  and g30121 (n16402, n_14102, n_14103);
  not g30122 (n_14104, n16401);
  not g30123 (n_14105, n16402);
  and g30124 (n16403, n_14104, n_14105);
  and g30125 (n16404, n_13726, n_13727);
  not g30126 (n_14106, n16404);
  and g30127 (n16405, n_13723, n_14106);
  and g30128 (n16406, n16403, n16405);
  not g30129 (n_14107, n16403);
  not g30130 (n_14108, n16405);
  and g30131 (n16407, n_14107, n_14108);
  not g30132 (n_14109, n16406);
  not g30133 (n_14110, n16407);
  and g30134 (n16408, n_14109, n_14110);
  and g30135 (n16409, \b[25] , n7446);
  and g30136 (n16410, \b[23] , n7787);
  and g30137 (n16411, \b[24] , n7441);
  and g30143 (n16414, n2485, n7449);
  not g30146 (n_14115, n16415);
  and g30147 (n16416, \a[47] , n_14115);
  not g30148 (n_14116, n16416);
  and g30149 (n16417, \a[47] , n_14116);
  and g30150 (n16418, n_14115, n_14116);
  not g30151 (n_14117, n16417);
  not g30152 (n_14118, n16418);
  and g30153 (n16419, n_14117, n_14118);
  not g30154 (n_14119, n16419);
  and g30155 (n16420, n16408, n_14119);
  not g30156 (n_14120, n16420);
  and g30157 (n16421, n16408, n_14120);
  and g30158 (n16422, n_14119, n_14120);
  not g30159 (n_14121, n16421);
  not g30160 (n_14122, n16422);
  and g30161 (n16423, n_14121, n_14122);
  and g30162 (n16424, n_13740, n_13745);
  and g30163 (n16425, n16423, n16424);
  not g30164 (n_14123, n16423);
  not g30165 (n_14124, n16424);
  and g30166 (n16426, n_14123, n_14124);
  not g30167 (n_14125, n16425);
  not g30168 (n_14126, n16426);
  and g30169 (n16427, n_14125, n_14126);
  and g30170 (n16428, \b[28] , n6595);
  and g30171 (n16429, \b[26] , n6902);
  and g30172 (n16430, \b[27] , n6590);
  and g30178 (n16433, n3189, n6598);
  not g30181 (n_14131, n16434);
  and g30182 (n16435, \a[44] , n_14131);
  not g30183 (n_14132, n16435);
  and g30184 (n16436, \a[44] , n_14132);
  and g30185 (n16437, n_14131, n_14132);
  not g30186 (n_14133, n16436);
  not g30187 (n_14134, n16437);
  and g30188 (n16438, n_14133, n_14134);
  not g30189 (n_14135, n16438);
  and g30190 (n16439, n16427, n_14135);
  not g30191 (n_14136, n16439);
  and g30192 (n16440, n16427, n_14136);
  and g30193 (n16441, n_14135, n_14136);
  not g30194 (n_14137, n16440);
  not g30195 (n_14138, n16441);
  and g30196 (n16442, n_14137, n_14138);
  and g30197 (n16443, n_13755, n_13761);
  and g30198 (n16444, n16442, n16443);
  not g30199 (n_14139, n16442);
  not g30200 (n_14140, n16443);
  and g30201 (n16445, n_14139, n_14140);
  not g30202 (n_14141, n16444);
  not g30203 (n_14142, n16445);
  and g30204 (n16446, n_14141, n_14142);
  and g30205 (n16447, \b[31] , n5777);
  and g30206 (n16448, \b[29] , n6059);
  and g30207 (n16449, \b[30] , n5772);
  and g30213 (n16452, n3796, n5780);
  not g30216 (n_14147, n16453);
  and g30217 (n16454, \a[41] , n_14147);
  not g30218 (n_14148, n16454);
  and g30219 (n16455, \a[41] , n_14148);
  and g30220 (n16456, n_14147, n_14148);
  not g30221 (n_14149, n16455);
  not g30222 (n_14150, n16456);
  and g30223 (n16457, n_14149, n_14150);
  not g30224 (n_14151, n16446);
  and g30225 (n16458, n_14151, n16457);
  not g30226 (n_14152, n16457);
  and g30227 (n16459, n16446, n_14152);
  not g30228 (n_14153, n16458);
  not g30229 (n_14154, n16459);
  and g30230 (n16460, n_14153, n_14154);
  not g30231 (n_14155, n16023);
  and g30232 (n16461, n_14155, n16460);
  not g30233 (n_14156, n16460);
  and g30234 (n16462, n16023, n_14156);
  not g30235 (n_14157, n16461);
  not g30236 (n_14158, n16462);
  and g30237 (n16463, n_14157, n_14158);
  not g30238 (n_14159, n16305);
  and g30239 (n16464, n_14159, n16463);
  not g30240 (n_14160, n16463);
  and g30241 (n16465, n16305, n_14160);
  not g30242 (n_14161, n16464);
  not g30243 (n_14162, n16465);
  and g30244 (n16466, n_14161, n_14162);
  not g30245 (n_14163, n16294);
  and g30246 (n16467, n_14163, n16466);
  not g30247 (n_14164, n16466);
  and g30248 (n16468, n16294, n_14164);
  not g30249 (n_14165, n16467);
  not g30250 (n_14166, n16468);
  and g30251 (n16469, n_14165, n_14166);
  not g30252 (n_14167, n16292);
  and g30253 (n16470, n_14167, n16469);
  not g30254 (n_14168, n16470);
  and g30255 (n16471, n_14167, n_14168);
  and g30256 (n16472, n16469, n_14168);
  not g30257 (n_14169, n16471);
  not g30258 (n_14170, n16472);
  and g30259 (n16473, n_14169, n_14170);
  not g30260 (n_14171, n16473);
  and g30261 (n16474, n16281, n_14171);
  not g30262 (n_14172, n16474);
  and g30263 (n16475, n16281, n_14172);
  and g30264 (n16476, n_14171, n_14172);
  not g30265 (n_14173, n16475);
  not g30266 (n_14174, n16476);
  and g30267 (n16477, n_14173, n_14174);
  not g30268 (n_14175, n16266);
  and g30269 (n16478, n_14175, n16477);
  not g30270 (n_14176, n16477);
  and g30271 (n16479, n16266, n_14176);
  not g30272 (n_14177, n16478);
  not g30273 (n_14178, n16479);
  and g30274 (n16480, n_14177, n_14178);
  not g30275 (n_14179, n16480);
  and g30276 (n16481, n16250, n_14179);
  not g30277 (n_14180, n16481);
  and g30278 (n16482, n16250, n_14180);
  and g30279 (n16483, n_14179, n_14180);
  not g30280 (n_14181, n16482);
  not g30281 (n_14182, n16483);
  and g30282 (n16484, n_14181, n_14182);
  not g30283 (n_14183, n16235);
  and g30284 (n16485, n_14183, n16484);
  not g30285 (n_14184, n16484);
  and g30286 (n16486, n16235, n_14184);
  not g30287 (n_14185, n16485);
  not g30288 (n_14186, n16486);
  and g30289 (n16487, n_14185, n_14186);
  not g30290 (n_14187, n16487);
  and g30291 (n16488, n16218, n_14187);
  not g30292 (n_14188, n16488);
  and g30293 (n16489, n16218, n_14188);
  and g30294 (n16490, n_14187, n_14188);
  not g30295 (n_14189, n16489);
  not g30296 (n_14190, n16490);
  and g30297 (n16491, n_14189, n_14190);
  not g30298 (n_14191, n16491);
  and g30299 (n16492, n16203, n_14191);
  not g30300 (n_14192, n16203);
  and g30301 (n16493, n_14192, n16491);
  not g30302 (n_14193, n16493);
  and g30303 (n16494, n16188, n_14193);
  not g30304 (n_14194, n16492);
  and g30305 (n16495, n_14194, n16494);
  not g30306 (n_14195, n16495);
  and g30307 (n16496, n16188, n_14195);
  and g30308 (n16497, n_14193, n_14195);
  and g30309 (n16498, n_14194, n16497);
  not g30310 (n_14196, n16496);
  not g30311 (n_14197, n16498);
  and g30312 (n16499, n_14196, n_14197);
  not g30313 (n_14198, n16499);
  and g30314 (n16500, n16173, n_14198);
  not g30315 (n_14199, n16173);
  and g30316 (n16501, n_14199, n16499);
  not g30317 (n_14200, n16501);
  and g30318 (n16502, n16158, n_14200);
  not g30319 (n_14201, n16500);
  and g30320 (n16503, n_14201, n16502);
  not g30321 (n_14202, n16503);
  and g30322 (n16504, n16158, n_14202);
  and g30323 (n16505, n_14200, n_14202);
  and g30324 (n16506, n_14201, n16505);
  not g30325 (n_14203, n16504);
  not g30326 (n_14204, n16506);
  and g30327 (n16507, n_14203, n_14204);
  and g30328 (n16508, n_13882, n_13883);
  not g30329 (n_14205, n16508);
  and g30330 (n16509, n_13575, n_14205);
  not g30331 (n_14206, n16507);
  not g30332 (n_14207, n16509);
  and g30333 (n16510, n_14206, n_14207);
  not g30334 (n_14208, n16510);
  and g30335 (n16511, n_14206, n_14208);
  and g30336 (n16512, n_14207, n_14208);
  not g30337 (n_14209, n16511);
  not g30338 (n_14210, n16512);
  and g30339 (n16513, n_14209, n_14210);
  and g30340 (n16514, n_13888, n_13892);
  not g30341 (n_14211, n16513);
  not g30342 (n_14212, n16514);
  and g30343 (n16515, n_14211, n_14212);
  and g30344 (n16516, n16513, n16514);
  not g30345 (n_14213, n16515);
  not g30346 (n_14214, n16516);
  and g30347 (\f[70] , n_14213, n_14214);
  and g30348 (n16518, n_14208, n_14213);
  and g30349 (n16519, n_13903, n_14202);
  and g30350 (n16520, n_13916, n_14201);
  and g30351 (n16521, \b[63] , n541);
  and g30352 (n16522, n514, n13797);
  not g30353 (n_14215, n16521);
  not g30354 (n_14216, n16522);
  and g30355 (n16523, n_14215, n_14216);
  not g30356 (n_14217, n16523);
  and g30357 (n16524, \a[8] , n_14217);
  not g30358 (n_14218, n16524);
  and g30359 (n16525, \a[8] , n_14218);
  and g30360 (n16526, n_14217, n_14218);
  not g30361 (n_14219, n16525);
  not g30362 (n_14220, n16526);
  and g30363 (n16527, n_14219, n_14220);
  not g30364 (n_14221, n16520);
  not g30365 (n_14222, n16527);
  and g30366 (n16528, n_14221, n_14222);
  not g30367 (n_14223, n16528);
  and g30368 (n16529, n_14221, n_14223);
  and g30369 (n16530, n_14222, n_14223);
  not g30370 (n_14224, n16529);
  not g30371 (n_14225, n16530);
  and g30372 (n16531, n_14224, n_14225);
  and g30373 (n16532, \b[56] , n1302);
  and g30374 (n16533, \b[54] , n1391);
  and g30375 (n16534, \b[55] , n1297);
  and g30381 (n16537, n1305, n10708);
  not g30384 (n_14230, n16538);
  and g30385 (n16539, \a[17] , n_14230);
  not g30386 (n_14231, n16539);
  and g30387 (n16540, \a[17] , n_14231);
  and g30388 (n16541, n_14230, n_14231);
  not g30389 (n_14232, n16540);
  not g30390 (n_14233, n16541);
  and g30391 (n16542, n_14232, n_14233);
  and g30392 (n16543, n_13952, n_14188);
  and g30393 (n16544, n16542, n16543);
  not g30394 (n_14234, n16542);
  not g30395 (n_14235, n16543);
  and g30396 (n16545, n_14234, n_14235);
  not g30397 (n_14236, n16544);
  not g30398 (n_14237, n16545);
  and g30399 (n16546, n_14236, n_14237);
  and g30400 (n16547, \b[50] , n2048);
  and g30401 (n16548, \b[48] , n2198);
  and g30402 (n16549, \b[49] , n2043);
  and g30408 (n16552, n2051, n8949);
  not g30411 (n_14242, n16553);
  and g30412 (n16554, \a[23] , n_14242);
  not g30413 (n_14243, n16554);
  and g30414 (n16555, \a[23] , n_14243);
  and g30415 (n16556, n_14242, n_14243);
  not g30416 (n_14244, n16555);
  not g30417 (n_14245, n16556);
  and g30418 (n16557, n_14244, n_14245);
  and g30419 (n16558, n_13978, n_14180);
  and g30420 (n16559, n16557, n16558);
  not g30421 (n_14246, n16557);
  not g30422 (n_14247, n16558);
  and g30423 (n16560, n_14246, n_14247);
  not g30424 (n_14248, n16559);
  not g30425 (n_14249, n16560);
  and g30426 (n16561, n_14248, n_14249);
  and g30427 (n16562, \b[47] , n2539);
  and g30428 (n16563, \b[45] , n2685);
  and g30429 (n16564, \b[46] , n2534);
  and g30435 (n16567, n2542, n7703);
  not g30438 (n_14254, n16568);
  and g30439 (n16569, \a[26] , n_14254);
  not g30440 (n_14255, n16569);
  and g30441 (n16570, \a[26] , n_14255);
  and g30442 (n16571, n_14254, n_14255);
  not g30443 (n_14256, n16570);
  not g30444 (n_14257, n16571);
  and g30445 (n16572, n_14256, n_14257);
  and g30446 (n16573, n_14175, n_14176);
  not g30447 (n_14258, n16573);
  and g30448 (n16574, n_13990, n_14258);
  not g30449 (n_14259, n16572);
  not g30450 (n_14260, n16574);
  and g30451 (n16575, n_14259, n_14260);
  not g30452 (n_14261, n16575);
  and g30453 (n16576, n_14259, n_14261);
  and g30454 (n16577, n_14260, n_14261);
  not g30455 (n_14262, n16576);
  not g30456 (n_14263, n16577);
  and g30457 (n16578, n_14262, n_14263);
  and g30458 (n16579, \b[41] , n3638);
  and g30459 (n16580, \b[39] , n3843);
  and g30460 (n16581, \b[40] , n3633);
  and g30466 (n16584, n3641, n6219);
  not g30469 (n_14268, n16585);
  and g30470 (n16586, \a[32] , n_14268);
  not g30471 (n_14269, n16586);
  and g30472 (n16587, \a[32] , n_14269);
  and g30473 (n16588, n_14268, n_14269);
  not g30474 (n_14270, n16587);
  not g30475 (n_14271, n16588);
  and g30476 (n16589, n_14270, n_14271);
  and g30477 (n16590, n_14165, n_14168);
  and g30478 (n16591, n16589, n16590);
  not g30479 (n_14272, n16589);
  not g30480 (n_14273, n16590);
  and g30481 (n16592, n_14272, n_14273);
  not g30482 (n_14274, n16591);
  not g30483 (n_14275, n16592);
  and g30484 (n16593, n_14274, n_14275);
  and g30485 (n16594, \b[35] , n5035);
  and g30486 (n16595, \b[33] , n5277);
  and g30487 (n16596, \b[34] , n5030);
  and g30493 (n16599, n4696, n5038);
  not g30496 (n_14280, n16600);
  and g30497 (n16601, \a[38] , n_14280);
  not g30498 (n_14281, n16601);
  and g30499 (n16602, \a[38] , n_14281);
  and g30500 (n16603, n_14280, n_14281);
  not g30501 (n_14282, n16602);
  not g30502 (n_14283, n16603);
  and g30503 (n16604, n_14282, n_14283);
  and g30504 (n16605, \b[26] , n7446);
  and g30505 (n16606, \b[24] , n7787);
  and g30506 (n16607, \b[25] , n7441);
  and g30512 (n16610, n2813, n7449);
  not g30515 (n_14288, n16611);
  and g30516 (n16612, \a[47] , n_14288);
  not g30517 (n_14289, n16612);
  and g30518 (n16613, \a[47] , n_14289);
  and g30519 (n16614, n_14288, n_14289);
  not g30520 (n_14290, n16613);
  not g30521 (n_14291, n16614);
  and g30522 (n16615, n_14290, n_14291);
  and g30523 (n16616, n_14093, n_14103);
  and g30524 (n16617, \b[23] , n8362);
  and g30525 (n16618, \b[21] , n8715);
  and g30526 (n16619, \b[22] , n8357);
  and g30532 (n16622, n2300, n8365);
  not g30535 (n_14296, n16623);
  and g30536 (n16624, \a[50] , n_14296);
  not g30537 (n_14297, n16624);
  and g30538 (n16625, \a[50] , n_14297);
  and g30539 (n16626, n_14296, n_14297);
  not g30540 (n_14298, n16625);
  not g30541 (n_14299, n16626);
  and g30542 (n16627, n_14298, n_14299);
  and g30543 (n16628, n_14077, n_14087);
  and g30544 (n16629, n_14044, n_14055);
  and g30545 (n16630, n_14027, n_14040);
  and g30546 (n16631, \b[7] , n13903);
  and g30547 (n16632, \b[8] , n_11555);
  not g30548 (n_14300, n16631);
  not g30549 (n_14301, n16632);
  and g30550 (n16633, n_14300, n_14301);
  not g30551 (n_14302, n16633);
  and g30552 (n16634, n16311, n_14302);
  and g30553 (n16635, n_14026, n16633);
  not g30554 (n_14303, n16630);
  not g30555 (n_14304, n16635);
  and g30556 (n16636, n_14303, n_14304);
  not g30557 (n_14305, n16634);
  and g30558 (n16637, n_14305, n16636);
  not g30559 (n_14306, n16637);
  and g30560 (n16638, n_14303, n_14306);
  and g30561 (n16639, n_14304, n_14306);
  and g30562 (n16640, n_14305, n16639);
  not g30563 (n_14307, n16638);
  not g30564 (n_14308, n16640);
  and g30565 (n16641, n_14307, n_14308);
  and g30566 (n16642, \b[11] , n12668);
  and g30567 (n16643, \b[9] , n13047);
  and g30568 (n16644, \b[10] , n12663);
  and g30574 (n16647, n818, n12671);
  not g30577 (n_14313, n16648);
  and g30578 (n16649, \a[62] , n_14313);
  not g30579 (n_14314, n16649);
  and g30580 (n16650, \a[62] , n_14314);
  and g30581 (n16651, n_14313, n_14314);
  not g30582 (n_14315, n16650);
  not g30583 (n_14316, n16651);
  and g30584 (n16652, n_14315, n_14316);
  not g30585 (n_14317, n16641);
  and g30586 (n16653, n_14317, n16652);
  not g30587 (n_14318, n16652);
  and g30588 (n16654, n16641, n_14318);
  not g30589 (n_14319, n16653);
  not g30590 (n_14320, n16654);
  and g30591 (n16655, n_14319, n_14320);
  and g30592 (n16656, \b[14] , n11531);
  and g30593 (n16657, \b[12] , n11896);
  and g30594 (n16658, \b[13] , n11526);
  and g30600 (n16661, n1034, n11534);
  not g30603 (n_14325, n16662);
  and g30604 (n16663, \a[59] , n_14325);
  not g30605 (n_14326, n16663);
  and g30606 (n16664, \a[59] , n_14326);
  and g30607 (n16665, n_14325, n_14326);
  not g30608 (n_14327, n16664);
  not g30609 (n_14328, n16665);
  and g30610 (n16666, n_14327, n_14328);
  not g30611 (n_14329, n16655);
  not g30612 (n_14330, n16666);
  and g30613 (n16667, n_14329, n_14330);
  and g30614 (n16668, n16655, n16666);
  not g30615 (n_14331, n16667);
  not g30616 (n_14332, n16668);
  and g30617 (n16669, n_14331, n_14332);
  not g30618 (n_14333, n16669);
  and g30619 (n16670, n16629, n_14333);
  not g30620 (n_14334, n16629);
  and g30621 (n16671, n_14334, n16669);
  not g30622 (n_14335, n16670);
  not g30623 (n_14336, n16671);
  and g30624 (n16672, n_14335, n_14336);
  and g30625 (n16673, \b[17] , n10426);
  and g30626 (n16674, \b[15] , n10796);
  and g30627 (n16675, \b[16] , n10421);
  and g30633 (n16678, n1356, n10429);
  not g30636 (n_14341, n16679);
  and g30637 (n16680, \a[56] , n_14341);
  not g30638 (n_14342, n16680);
  and g30639 (n16681, \a[56] , n_14342);
  and g30640 (n16682, n_14341, n_14342);
  not g30641 (n_14343, n16681);
  not g30642 (n_14344, n16682);
  and g30643 (n16683, n_14343, n_14344);
  not g30644 (n_14345, n16683);
  and g30645 (n16684, n16672, n_14345);
  not g30646 (n_14346, n16684);
  and g30647 (n16685, n16672, n_14346);
  and g30648 (n16686, n_14345, n_14346);
  not g30649 (n_14347, n16685);
  not g30650 (n_14348, n16686);
  and g30651 (n16687, n_14347, n_14348);
  and g30652 (n16688, n_14061, n_14071);
  and g30653 (n16689, n16687, n16688);
  not g30654 (n_14349, n16687);
  not g30655 (n_14350, n16688);
  and g30656 (n16690, n_14349, n_14350);
  not g30657 (n_14351, n16689);
  not g30658 (n_14352, n16690);
  and g30659 (n16691, n_14351, n_14352);
  and g30660 (n16692, \b[20] , n9339);
  and g30661 (n16693, \b[18] , n9732);
  and g30662 (n16694, \b[19] , n9334);
  and g30668 (n16697, n1846, n9342);
  not g30671 (n_14357, n16698);
  and g30672 (n16699, \a[53] , n_14357);
  not g30673 (n_14358, n16699);
  and g30674 (n16700, \a[53] , n_14358);
  and g30675 (n16701, n_14357, n_14358);
  not g30676 (n_14359, n16700);
  not g30677 (n_14360, n16701);
  and g30678 (n16702, n_14359, n_14360);
  not g30679 (n_14361, n16691);
  and g30680 (n16703, n_14361, n16702);
  not g30681 (n_14362, n16702);
  and g30682 (n16704, n16691, n_14362);
  not g30683 (n_14363, n16703);
  not g30684 (n_14364, n16704);
  and g30685 (n16705, n_14363, n_14364);
  not g30686 (n_14365, n16628);
  and g30687 (n16706, n_14365, n16705);
  not g30688 (n_14366, n16706);
  and g30689 (n16707, n_14365, n_14366);
  and g30690 (n16708, n16705, n_14366);
  not g30691 (n_14367, n16707);
  not g30692 (n_14368, n16708);
  and g30693 (n16709, n_14367, n_14368);
  not g30694 (n_14369, n16627);
  not g30695 (n_14370, n16709);
  and g30696 (n16710, n_14369, n_14370);
  and g30697 (n16711, n16627, n_14368);
  and g30698 (n16712, n_14367, n16711);
  not g30699 (n_14371, n16710);
  not g30700 (n_14372, n16712);
  and g30701 (n16713, n_14371, n_14372);
  not g30702 (n_14373, n16616);
  and g30703 (n16714, n_14373, n16713);
  not g30704 (n_14374, n16713);
  and g30705 (n16715, n16616, n_14374);
  not g30706 (n_14375, n16714);
  not g30707 (n_14376, n16715);
  and g30708 (n16716, n_14375, n_14376);
  not g30709 (n_14377, n16615);
  and g30710 (n16717, n_14377, n16716);
  not g30711 (n_14378, n16717);
  and g30712 (n16718, n16716, n_14378);
  and g30713 (n16719, n_14377, n_14378);
  not g30714 (n_14379, n16718);
  not g30715 (n_14380, n16719);
  and g30716 (n16720, n_14379, n_14380);
  and g30717 (n16721, n_14110, n_14120);
  and g30718 (n16722, n16720, n16721);
  not g30719 (n_14381, n16720);
  not g30720 (n_14382, n16721);
  and g30721 (n16723, n_14381, n_14382);
  not g30722 (n_14383, n16722);
  not g30723 (n_14384, n16723);
  and g30724 (n16724, n_14383, n_14384);
  and g30725 (n16725, \b[29] , n6595);
  and g30726 (n16726, \b[27] , n6902);
  and g30727 (n16727, \b[28] , n6590);
  and g30733 (n16730, n3383, n6598);
  not g30736 (n_14389, n16731);
  and g30737 (n16732, \a[44] , n_14389);
  not g30738 (n_14390, n16732);
  and g30739 (n16733, \a[44] , n_14390);
  and g30740 (n16734, n_14389, n_14390);
  not g30741 (n_14391, n16733);
  not g30742 (n_14392, n16734);
  and g30743 (n16735, n_14391, n_14392);
  not g30744 (n_14393, n16735);
  and g30745 (n16736, n16724, n_14393);
  not g30746 (n_14394, n16736);
  and g30747 (n16737, n16724, n_14394);
  and g30748 (n16738, n_14393, n_14394);
  not g30749 (n_14395, n16737);
  not g30750 (n_14396, n16738);
  and g30751 (n16739, n_14395, n_14396);
  and g30752 (n16740, n_14126, n_14136);
  and g30753 (n16741, n16739, n16740);
  not g30754 (n_14397, n16739);
  not g30755 (n_14398, n16740);
  and g30756 (n16742, n_14397, n_14398);
  not g30757 (n_14399, n16741);
  not g30758 (n_14400, n16742);
  and g30759 (n16743, n_14399, n_14400);
  and g30760 (n16744, \b[32] , n5777);
  and g30761 (n16745, \b[30] , n6059);
  and g30762 (n16746, \b[31] , n5772);
  and g30768 (n16749, n4013, n5780);
  not g30771 (n_14405, n16750);
  and g30772 (n16751, \a[41] , n_14405);
  not g30773 (n_14406, n16751);
  and g30774 (n16752, \a[41] , n_14406);
  and g30775 (n16753, n_14405, n_14406);
  not g30776 (n_14407, n16752);
  not g30777 (n_14408, n16753);
  and g30778 (n16754, n_14407, n_14408);
  not g30779 (n_14409, n16743);
  and g30780 (n16755, n_14409, n16754);
  not g30781 (n_14410, n16754);
  and g30782 (n16756, n16743, n_14410);
  not g30783 (n_14411, n16755);
  not g30784 (n_14412, n16756);
  and g30785 (n16757, n_14411, n_14412);
  and g30786 (n16758, n_14142, n_14154);
  not g30787 (n_14413, n16758);
  and g30788 (n16759, n16757, n_14413);
  not g30789 (n_14414, n16757);
  and g30790 (n16760, n_14414, n16758);
  not g30791 (n_14415, n16759);
  not g30792 (n_14416, n16760);
  and g30793 (n16761, n_14415, n_14416);
  not g30794 (n_14417, n16604);
  and g30795 (n16762, n_14417, n16761);
  not g30796 (n_14418, n16762);
  and g30797 (n16763, n16761, n_14418);
  and g30798 (n16764, n_14417, n_14418);
  not g30799 (n_14419, n16763);
  not g30800 (n_14420, n16764);
  and g30801 (n16765, n_14419, n_14420);
  and g30802 (n16766, n_14157, n_14161);
  and g30803 (n16767, n16765, n16766);
  not g30804 (n_14421, n16765);
  not g30805 (n_14422, n16766);
  and g30806 (n16768, n_14421, n_14422);
  not g30807 (n_14423, n16767);
  not g30808 (n_14424, n16768);
  and g30809 (n16769, n_14423, n_14424);
  and g30810 (n16770, \b[38] , n4287);
  and g30811 (n16771, \b[36] , n4532);
  and g30812 (n16772, \b[37] , n4282);
  and g30818 (n16775, n4290, n5205);
  not g30821 (n_14429, n16776);
  and g30822 (n16777, \a[35] , n_14429);
  not g30823 (n_14430, n16777);
  and g30824 (n16778, \a[35] , n_14430);
  and g30825 (n16779, n_14429, n_14430);
  not g30826 (n_14431, n16778);
  not g30827 (n_14432, n16779);
  and g30828 (n16780, n_14431, n_14432);
  not g30829 (n_14433, n16780);
  and g30830 (n16781, n16769, n_14433);
  not g30831 (n_14434, n16769);
  and g30832 (n16782, n_14434, n16780);
  not g30833 (n_14435, n16782);
  and g30834 (n16783, n16593, n_14435);
  not g30835 (n_14436, n16781);
  and g30836 (n16784, n_14436, n16783);
  not g30837 (n_14437, n16784);
  and g30838 (n16785, n16593, n_14437);
  and g30839 (n16786, n_14435, n_14437);
  and g30840 (n16787, n_14436, n16786);
  not g30841 (n_14438, n16785);
  not g30842 (n_14439, n16787);
  and g30843 (n16788, n_14438, n_14439);
  and g30844 (n16789, n_14004, n_14172);
  and g30845 (n16790, \b[44] , n3050);
  and g30846 (n16791, \b[42] , n3243);
  and g30847 (n16792, \b[43] , n3045);
  not g30848 (n_14440, n16791);
  not g30849 (n_14441, n16792);
  and g30850 (n16793, n_14440, n_14441);
  not g30851 (n_14442, n16790);
  and g30852 (n16794, n_14442, n16793);
  and g30853 (n16795, n_12601, n16794);
  and g30854 (n16796, n_13499, n16794);
  not g30855 (n_14443, n16795);
  not g30856 (n_14444, n16796);
  and g30857 (n16797, n_14443, n_14444);
  not g30858 (n_14445, n16797);
  and g30859 (n16798, \a[29] , n_14445);
  and g30860 (n16799, n_2476, n16797);
  not g30861 (n_14446, n16798);
  not g30862 (n_14447, n16799);
  and g30863 (n16800, n_14446, n_14447);
  not g30864 (n_14448, n16789);
  not g30865 (n_14449, n16800);
  and g30866 (n16801, n_14448, n_14449);
  not g30867 (n_14450, n16801);
  and g30868 (n16802, n_14448, n_14450);
  and g30869 (n16803, n_14449, n_14450);
  not g30870 (n_14451, n16802);
  not g30871 (n_14452, n16803);
  and g30872 (n16804, n_14451, n_14452);
  not g30873 (n_14453, n16788);
  not g30874 (n_14454, n16804);
  and g30875 (n16805, n_14453, n_14454);
  not g30876 (n_14455, n16805);
  and g30877 (n16806, n_14453, n_14455);
  and g30878 (n16807, n_14454, n_14455);
  not g30879 (n_14456, n16806);
  not g30880 (n_14457, n16807);
  and g30881 (n16808, n_14456, n_14457);
  not g30882 (n_14458, n16578);
  not g30883 (n_14459, n16808);
  and g30884 (n16809, n_14458, n_14459);
  not g30885 (n_14460, n16809);
  and g30886 (n16810, n_14458, n_14460);
  and g30887 (n16811, n_14459, n_14460);
  not g30888 (n_14461, n16810);
  not g30889 (n_14462, n16811);
  and g30890 (n16812, n_14461, n_14462);
  not g30891 (n_14463, n16561);
  and g30892 (n16813, n_14463, n16812);
  not g30893 (n_14464, n16812);
  and g30894 (n16814, n16561, n_14464);
  not g30895 (n_14465, n16813);
  not g30896 (n_14466, n16814);
  and g30897 (n16815, n_14465, n_14466);
  and g30898 (n16816, n_14183, n_14184);
  not g30899 (n_14467, n16816);
  and g30900 (n16817, n_13964, n_14467);
  and g30901 (n16818, \b[53] , n1627);
  and g30902 (n16819, \b[51] , n1763);
  and g30903 (n16820, \b[52] , n1622);
  not g30904 (n_14468, n16819);
  not g30905 (n_14469, n16820);
  and g30906 (n16821, n_14468, n_14469);
  not g30907 (n_14470, n16818);
  and g30908 (n16822, n_14470, n16821);
  not g30909 (n_14471, n1630);
  and g30910 (n16823, n_14471, n16822);
  and g30911 (n16824, n_13261, n16822);
  not g30912 (n_14472, n16823);
  not g30913 (n_14473, n16824);
  and g30914 (n16825, n_14472, n_14473);
  not g30915 (n_14474, n16825);
  and g30916 (n16826, \a[20] , n_14474);
  and g30917 (n16827, n_1221, n16825);
  not g30918 (n_14475, n16826);
  not g30919 (n_14476, n16827);
  and g30920 (n16828, n_14475, n_14476);
  not g30921 (n_14477, n16817);
  not g30922 (n_14478, n16828);
  and g30923 (n16829, n_14477, n_14478);
  not g30924 (n_14479, n16829);
  and g30925 (n16830, n_14477, n_14479);
  and g30926 (n16831, n_14478, n_14479);
  not g30927 (n_14480, n16830);
  not g30928 (n_14481, n16831);
  and g30929 (n16832, n_14480, n_14481);
  not g30930 (n_14482, n16832);
  and g30931 (n16833, n16815, n_14482);
  not g30932 (n_14483, n16833);
  and g30933 (n16834, n16815, n_14483);
  and g30934 (n16835, n_14482, n_14483);
  not g30935 (n_14484, n16834);
  not g30936 (n_14485, n16835);
  and g30937 (n16836, n_14484, n_14485);
  not g30938 (n_14486, n16836);
  and g30939 (n16837, n16546, n_14486);
  not g30940 (n_14487, n16837);
  and g30941 (n16838, n16546, n_14487);
  and g30942 (n16839, n_14486, n_14487);
  not g30943 (n_14488, n16838);
  not g30944 (n_14489, n16839);
  and g30945 (n16840, n_14488, n_14489);
  and g30946 (n16841, \b[59] , n951);
  and g30947 (n16842, \b[57] , n1056);
  and g30948 (n16843, \b[58] , n946);
  and g30954 (n16846, n954, n12179);
  not g30957 (n_14494, n16847);
  and g30958 (n16848, \a[14] , n_14494);
  not g30959 (n_14495, n16848);
  and g30960 (n16849, \a[14] , n_14495);
  and g30961 (n16850, n_14494, n_14495);
  not g30962 (n_14496, n16849);
  not g30963 (n_14497, n16850);
  and g30964 (n16851, n_14496, n_14497);
  and g30965 (n16852, n_13940, n_14194);
  not g30966 (n_14498, n16851);
  not g30967 (n_14499, n16852);
  and g30968 (n16853, n_14498, n_14499);
  not g30969 (n_14500, n16853);
  and g30970 (n16854, n_14498, n_14500);
  and g30971 (n16855, n_14499, n_14500);
  not g30972 (n_14501, n16854);
  not g30973 (n_14502, n16855);
  and g30974 (n16856, n_14501, n_14502);
  not g30975 (n_14503, n16840);
  and g30976 (n16857, n_14503, n16856);
  not g30977 (n_14504, n16856);
  and g30978 (n16858, n16840, n_14504);
  not g30979 (n_14505, n16857);
  not g30980 (n_14506, n16858);
  and g30981 (n16859, n_14505, n_14506);
  and g30982 (n16860, n_13927, n_14195);
  and g30983 (n16861, \b[62] , n700);
  and g30984 (n16862, \b[60] , n767);
  and g30985 (n16863, \b[61] , n695);
  not g30986 (n_14507, n16862);
  not g30987 (n_14508, n16863);
  and g30988 (n16864, n_14507, n_14508);
  not g30989 (n_14509, n16861);
  and g30990 (n16865, n_14509, n16864);
  and g30991 (n16866, n_13159, n16865);
  and g30992 (n16867, n_13538, n16865);
  not g30993 (n_14510, n16866);
  not g30994 (n_14511, n16867);
  and g30995 (n16868, n_14510, n_14511);
  not g30996 (n_14512, n16868);
  and g30997 (n16869, \a[11] , n_14512);
  and g30998 (n16870, n_400, n16868);
  not g30999 (n_14513, n16869);
  not g31000 (n_14514, n16870);
  and g31001 (n16871, n_14513, n_14514);
  not g31002 (n_14515, n16860);
  not g31003 (n_14516, n16871);
  and g31004 (n16872, n_14515, n_14516);
  not g31005 (n_14517, n16872);
  and g31006 (n16873, n_14515, n_14517);
  and g31007 (n16874, n_14516, n_14517);
  not g31008 (n_14518, n16873);
  not g31009 (n_14519, n16874);
  and g31010 (n16875, n_14518, n_14519);
  not g31011 (n_14520, n16859);
  not g31012 (n_14521, n16875);
  and g31013 (n16876, n_14520, n_14521);
  and g31014 (n16877, n16859, n_14519);
  and g31015 (n16878, n_14518, n16877);
  not g31016 (n_14522, n16876);
  not g31017 (n_14523, n16878);
  and g31018 (n16879, n_14522, n_14523);
  not g31019 (n_14524, n16531);
  and g31020 (n16880, n_14524, n16879);
  not g31021 (n_14525, n16879);
  and g31022 (n16881, n16531, n_14525);
  not g31023 (n_14526, n16880);
  not g31024 (n_14527, n16881);
  and g31025 (n16882, n_14526, n_14527);
  not g31026 (n_14528, n16519);
  and g31027 (n16883, n_14528, n16882);
  not g31028 (n_14529, n16883);
  and g31029 (n16884, n_14528, n_14529);
  and g31030 (n16885, n16882, n_14529);
  not g31031 (n_14530, n16884);
  not g31032 (n_14531, n16885);
  and g31033 (n16886, n_14530, n_14531);
  not g31034 (n_14532, n16518);
  not g31035 (n_14533, n16886);
  and g31036 (n16887, n_14532, n_14533);
  and g31037 (n16888, n16518, n_14531);
  and g31038 (n16889, n_14530, n16888);
  not g31039 (n_14534, n16887);
  not g31040 (n_14535, n16889);
  and g31041 (\f[71] , n_14534, n_14535);
  and g31042 (n16891, n_14529, n_14534);
  and g31043 (n16892, n_14223, n_14526);
  and g31044 (n16893, n_14517, n_14522);
  and g31045 (n16894, \b[63] , n700);
  and g31046 (n16895, \b[61] , n767);
  and g31047 (n16896, \b[62] , n695);
  and g31053 (n16899, n703, n13771);
  not g31056 (n_14540, n16900);
  and g31057 (n16901, \a[11] , n_14540);
  not g31058 (n_14541, n16901);
  and g31059 (n16902, \a[11] , n_14541);
  and g31060 (n16903, n_14540, n_14541);
  not g31061 (n_14542, n16902);
  not g31062 (n_14543, n16903);
  and g31063 (n16904, n_14542, n_14543);
  not g31064 (n_14544, n16893);
  not g31065 (n_14545, n16904);
  and g31066 (n16905, n_14544, n_14545);
  not g31067 (n_14546, n16905);
  and g31068 (n16906, n_14544, n_14546);
  and g31069 (n16907, n_14545, n_14546);
  not g31070 (n_14547, n16906);
  not g31071 (n_14548, n16907);
  and g31072 (n16908, n_14547, n_14548);
  and g31073 (n16909, n_14503, n_14504);
  not g31074 (n_14549, n16909);
  and g31075 (n16910, n_14500, n_14549);
  and g31076 (n16911, \b[60] , n951);
  and g31077 (n16912, \b[58] , n1056);
  and g31078 (n16913, \b[59] , n946);
  and g31084 (n16916, n954, n12211);
  not g31087 (n_14554, n16917);
  and g31088 (n16918, \a[14] , n_14554);
  not g31089 (n_14555, n16918);
  and g31090 (n16919, \a[14] , n_14555);
  and g31091 (n16920, n_14554, n_14555);
  not g31092 (n_14556, n16919);
  not g31093 (n_14557, n16920);
  and g31094 (n16921, n_14556, n_14557);
  not g31095 (n_14558, n16910);
  and g31096 (n16922, n_14558, n16921);
  not g31097 (n_14559, n16921);
  and g31098 (n16923, n16910, n_14559);
  not g31099 (n_14560, n16922);
  not g31100 (n_14561, n16923);
  and g31101 (n16924, n_14560, n_14561);
  and g31102 (n16925, \b[57] , n1302);
  and g31103 (n16926, \b[55] , n1391);
  and g31104 (n16927, \b[56] , n1297);
  and g31110 (n16930, n1305, n11410);
  not g31113 (n_14566, n16931);
  and g31114 (n16932, \a[17] , n_14566);
  not g31115 (n_14567, n16932);
  and g31116 (n16933, \a[17] , n_14567);
  and g31117 (n16934, n_14566, n_14567);
  not g31118 (n_14568, n16933);
  not g31119 (n_14569, n16934);
  and g31120 (n16935, n_14568, n_14569);
  and g31121 (n16936, n_14237, n_14487);
  and g31122 (n16937, n16935, n16936);
  not g31123 (n_14570, n16935);
  not g31124 (n_14571, n16936);
  and g31125 (n16938, n_14570, n_14571);
  not g31126 (n_14572, n16937);
  not g31127 (n_14573, n16938);
  and g31128 (n16939, n_14572, n_14573);
  and g31129 (n16940, n_14479, n_14483);
  and g31130 (n16941, \b[54] , n1627);
  and g31131 (n16942, \b[52] , n1763);
  and g31132 (n16943, \b[53] , n1622);
  and g31138 (n16946, n1630, n9998);
  not g31141 (n_14578, n16947);
  and g31142 (n16948, \a[20] , n_14578);
  not g31143 (n_14579, n16948);
  and g31144 (n16949, \a[20] , n_14579);
  and g31145 (n16950, n_14578, n_14579);
  not g31146 (n_14580, n16949);
  not g31147 (n_14581, n16950);
  and g31148 (n16951, n_14580, n_14581);
  not g31149 (n_14582, n16940);
  not g31150 (n_14583, n16951);
  and g31151 (n16952, n_14582, n_14583);
  not g31152 (n_14584, n16952);
  and g31153 (n16953, n_14582, n_14584);
  and g31154 (n16954, n_14583, n_14584);
  not g31155 (n_14585, n16953);
  not g31156 (n_14586, n16954);
  and g31157 (n16955, n_14585, n_14586);
  and g31158 (n16956, \b[48] , n2539);
  and g31159 (n16957, \b[46] , n2685);
  and g31160 (n16958, \b[47] , n2534);
  and g31166 (n16961, n2542, n8009);
  not g31169 (n_14591, n16962);
  and g31170 (n16963, \a[26] , n_14591);
  not g31171 (n_14592, n16963);
  and g31172 (n16964, \a[26] , n_14592);
  and g31173 (n16965, n_14591, n_14592);
  not g31174 (n_14593, n16964);
  not g31175 (n_14594, n16965);
  and g31176 (n16966, n_14593, n_14594);
  and g31177 (n16967, n_14261, n_14460);
  and g31178 (n16968, n16966, n16967);
  not g31179 (n_14595, n16966);
  not g31180 (n_14596, n16967);
  and g31181 (n16969, n_14595, n_14596);
  not g31182 (n_14597, n16968);
  not g31183 (n_14598, n16969);
  and g31184 (n16970, n_14597, n_14598);
  and g31185 (n16971, n_14450, n_14455);
  and g31186 (n16972, \b[45] , n3050);
  and g31187 (n16973, \b[43] , n3243);
  and g31188 (n16974, \b[44] , n3045);
  and g31194 (n16977, n3053, n7361);
  not g31197 (n_14603, n16978);
  and g31198 (n16979, \a[29] , n_14603);
  not g31199 (n_14604, n16979);
  and g31200 (n16980, \a[29] , n_14604);
  and g31201 (n16981, n_14603, n_14604);
  not g31202 (n_14605, n16980);
  not g31203 (n_14606, n16981);
  and g31204 (n16982, n_14605, n_14606);
  not g31205 (n_14607, n16971);
  not g31206 (n_14608, n16982);
  and g31207 (n16983, n_14607, n_14608);
  not g31208 (n_14609, n16983);
  and g31209 (n16984, n_14607, n_14609);
  and g31210 (n16985, n_14608, n_14609);
  not g31211 (n_14610, n16984);
  not g31212 (n_14611, n16985);
  and g31213 (n16986, n_14610, n_14611);
  and g31214 (n16987, n_14275, n_14437);
  and g31215 (n16988, \b[42] , n3638);
  and g31216 (n16989, \b[40] , n3843);
  and g31217 (n16990, \b[41] , n3633);
  and g31223 (n16993, n3641, n6489);
  not g31226 (n_14616, n16994);
  and g31227 (n16995, \a[32] , n_14616);
  not g31228 (n_14617, n16995);
  and g31229 (n16996, \a[32] , n_14617);
  and g31230 (n16997, n_14616, n_14617);
  not g31231 (n_14618, n16996);
  not g31232 (n_14619, n16997);
  and g31233 (n16998, n_14618, n_14619);
  not g31234 (n_14620, n16987);
  not g31235 (n_14621, n16998);
  and g31236 (n16999, n_14620, n_14621);
  not g31237 (n_14622, n16999);
  and g31238 (n17000, n_14620, n_14622);
  and g31239 (n17001, n_14621, n_14622);
  not g31240 (n_14623, n17000);
  not g31241 (n_14624, n17001);
  and g31242 (n17002, n_14623, n_14624);
  and g31243 (n17003, n_14415, n_14418);
  and g31244 (n17004, n_14400, n_14412);
  and g31245 (n17005, n_14384, n_14394);
  and g31246 (n17006, n_14366, n_14371);
  and g31247 (n17007, \b[24] , n8362);
  and g31248 (n17008, \b[22] , n8715);
  and g31249 (n17009, \b[23] , n8357);
  and g31255 (n17012, n2458, n8365);
  not g31258 (n_14629, n17013);
  and g31259 (n17014, \a[50] , n_14629);
  not g31260 (n_14630, n17014);
  and g31261 (n17015, \a[50] , n_14630);
  and g31262 (n17016, n_14629, n_14630);
  not g31263 (n_14631, n17015);
  not g31264 (n_14632, n17016);
  and g31265 (n17017, n_14631, n_14632);
  and g31266 (n17018, \b[18] , n10426);
  and g31267 (n17019, \b[16] , n10796);
  and g31268 (n17020, \b[17] , n10421);
  and g31274 (n17023, n1566, n10429);
  not g31277 (n_14637, n17024);
  and g31278 (n17025, \a[56] , n_14637);
  not g31279 (n_14638, n17025);
  and g31280 (n17026, \a[56] , n_14638);
  and g31281 (n17027, n_14637, n_14638);
  not g31282 (n_14639, n17026);
  not g31283 (n_14640, n17027);
  and g31284 (n17028, n_14639, n_14640);
  and g31285 (n17029, n_14317, n_14318);
  not g31286 (n_14641, n17029);
  and g31287 (n17030, n_14331, n_14641);
  and g31288 (n17031, \b[12] , n12668);
  and g31289 (n17032, \b[10] , n13047);
  and g31290 (n17033, \b[11] , n12663);
  and g31296 (n17036, n842, n12671);
  not g31299 (n_14646, n17037);
  and g31300 (n17038, \a[62] , n_14646);
  not g31301 (n_14647, n17038);
  and g31302 (n17039, \a[62] , n_14647);
  and g31303 (n17040, n_14646, n_14647);
  not g31304 (n_14648, n17039);
  not g31305 (n_14649, n17040);
  and g31306 (n17041, n_14648, n_14649);
  and g31307 (n17042, \b[8] , n13903);
  and g31308 (n17043, \b[9] , n_11555);
  not g31309 (n_14650, n17042);
  not g31310 (n_14651, n17043);
  and g31311 (n17044, n_14650, n_14651);
  and g31312 (n17045, \a[8] , n_14302);
  and g31313 (n17046, n_234, n16633);
  not g31314 (n_14652, n17045);
  not g31315 (n_14653, n17046);
  and g31316 (n17047, n_14652, n_14653);
  not g31317 (n_14654, n17044);
  not g31318 (n_14655, n17047);
  and g31319 (n17048, n_14654, n_14655);
  and g31320 (n17049, n17044, n17047);
  not g31321 (n_14656, n17048);
  not g31322 (n_14657, n17049);
  and g31323 (n17050, n_14656, n_14657);
  not g31324 (n_14658, n16639);
  and g31325 (n17051, n_14658, n17050);
  not g31326 (n_14659, n17050);
  and g31327 (n17052, n16639, n_14659);
  not g31328 (n_14660, n17051);
  not g31329 (n_14661, n17052);
  and g31330 (n17053, n_14660, n_14661);
  and g31331 (n17054, n17041, n17053);
  not g31332 (n_14662, n17041);
  not g31333 (n_14663, n17053);
  and g31334 (n17055, n_14662, n_14663);
  not g31335 (n_14664, n17054);
  not g31336 (n_14665, n17055);
  and g31337 (n17056, n_14664, n_14665);
  and g31338 (n17057, \b[15] , n11531);
  and g31339 (n17058, \b[13] , n11896);
  and g31340 (n17059, \b[14] , n11526);
  and g31346 (n17062, n1131, n11534);
  not g31349 (n_14670, n17063);
  and g31350 (n17064, \a[59] , n_14670);
  not g31351 (n_14671, n17064);
  and g31352 (n17065, \a[59] , n_14671);
  and g31353 (n17066, n_14670, n_14671);
  not g31354 (n_14672, n17065);
  not g31355 (n_14673, n17066);
  and g31356 (n17067, n_14672, n_14673);
  not g31357 (n_14674, n17056);
  not g31358 (n_14675, n17067);
  and g31359 (n17068, n_14674, n_14675);
  and g31360 (n17069, n17056, n17067);
  not g31361 (n_14676, n17068);
  not g31362 (n_14677, n17069);
  and g31363 (n17070, n_14676, n_14677);
  not g31364 (n_14678, n17030);
  and g31365 (n17071, n_14678, n17070);
  not g31366 (n_14679, n17070);
  and g31367 (n17072, n17030, n_14679);
  not g31368 (n_14680, n17071);
  not g31369 (n_14681, n17072);
  and g31370 (n17073, n_14680, n_14681);
  not g31371 (n_14682, n17028);
  and g31372 (n17074, n_14682, n17073);
  not g31373 (n_14683, n17074);
  and g31374 (n17075, n17073, n_14683);
  and g31375 (n17076, n_14682, n_14683);
  not g31376 (n_14684, n17075);
  not g31377 (n_14685, n17076);
  and g31378 (n17077, n_14684, n_14685);
  and g31379 (n17078, n_14336, n_14346);
  and g31380 (n17079, n17077, n17078);
  not g31381 (n_14686, n17077);
  not g31382 (n_14687, n17078);
  and g31383 (n17080, n_14686, n_14687);
  not g31384 (n_14688, n17079);
  not g31385 (n_14689, n17080);
  and g31386 (n17081, n_14688, n_14689);
  and g31387 (n17082, \b[21] , n9339);
  and g31388 (n17083, \b[19] , n9732);
  and g31389 (n17084, \b[20] , n9334);
  and g31395 (n17087, n1984, n9342);
  not g31398 (n_14694, n17088);
  and g31399 (n17089, \a[53] , n_14694);
  not g31400 (n_14695, n17089);
  and g31401 (n17090, \a[53] , n_14695);
  and g31402 (n17091, n_14694, n_14695);
  not g31403 (n_14696, n17090);
  not g31404 (n_14697, n17091);
  and g31405 (n17092, n_14696, n_14697);
  not g31406 (n_14698, n17092);
  and g31407 (n17093, n17081, n_14698);
  not g31408 (n_14699, n17093);
  and g31409 (n17094, n17081, n_14699);
  and g31410 (n17095, n_14698, n_14699);
  not g31411 (n_14700, n17094);
  not g31412 (n_14701, n17095);
  and g31413 (n17096, n_14700, n_14701);
  and g31414 (n17097, n_14352, n_14364);
  not g31415 (n_14702, n17096);
  not g31416 (n_14703, n17097);
  and g31417 (n17098, n_14702, n_14703);
  and g31418 (n17099, n17096, n17097);
  not g31419 (n_14704, n17098);
  not g31420 (n_14705, n17099);
  and g31421 (n17100, n_14704, n_14705);
  not g31422 (n_14706, n17017);
  and g31423 (n17101, n_14706, n17100);
  not g31424 (n_14707, n17101);
  and g31425 (n17102, n_14706, n_14707);
  and g31426 (n17103, n17100, n_14707);
  not g31427 (n_14708, n17102);
  not g31428 (n_14709, n17103);
  and g31429 (n17104, n_14708, n_14709);
  not g31430 (n_14710, n17006);
  not g31431 (n_14711, n17104);
  and g31432 (n17105, n_14710, n_14711);
  not g31433 (n_14712, n17105);
  and g31434 (n17106, n_14710, n_14712);
  and g31435 (n17107, n_14711, n_14712);
  not g31436 (n_14713, n17106);
  not g31437 (n_14714, n17107);
  and g31438 (n17108, n_14713, n_14714);
  and g31439 (n17109, \b[27] , n7446);
  and g31440 (n17110, \b[25] , n7787);
  and g31441 (n17111, \b[26] , n7441);
  and g31447 (n17114, n2990, n7449);
  not g31450 (n_14719, n17115);
  and g31451 (n17116, \a[47] , n_14719);
  not g31452 (n_14720, n17116);
  and g31453 (n17117, \a[47] , n_14720);
  and g31454 (n17118, n_14719, n_14720);
  not g31455 (n_14721, n17117);
  not g31456 (n_14722, n17118);
  and g31457 (n17119, n_14721, n_14722);
  not g31458 (n_14723, n17108);
  not g31459 (n_14724, n17119);
  and g31460 (n17120, n_14723, n_14724);
  not g31461 (n_14725, n17120);
  and g31462 (n17121, n_14723, n_14725);
  and g31463 (n17122, n_14724, n_14725);
  not g31464 (n_14726, n17121);
  not g31465 (n_14727, n17122);
  and g31466 (n17123, n_14726, n_14727);
  and g31467 (n17124, n_14375, n_14378);
  and g31468 (n17125, n17123, n17124);
  not g31469 (n_14728, n17123);
  not g31470 (n_14729, n17124);
  and g31471 (n17126, n_14728, n_14729);
  not g31472 (n_14730, n17125);
  not g31473 (n_14731, n17126);
  and g31474 (n17127, n_14730, n_14731);
  and g31475 (n17128, \b[30] , n6595);
  and g31476 (n17129, \b[28] , n6902);
  and g31477 (n17130, \b[29] , n6590);
  and g31483 (n17133, n3577, n6598);
  not g31486 (n_14736, n17134);
  and g31487 (n17135, \a[44] , n_14736);
  not g31488 (n_14737, n17135);
  and g31489 (n17136, \a[44] , n_14737);
  and g31490 (n17137, n_14736, n_14737);
  not g31491 (n_14738, n17136);
  not g31492 (n_14739, n17137);
  and g31493 (n17138, n_14738, n_14739);
  not g31494 (n_14740, n17138);
  and g31495 (n17139, n17127, n_14740);
  not g31496 (n_14741, n17127);
  and g31497 (n17140, n_14741, n17138);
  not g31498 (n_14742, n17005);
  not g31499 (n_14743, n17140);
  and g31500 (n17141, n_14742, n_14743);
  not g31501 (n_14744, n17139);
  and g31502 (n17142, n_14744, n17141);
  not g31503 (n_14745, n17142);
  and g31504 (n17143, n_14742, n_14745);
  and g31505 (n17144, n_14744, n_14745);
  and g31506 (n17145, n_14743, n17144);
  not g31507 (n_14746, n17143);
  not g31508 (n_14747, n17145);
  and g31509 (n17146, n_14746, n_14747);
  and g31510 (n17147, \b[33] , n5777);
  and g31511 (n17148, \b[31] , n6059);
  and g31512 (n17149, \b[32] , n5772);
  and g31518 (n17152, n4223, n5780);
  not g31521 (n_14752, n17153);
  and g31522 (n17154, \a[41] , n_14752);
  not g31523 (n_14753, n17154);
  and g31524 (n17155, \a[41] , n_14753);
  and g31525 (n17156, n_14752, n_14753);
  not g31526 (n_14754, n17155);
  not g31527 (n_14755, n17156);
  and g31528 (n17157, n_14754, n_14755);
  not g31529 (n_14756, n17146);
  not g31530 (n_14757, n17157);
  and g31531 (n17158, n_14756, n_14757);
  not g31532 (n_14758, n17158);
  and g31533 (n17159, n_14756, n_14758);
  and g31534 (n17160, n_14757, n_14758);
  not g31535 (n_14759, n17159);
  not g31536 (n_14760, n17160);
  and g31537 (n17161, n_14759, n_14760);
  not g31538 (n_14761, n17004);
  and g31539 (n17162, n_14761, n17161);
  not g31540 (n_14762, n17161);
  and g31541 (n17163, n17004, n_14762);
  not g31542 (n_14763, n17162);
  not g31543 (n_14764, n17163);
  and g31544 (n17164, n_14763, n_14764);
  and g31545 (n17165, \b[36] , n5035);
  and g31546 (n17166, \b[34] , n5277);
  and g31547 (n17167, \b[35] , n5030);
  and g31553 (n17170, n4922, n5038);
  not g31556 (n_14769, n17171);
  and g31557 (n17172, \a[38] , n_14769);
  not g31558 (n_14770, n17172);
  and g31559 (n17173, \a[38] , n_14770);
  and g31560 (n17174, n_14769, n_14770);
  not g31561 (n_14771, n17173);
  not g31562 (n_14772, n17174);
  and g31563 (n17175, n_14771, n_14772);
  not g31564 (n_14773, n17164);
  not g31565 (n_14774, n17175);
  and g31566 (n17176, n_14773, n_14774);
  and g31567 (n17177, n17164, n17175);
  not g31568 (n_14775, n17176);
  not g31569 (n_14776, n17177);
  and g31570 (n17178, n_14775, n_14776);
  not g31571 (n_14777, n17178);
  and g31572 (n17179, n17003, n_14777);
  not g31573 (n_14778, n17003);
  and g31574 (n17180, n_14778, n17178);
  not g31575 (n_14779, n17179);
  not g31576 (n_14780, n17180);
  and g31577 (n17181, n_14779, n_14780);
  and g31578 (n17182, \b[39] , n4287);
  and g31579 (n17183, \b[37] , n4532);
  and g31580 (n17184, \b[38] , n4282);
  and g31586 (n17187, n4290, n5451);
  not g31589 (n_14785, n17188);
  and g31590 (n17189, \a[35] , n_14785);
  not g31591 (n_14786, n17189);
  and g31592 (n17190, \a[35] , n_14786);
  and g31593 (n17191, n_14785, n_14786);
  not g31594 (n_14787, n17190);
  not g31595 (n_14788, n17191);
  and g31596 (n17192, n_14787, n_14788);
  not g31597 (n_14789, n17192);
  and g31598 (n17193, n17181, n_14789);
  not g31599 (n_14790, n17193);
  and g31600 (n17194, n17181, n_14790);
  and g31601 (n17195, n_14789, n_14790);
  not g31602 (n_14791, n17194);
  not g31603 (n_14792, n17195);
  and g31604 (n17196, n_14791, n_14792);
  and g31605 (n17197, n_14424, n_14436);
  not g31606 (n_14793, n17196);
  not g31607 (n_14794, n17197);
  and g31608 (n17198, n_14793, n_14794);
  not g31609 (n_14795, n17198);
  and g31610 (n17199, n_14793, n_14795);
  and g31611 (n17200, n_14794, n_14795);
  not g31612 (n_14796, n17199);
  not g31613 (n_14797, n17200);
  and g31614 (n17201, n_14796, n_14797);
  not g31615 (n_14798, n17002);
  not g31616 (n_14799, n17201);
  and g31617 (n17202, n_14798, n_14799);
  not g31618 (n_14800, n17202);
  and g31619 (n17203, n_14798, n_14800);
  and g31620 (n17204, n_14799, n_14800);
  not g31621 (n_14801, n17203);
  not g31622 (n_14802, n17204);
  and g31623 (n17205, n_14801, n_14802);
  not g31624 (n_14803, n16986);
  and g31625 (n17206, n_14803, n17205);
  not g31626 (n_14804, n17205);
  and g31627 (n17207, n16986, n_14804);
  not g31628 (n_14805, n17206);
  not g31629 (n_14806, n17207);
  and g31630 (n17208, n_14805, n_14806);
  not g31631 (n_14807, n17208);
  and g31632 (n17209, n16970, n_14807);
  not g31633 (n_14808, n17209);
  and g31634 (n17210, n16970, n_14808);
  and g31635 (n17211, n_14807, n_14808);
  not g31636 (n_14809, n17210);
  not g31637 (n_14810, n17211);
  and g31638 (n17212, n_14809, n_14810);
  and g31639 (n17213, \b[51] , n2048);
  and g31640 (n17214, \b[49] , n2198);
  and g31641 (n17215, \b[50] , n2043);
  and g31647 (n17218, n2051, n8976);
  not g31650 (n_14815, n17219);
  and g31651 (n17220, \a[23] , n_14815);
  not g31652 (n_14816, n17220);
  and g31653 (n17221, \a[23] , n_14816);
  and g31654 (n17222, n_14815, n_14816);
  not g31655 (n_14817, n17221);
  not g31656 (n_14818, n17222);
  and g31657 (n17223, n_14817, n_14818);
  and g31658 (n17224, n_14249, n_14466);
  not g31659 (n_14819, n17223);
  not g31660 (n_14820, n17224);
  and g31661 (n17225, n_14819, n_14820);
  and g31662 (n17226, n17223, n17224);
  not g31663 (n_14821, n17225);
  not g31664 (n_14822, n17226);
  and g31665 (n17227, n_14821, n_14822);
  not g31666 (n_14823, n17212);
  and g31667 (n17228, n_14823, n17227);
  not g31668 (n_14824, n17228);
  and g31669 (n17229, n_14823, n_14824);
  and g31670 (n17230, n17227, n_14824);
  not g31671 (n_14825, n17229);
  not g31672 (n_14826, n17230);
  and g31673 (n17231, n_14825, n_14826);
  not g31674 (n_14827, n16955);
  not g31675 (n_14828, n17231);
  and g31676 (n17232, n_14827, n_14828);
  not g31677 (n_14829, n17232);
  and g31678 (n17233, n_14827, n_14829);
  and g31679 (n17234, n_14828, n_14829);
  not g31680 (n_14830, n17233);
  not g31681 (n_14831, n17234);
  and g31682 (n17235, n_14830, n_14831);
  not g31683 (n_14832, n17235);
  and g31684 (n17236, n16939, n_14832);
  not g31685 (n_14833, n16939);
  and g31686 (n17237, n_14833, n17235);
  not g31687 (n_14834, n16924);
  not g31688 (n_14835, n17237);
  and g31689 (n17238, n_14834, n_14835);
  not g31690 (n_14836, n17236);
  and g31691 (n17239, n_14836, n17238);
  not g31692 (n_14837, n17239);
  and g31693 (n17240, n_14834, n_14837);
  and g31694 (n17241, n_14835, n_14837);
  and g31695 (n17242, n_14836, n17241);
  not g31696 (n_14838, n17240);
  not g31697 (n_14839, n17242);
  and g31698 (n17243, n_14838, n_14839);
  not g31699 (n_14840, n16908);
  and g31700 (n17244, n_14840, n17243);
  not g31701 (n_14841, n17243);
  and g31702 (n17245, n16908, n_14841);
  not g31703 (n_14842, n17244);
  not g31704 (n_14843, n17245);
  and g31705 (n17246, n_14842, n_14843);
  not g31706 (n_14844, n16892);
  not g31707 (n_14845, n17246);
  and g31708 (n17247, n_14844, n_14845);
  not g31709 (n_14846, n17247);
  and g31710 (n17248, n_14844, n_14846);
  and g31711 (n17249, n_14845, n_14846);
  not g31712 (n_14847, n17248);
  not g31713 (n_14848, n17249);
  and g31714 (n17250, n_14847, n_14848);
  not g31715 (n_14849, n16891);
  not g31716 (n_14850, n17250);
  and g31717 (n17251, n_14849, n_14850);
  and g31718 (n17252, n16891, n_14848);
  and g31719 (n17253, n_14847, n17252);
  not g31720 (n_14851, n17251);
  not g31721 (n_14852, n17253);
  and g31722 (\f[72] , n_14851, n_14852);
  and g31723 (n17255, n_14846, n_14851);
  and g31724 (n17256, n_14840, n_14841);
  not g31725 (n_14853, n17256);
  and g31726 (n17257, n_14546, n_14853);
  and g31727 (n17258, \b[61] , n951);
  and g31728 (n17259, \b[59] , n1056);
  and g31729 (n17260, \b[60] , n946);
  and g31735 (n17263, n954, n12969);
  not g31738 (n_14858, n17264);
  and g31739 (n17265, \a[14] , n_14858);
  not g31740 (n_14859, n17265);
  and g31741 (n17266, \a[14] , n_14859);
  and g31742 (n17267, n_14858, n_14859);
  not g31743 (n_14860, n17266);
  not g31744 (n_14861, n17267);
  and g31745 (n17268, n_14860, n_14861);
  and g31746 (n17269, n_14573, n_14836);
  not g31747 (n_14862, n17268);
  not g31748 (n_14863, n17269);
  and g31749 (n17270, n_14862, n_14863);
  not g31750 (n_14864, n17270);
  and g31751 (n17271, n_14862, n_14864);
  and g31752 (n17272, n_14863, n_14864);
  not g31753 (n_14865, n17271);
  not g31754 (n_14866, n17272);
  and g31755 (n17273, n_14865, n_14866);
  and g31756 (n17274, \b[55] , n1627);
  and g31757 (n17275, \b[53] , n1763);
  and g31758 (n17276, \b[54] , n1622);
  and g31764 (n17279, n1630, n10684);
  not g31767 (n_14871, n17280);
  and g31768 (n17281, \a[20] , n_14871);
  not g31769 (n_14872, n17281);
  and g31770 (n17282, \a[20] , n_14872);
  and g31771 (n17283, n_14871, n_14872);
  not g31772 (n_14873, n17282);
  not g31773 (n_14874, n17283);
  and g31774 (n17284, n_14873, n_14874);
  and g31775 (n17285, n_14821, n_14824);
  and g31776 (n17286, n17284, n17285);
  not g31777 (n_14875, n17284);
  not g31778 (n_14876, n17285);
  and g31779 (n17287, n_14875, n_14876);
  not g31780 (n_14877, n17286);
  not g31781 (n_14878, n17287);
  and g31782 (n17288, n_14877, n_14878);
  and g31783 (n17289, \b[52] , n2048);
  and g31784 (n17290, \b[50] , n2198);
  and g31785 (n17291, \b[51] , n2043);
  and g31791 (n17294, n2051, n9628);
  not g31794 (n_14883, n17295);
  and g31795 (n17296, \a[23] , n_14883);
  not g31796 (n_14884, n17296);
  and g31797 (n17297, \a[23] , n_14884);
  and g31798 (n17298, n_14883, n_14884);
  not g31799 (n_14885, n17297);
  not g31800 (n_14886, n17298);
  and g31801 (n17299, n_14885, n_14886);
  and g31802 (n17300, n_14598, n_14808);
  and g31803 (n17301, n17299, n17300);
  not g31804 (n_14887, n17299);
  not g31805 (n_14888, n17300);
  and g31806 (n17302, n_14887, n_14888);
  not g31807 (n_14889, n17301);
  not g31808 (n_14890, n17302);
  and g31809 (n17303, n_14889, n_14890);
  and g31810 (n17304, \b[49] , n2539);
  and g31811 (n17305, \b[47] , n2685);
  and g31812 (n17306, \b[48] , n2534);
  and g31818 (n17309, n2542, n8625);
  not g31821 (n_14895, n17310);
  and g31822 (n17311, \a[26] , n_14895);
  not g31823 (n_14896, n17311);
  and g31824 (n17312, \a[26] , n_14896);
  and g31825 (n17313, n_14895, n_14896);
  not g31826 (n_14897, n17312);
  not g31827 (n_14898, n17313);
  and g31828 (n17314, n_14897, n_14898);
  and g31829 (n17315, n_14803, n_14804);
  not g31830 (n_14899, n17315);
  and g31831 (n17316, n_14609, n_14899);
  not g31832 (n_14900, n17314);
  not g31833 (n_14901, n17316);
  and g31834 (n17317, n_14900, n_14901);
  not g31835 (n_14902, n17317);
  and g31836 (n17318, n_14900, n_14902);
  and g31837 (n17319, n_14901, n_14902);
  not g31838 (n_14903, n17318);
  not g31839 (n_14904, n17319);
  and g31840 (n17320, n_14903, n_14904);
  and g31841 (n17321, \b[43] , n3638);
  and g31842 (n17322, \b[41] , n3843);
  and g31843 (n17323, \b[42] , n3633);
  and g31849 (n17326, n3641, n6515);
  not g31852 (n_14909, n17327);
  and g31853 (n17328, \a[32] , n_14909);
  not g31854 (n_14910, n17328);
  and g31855 (n17329, \a[32] , n_14910);
  and g31856 (n17330, n_14909, n_14910);
  not g31857 (n_14911, n17329);
  not g31858 (n_14912, n17330);
  and g31859 (n17331, n_14911, n_14912);
  and g31860 (n17332, n_14790, n_14795);
  and g31861 (n17333, n17331, n17332);
  not g31862 (n_14913, n17331);
  not g31863 (n_14914, n17332);
  and g31864 (n17334, n_14913, n_14914);
  not g31865 (n_14915, n17333);
  not g31866 (n_14916, n17334);
  and g31867 (n17335, n_14915, n_14916);
  and g31868 (n17336, \b[40] , n4287);
  and g31869 (n17337, \b[38] , n4532);
  and g31870 (n17338, \b[39] , n4282);
  and g31876 (n17341, n4290, n5955);
  not g31879 (n_14921, n17342);
  and g31880 (n17343, \a[35] , n_14921);
  not g31881 (n_14922, n17343);
  and g31882 (n17344, \a[35] , n_14922);
  and g31883 (n17345, n_14921, n_14922);
  not g31884 (n_14923, n17344);
  not g31885 (n_14924, n17345);
  and g31886 (n17346, n_14923, n_14924);
  and g31887 (n17347, n_14775, n_14780);
  and g31888 (n17348, \b[37] , n5035);
  and g31889 (n17349, \b[35] , n5277);
  and g31890 (n17350, \b[36] , n5030);
  and g31896 (n17353, n5038, n5181);
  not g31899 (n_14929, n17354);
  and g31900 (n17355, \a[38] , n_14929);
  not g31901 (n_14930, n17355);
  and g31902 (n17356, \a[38] , n_14930);
  and g31903 (n17357, n_14929, n_14930);
  not g31904 (n_14931, n17356);
  not g31905 (n_14932, n17357);
  and g31906 (n17358, n_14931, n_14932);
  and g31907 (n17359, n_14761, n_14762);
  not g31908 (n_14933, n17359);
  and g31909 (n17360, n_14758, n_14933);
  and g31910 (n17361, \b[34] , n5777);
  and g31911 (n17362, \b[32] , n6059);
  and g31912 (n17363, \b[33] , n5772);
  and g31918 (n17366, n4466, n5780);
  not g31921 (n_14938, n17367);
  and g31922 (n17368, \a[41] , n_14938);
  not g31923 (n_14939, n17368);
  and g31924 (n17369, \a[41] , n_14939);
  and g31925 (n17370, n_14938, n_14939);
  not g31926 (n_14940, n17369);
  not g31927 (n_14941, n17370);
  and g31928 (n17371, n_14940, n_14941);
  and g31929 (n17372, \b[13] , n12668);
  and g31930 (n17373, \b[11] , n13047);
  and g31931 (n17374, \b[12] , n12663);
  and g31937 (n17377, n1008, n12671);
  not g31940 (n_14946, n17378);
  and g31941 (n17379, \a[62] , n_14946);
  not g31942 (n_14947, n17379);
  and g31943 (n17380, \a[62] , n_14947);
  and g31944 (n17381, n_14946, n_14947);
  not g31945 (n_14948, n17380);
  not g31946 (n_14949, n17381);
  and g31947 (n17382, n_14948, n_14949);
  and g31948 (n17383, \b[9] , n13903);
  and g31949 (n17384, \b[10] , n_11555);
  not g31950 (n_14950, n17383);
  not g31951 (n_14951, n17384);
  and g31952 (n17385, n_14950, n_14951);
  and g31953 (n17386, n_234, n_14302);
  not g31954 (n_14952, n17386);
  and g31955 (n17387, n_14656, n_14952);
  not g31956 (n_14953, n17387);
  and g31957 (n17388, n17385, n_14953);
  not g31958 (n_14954, n17388);
  and g31959 (n17389, n17385, n_14954);
  and g31960 (n17390, n_14953, n_14954);
  not g31961 (n_14955, n17389);
  not g31962 (n_14956, n17390);
  and g31963 (n17391, n_14955, n_14956);
  not g31964 (n_14957, n17382);
  not g31965 (n_14958, n17391);
  and g31966 (n17392, n_14957, n_14958);
  not g31967 (n_14959, n17392);
  and g31968 (n17393, n_14957, n_14959);
  and g31969 (n17394, n_14958, n_14959);
  not g31970 (n_14960, n17393);
  not g31971 (n_14961, n17394);
  and g31972 (n17395, n_14960, n_14961);
  and g31973 (n17396, n_14662, n17053);
  not g31974 (n_14962, n17396);
  and g31975 (n17397, n_14660, n_14962);
  not g31976 (n_14963, n17395);
  not g31977 (n_14964, n17397);
  and g31978 (n17398, n_14963, n_14964);
  not g31979 (n_14965, n17398);
  and g31980 (n17399, n_14963, n_14965);
  and g31981 (n17400, n_14964, n_14965);
  not g31982 (n_14966, n17399);
  not g31983 (n_14967, n17400);
  and g31984 (n17401, n_14966, n_14967);
  and g31985 (n17402, \b[16] , n11531);
  and g31986 (n17403, \b[14] , n11896);
  and g31987 (n17404, \b[15] , n11526);
  and g31993 (n17407, n1237, n11534);
  not g31996 (n_14972, n17408);
  and g31997 (n17409, \a[59] , n_14972);
  not g31998 (n_14973, n17409);
  and g31999 (n17410, \a[59] , n_14973);
  and g32000 (n17411, n_14972, n_14973);
  not g32001 (n_14974, n17410);
  not g32002 (n_14975, n17411);
  and g32003 (n17412, n_14974, n_14975);
  not g32004 (n_14976, n17401);
  not g32005 (n_14977, n17412);
  and g32006 (n17413, n_14976, n_14977);
  not g32007 (n_14978, n17413);
  and g32008 (n17414, n_14976, n_14978);
  and g32009 (n17415, n_14977, n_14978);
  not g32010 (n_14979, n17414);
  not g32011 (n_14980, n17415);
  and g32012 (n17416, n_14979, n_14980);
  and g32013 (n17417, n_14676, n_14680);
  and g32014 (n17418, n17416, n17417);
  not g32015 (n_14981, n17416);
  not g32016 (n_14982, n17417);
  and g32017 (n17419, n_14981, n_14982);
  not g32018 (n_14983, n17418);
  not g32019 (n_14984, n17419);
  and g32020 (n17420, n_14983, n_14984);
  and g32021 (n17421, \b[19] , n10426);
  and g32022 (n17422, \b[17] , n10796);
  and g32023 (n17423, \b[18] , n10421);
  and g32029 (n17426, n1708, n10429);
  not g32032 (n_14989, n17427);
  and g32033 (n17428, \a[56] , n_14989);
  not g32034 (n_14990, n17428);
  and g32035 (n17429, \a[56] , n_14990);
  and g32036 (n17430, n_14989, n_14990);
  not g32037 (n_14991, n17429);
  not g32038 (n_14992, n17430);
  and g32039 (n17431, n_14991, n_14992);
  not g32040 (n_14993, n17431);
  and g32041 (n17432, n17420, n_14993);
  not g32042 (n_14994, n17432);
  and g32043 (n17433, n17420, n_14994);
  and g32044 (n17434, n_14993, n_14994);
  not g32045 (n_14995, n17433);
  not g32046 (n_14996, n17434);
  and g32047 (n17435, n_14995, n_14996);
  and g32048 (n17436, n_14683, n_14689);
  and g32049 (n17437, n17435, n17436);
  not g32050 (n_14997, n17435);
  not g32051 (n_14998, n17436);
  and g32052 (n17438, n_14997, n_14998);
  not g32053 (n_14999, n17437);
  not g32054 (n_15000, n17438);
  and g32055 (n17439, n_14999, n_15000);
  and g32056 (n17440, \b[22] , n9339);
  and g32057 (n17441, \b[20] , n9732);
  and g32058 (n17442, \b[21] , n9334);
  and g32064 (n17445, n2145, n9342);
  not g32067 (n_15005, n17446);
  and g32068 (n17447, \a[53] , n_15005);
  not g32069 (n_15006, n17447);
  and g32070 (n17448, \a[53] , n_15006);
  and g32071 (n17449, n_15005, n_15006);
  not g32072 (n_15007, n17448);
  not g32073 (n_15008, n17449);
  and g32074 (n17450, n_15007, n_15008);
  not g32075 (n_15009, n17450);
  and g32076 (n17451, n17439, n_15009);
  not g32077 (n_15010, n17451);
  and g32078 (n17452, n17439, n_15010);
  and g32079 (n17453, n_15009, n_15010);
  not g32080 (n_15011, n17452);
  not g32081 (n_15012, n17453);
  and g32082 (n17454, n_15011, n_15012);
  and g32083 (n17455, n_14699, n_14704);
  and g32084 (n17456, n17454, n17455);
  not g32085 (n_15013, n17454);
  not g32086 (n_15014, n17455);
  and g32087 (n17457, n_15013, n_15014);
  not g32088 (n_15015, n17456);
  not g32089 (n_15016, n17457);
  and g32090 (n17458, n_15015, n_15016);
  and g32091 (n17459, \b[25] , n8362);
  and g32092 (n17460, \b[23] , n8715);
  and g32093 (n17461, \b[24] , n8357);
  and g32099 (n17464, n2485, n8365);
  not g32102 (n_15021, n17465);
  and g32103 (n17466, \a[50] , n_15021);
  not g32104 (n_15022, n17466);
  and g32105 (n17467, \a[50] , n_15022);
  and g32106 (n17468, n_15021, n_15022);
  not g32107 (n_15023, n17467);
  not g32108 (n_15024, n17468);
  and g32109 (n17469, n_15023, n_15024);
  not g32110 (n_15025, n17469);
  and g32111 (n17470, n17458, n_15025);
  not g32112 (n_15026, n17470);
  and g32113 (n17471, n17458, n_15026);
  and g32114 (n17472, n_15025, n_15026);
  not g32115 (n_15027, n17471);
  not g32116 (n_15028, n17472);
  and g32117 (n17473, n_15027, n_15028);
  and g32118 (n17474, n_14707, n_14712);
  and g32119 (n17475, n17473, n17474);
  not g32120 (n_15029, n17473);
  not g32121 (n_15030, n17474);
  and g32122 (n17476, n_15029, n_15030);
  not g32123 (n_15031, n17475);
  not g32124 (n_15032, n17476);
  and g32125 (n17477, n_15031, n_15032);
  and g32126 (n17478, \b[28] , n7446);
  and g32127 (n17479, \b[26] , n7787);
  and g32128 (n17480, \b[27] , n7441);
  and g32134 (n17483, n3189, n7449);
  not g32137 (n_15037, n17484);
  and g32138 (n17485, \a[47] , n_15037);
  not g32139 (n_15038, n17485);
  and g32140 (n17486, \a[47] , n_15038);
  and g32141 (n17487, n_15037, n_15038);
  not g32142 (n_15039, n17486);
  not g32143 (n_15040, n17487);
  and g32144 (n17488, n_15039, n_15040);
  not g32145 (n_15041, n17488);
  and g32146 (n17489, n17477, n_15041);
  not g32147 (n_15042, n17489);
  and g32148 (n17490, n17477, n_15042);
  and g32149 (n17491, n_15041, n_15042);
  not g32150 (n_15043, n17490);
  not g32151 (n_15044, n17491);
  and g32152 (n17492, n_15043, n_15044);
  and g32153 (n17493, n_14725, n_14731);
  and g32154 (n17494, n17492, n17493);
  not g32155 (n_15045, n17492);
  not g32156 (n_15046, n17493);
  and g32157 (n17495, n_15045, n_15046);
  not g32158 (n_15047, n17494);
  not g32159 (n_15048, n17495);
  and g32160 (n17496, n_15047, n_15048);
  and g32161 (n17497, \b[31] , n6595);
  and g32162 (n17498, \b[29] , n6902);
  and g32163 (n17499, \b[30] , n6590);
  and g32169 (n17502, n3796, n6598);
  not g32172 (n_15053, n17503);
  and g32173 (n17504, \a[44] , n_15053);
  not g32174 (n_15054, n17504);
  and g32175 (n17505, \a[44] , n_15054);
  and g32176 (n17506, n_15053, n_15054);
  not g32177 (n_15055, n17505);
  not g32178 (n_15056, n17506);
  and g32179 (n17507, n_15055, n_15056);
  not g32180 (n_15057, n17496);
  and g32181 (n17508, n_15057, n17507);
  not g32182 (n_15058, n17507);
  and g32183 (n17509, n17496, n_15058);
  not g32184 (n_15059, n17508);
  not g32185 (n_15060, n17509);
  and g32186 (n17510, n_15059, n_15060);
  not g32187 (n_15061, n17144);
  and g32188 (n17511, n_15061, n17510);
  not g32189 (n_15062, n17510);
  and g32190 (n17512, n17144, n_15062);
  not g32191 (n_15063, n17511);
  not g32192 (n_15064, n17512);
  and g32193 (n17513, n_15063, n_15064);
  not g32194 (n_15065, n17371);
  and g32195 (n17514, n_15065, n17513);
  not g32196 (n_15066, n17513);
  and g32197 (n17515, n17371, n_15066);
  not g32198 (n_15067, n17514);
  not g32199 (n_15068, n17515);
  and g32200 (n17516, n_15067, n_15068);
  not g32201 (n_15069, n17360);
  and g32202 (n17517, n_15069, n17516);
  not g32203 (n_15070, n17517);
  and g32204 (n17518, n_15069, n_15070);
  and g32205 (n17519, n17516, n_15070);
  not g32206 (n_15071, n17518);
  not g32207 (n_15072, n17519);
  and g32208 (n17520, n_15071, n_15072);
  not g32209 (n_15073, n17358);
  not g32210 (n_15074, n17520);
  and g32211 (n17521, n_15073, n_15074);
  and g32212 (n17522, n17358, n_15072);
  and g32213 (n17523, n_15071, n17522);
  not g32214 (n_15075, n17521);
  not g32215 (n_15076, n17523);
  and g32216 (n17524, n_15075, n_15076);
  not g32217 (n_15077, n17347);
  and g32218 (n17525, n_15077, n17524);
  not g32219 (n_15078, n17525);
  and g32220 (n17526, n_15077, n_15078);
  and g32221 (n17527, n17524, n_15078);
  not g32222 (n_15079, n17526);
  not g32223 (n_15080, n17527);
  and g32224 (n17528, n_15079, n_15080);
  not g32225 (n_15081, n17346);
  not g32226 (n_15082, n17528);
  and g32227 (n17529, n_15081, n_15082);
  not g32228 (n_15083, n17529);
  and g32229 (n17530, n_15081, n_15083);
  and g32230 (n17531, n_15082, n_15083);
  not g32231 (n_15084, n17530);
  not g32232 (n_15085, n17531);
  and g32233 (n17532, n_15084, n_15085);
  not g32234 (n_15086, n17532);
  and g32235 (n17533, n17335, n_15086);
  not g32236 (n_15087, n17533);
  and g32237 (n17534, n17335, n_15087);
  and g32238 (n17535, n_15086, n_15087);
  not g32239 (n_15088, n17534);
  not g32240 (n_15089, n17535);
  and g32241 (n17536, n_15088, n_15089);
  and g32242 (n17537, n_14622, n_14800);
  and g32243 (n17538, \b[46] , n3050);
  and g32244 (n17539, \b[44] , n3243);
  and g32245 (n17540, \b[45] , n3045);
  not g32246 (n_15090, n17539);
  not g32247 (n_15091, n17540);
  and g32248 (n17541, n_15090, n_15091);
  not g32249 (n_15092, n17538);
  and g32250 (n17542, n_15092, n17541);
  and g32251 (n17543, n_12601, n17542);
  and g32252 (n17544, n_13970, n17542);
  not g32253 (n_15093, n17543);
  not g32254 (n_15094, n17544);
  and g32255 (n17545, n_15093, n_15094);
  not g32256 (n_15095, n17545);
  and g32257 (n17546, \a[29] , n_15095);
  and g32258 (n17547, n_2476, n17545);
  not g32259 (n_15096, n17546);
  not g32260 (n_15097, n17547);
  and g32261 (n17548, n_15096, n_15097);
  not g32262 (n_15098, n17537);
  not g32263 (n_15099, n17548);
  and g32264 (n17549, n_15098, n_15099);
  not g32265 (n_15100, n17549);
  and g32266 (n17550, n_15098, n_15100);
  and g32267 (n17551, n_15099, n_15100);
  not g32268 (n_15101, n17550);
  not g32269 (n_15102, n17551);
  and g32270 (n17552, n_15101, n_15102);
  not g32271 (n_15103, n17536);
  not g32272 (n_15104, n17552);
  and g32273 (n17553, n_15103, n_15104);
  not g32274 (n_15105, n17553);
  and g32275 (n17554, n_15103, n_15105);
  and g32276 (n17555, n_15104, n_15105);
  not g32277 (n_15106, n17554);
  not g32278 (n_15107, n17555);
  and g32279 (n17556, n_15106, n_15107);
  not g32280 (n_15108, n17320);
  not g32281 (n_15109, n17556);
  and g32282 (n17557, n_15108, n_15109);
  not g32283 (n_15110, n17557);
  and g32284 (n17558, n_15108, n_15110);
  and g32285 (n17559, n_15109, n_15110);
  not g32286 (n_15111, n17558);
  not g32287 (n_15112, n17559);
  and g32288 (n17560, n_15111, n_15112);
  not g32289 (n_15113, n17560);
  and g32290 (n17561, n17303, n_15113);
  not g32291 (n_15114, n17303);
  and g32292 (n17562, n_15114, n17560);
  not g32293 (n_15115, n17562);
  and g32294 (n17563, n17288, n_15115);
  not g32295 (n_15116, n17561);
  and g32296 (n17564, n_15116, n17563);
  not g32297 (n_15117, n17564);
  and g32298 (n17565, n17288, n_15117);
  and g32299 (n17566, n_15115, n_15117);
  and g32300 (n17567, n_15116, n17566);
  not g32301 (n_15118, n17565);
  not g32302 (n_15119, n17567);
  and g32303 (n17568, n_15118, n_15119);
  and g32304 (n17569, n_14584, n_14829);
  and g32305 (n17570, \b[58] , n1302);
  and g32306 (n17571, \b[56] , n1391);
  and g32307 (n17572, \b[57] , n1297);
  not g32308 (n_15120, n17571);
  not g32309 (n_15121, n17572);
  and g32310 (n17573, n_15120, n_15121);
  not g32311 (n_15122, n17570);
  and g32312 (n17574, n_15122, n17573);
  and g32313 (n17575, n_13260, n17574);
  and g32314 (n17576, n_13160, n17574);
  not g32315 (n_15123, n17575);
  not g32316 (n_15124, n17576);
  and g32317 (n17577, n_15123, n_15124);
  not g32318 (n_15125, n17577);
  and g32319 (n17578, \a[17] , n_15125);
  and g32320 (n17579, n_926, n17577);
  not g32321 (n_15126, n17578);
  not g32322 (n_15127, n17579);
  and g32323 (n17580, n_15126, n_15127);
  not g32324 (n_15128, n17569);
  not g32325 (n_15129, n17580);
  and g32326 (n17581, n_15128, n_15129);
  not g32327 (n_15130, n17581);
  and g32328 (n17582, n_15128, n_15130);
  and g32329 (n17583, n_15129, n_15130);
  not g32330 (n_15131, n17582);
  not g32331 (n_15132, n17583);
  and g32332 (n17584, n_15131, n_15132);
  not g32333 (n_15133, n17568);
  not g32334 (n_15134, n17584);
  and g32335 (n17585, n_15133, n_15134);
  not g32336 (n_15135, n17585);
  and g32337 (n17586, n_15133, n_15135);
  and g32338 (n17587, n_15134, n_15135);
  not g32339 (n_15136, n17586);
  not g32340 (n_15137, n17587);
  and g32341 (n17588, n_15136, n_15137);
  not g32342 (n_15138, n17273);
  not g32343 (n_15139, n17588);
  and g32344 (n17589, n_15138, n_15139);
  not g32345 (n_15140, n17589);
  and g32346 (n17590, n_15138, n_15140);
  and g32347 (n17591, n_15139, n_15140);
  not g32348 (n_15141, n17590);
  not g32349 (n_15142, n17591);
  and g32350 (n17592, n_15141, n_15142);
  and g32351 (n17593, n_14558, n_14559);
  not g32352 (n_15143, n17593);
  and g32353 (n17594, n_14837, n_15143);
  and g32354 (n17595, \b[62] , n767);
  and g32355 (n17596, \b[63] , n695);
  not g32356 (n_15144, n17595);
  not g32357 (n_15145, n17596);
  and g32358 (n17597, n_15144, n_15145);
  and g32359 (n17598, n_13159, n17597);
  and g32360 (n17599, n13800, n17597);
  not g32361 (n_15146, n17598);
  not g32362 (n_15147, n17599);
  and g32363 (n17600, n_15146, n_15147);
  not g32364 (n_15148, n17600);
  and g32365 (n17601, \a[11] , n_15148);
  and g32366 (n17602, n_400, n17600);
  not g32367 (n_15149, n17601);
  not g32368 (n_15150, n17602);
  and g32369 (n17603, n_15149, n_15150);
  not g32370 (n_15151, n17594);
  not g32371 (n_15152, n17603);
  and g32372 (n17604, n_15151, n_15152);
  not g32373 (n_15153, n17604);
  and g32374 (n17605, n_15151, n_15153);
  and g32375 (n17606, n_15152, n_15153);
  not g32376 (n_15154, n17605);
  not g32377 (n_15155, n17606);
  and g32378 (n17607, n_15154, n_15155);
  not g32379 (n_15156, n17592);
  not g32380 (n_15157, n17607);
  and g32381 (n17608, n_15156, n_15157);
  and g32382 (n17609, n17592, n_15155);
  and g32383 (n17610, n_15154, n17609);
  not g32384 (n_15158, n17608);
  not g32385 (n_15159, n17610);
  and g32386 (n17611, n_15158, n_15159);
  not g32387 (n_15160, n17257);
  and g32388 (n17612, n_15160, n17611);
  not g32389 (n_15161, n17612);
  and g32390 (n17613, n_15160, n_15161);
  and g32391 (n17614, n17611, n_15161);
  not g32392 (n_15162, n17613);
  not g32393 (n_15163, n17614);
  and g32394 (n17615, n_15162, n_15163);
  not g32395 (n_15164, n17255);
  not g32396 (n_15165, n17615);
  and g32397 (n17616, n_15164, n_15165);
  and g32398 (n17617, n17255, n_15163);
  and g32399 (n17618, n_15162, n17617);
  not g32400 (n_15166, n17616);
  not g32401 (n_15167, n17618);
  and g32402 (\f[73] , n_15166, n_15167);
  and g32403 (n17620, n_15161, n_15166);
  and g32404 (n17621, n_15153, n_15158);
  and g32405 (n17622, n_14864, n_15140);
  and g32406 (n17623, \b[63] , n767);
  and g32407 (n17624, n703, n13797);
  not g32408 (n_15168, n17623);
  not g32409 (n_15169, n17624);
  and g32410 (n17625, n_15168, n_15169);
  not g32411 (n_15170, n17625);
  and g32412 (n17626, \a[11] , n_15170);
  not g32413 (n_15171, n17626);
  and g32414 (n17627, \a[11] , n_15171);
  and g32415 (n17628, n_15170, n_15171);
  not g32416 (n_15172, n17627);
  not g32417 (n_15173, n17628);
  and g32418 (n17629, n_15172, n_15173);
  not g32419 (n_15174, n17622);
  not g32420 (n_15175, n17629);
  and g32421 (n17630, n_15174, n_15175);
  not g32422 (n_15176, n17630);
  and g32423 (n17631, n_15174, n_15176);
  and g32424 (n17632, n_15175, n_15176);
  not g32425 (n_15177, n17631);
  not g32426 (n_15178, n17632);
  and g32427 (n17633, n_15177, n_15178);
  and g32428 (n17634, n_15130, n_15135);
  and g32429 (n17635, \b[62] , n951);
  and g32430 (n17636, \b[60] , n1056);
  and g32431 (n17637, \b[61] , n946);
  not g32432 (n_15179, n17636);
  not g32433 (n_15180, n17637);
  and g32434 (n17638, n_15179, n_15180);
  not g32435 (n_15181, n17635);
  and g32436 (n17639, n_15181, n17638);
  and g32437 (n17640, n_12819, n17639);
  and g32438 (n17641, n_13538, n17639);
  not g32439 (n_15182, n17640);
  not g32440 (n_15183, n17641);
  and g32441 (n17642, n_15182, n_15183);
  not g32442 (n_15184, n17642);
  and g32443 (n17643, \a[14] , n_15184);
  and g32444 (n17644, n_623, n17642);
  not g32445 (n_15185, n17643);
  not g32446 (n_15186, n17644);
  and g32447 (n17645, n_15185, n_15186);
  not g32448 (n_15187, n17634);
  not g32449 (n_15188, n17645);
  and g32450 (n17646, n_15187, n_15188);
  and g32451 (n17647, n17634, n17645);
  not g32452 (n_15189, n17646);
  not g32453 (n_15190, n17647);
  and g32454 (n17648, n_15189, n_15190);
  and g32455 (n17649, \b[59] , n1302);
  and g32456 (n17650, \b[57] , n1391);
  and g32457 (n17651, \b[58] , n1297);
  and g32463 (n17654, n1305, n12179);
  not g32466 (n_15195, n17655);
  and g32467 (n17656, \a[17] , n_15195);
  not g32468 (n_15196, n17656);
  and g32469 (n17657, \a[17] , n_15196);
  and g32470 (n17658, n_15195, n_15196);
  not g32471 (n_15197, n17657);
  not g32472 (n_15198, n17658);
  and g32473 (n17659, n_15197, n_15198);
  and g32474 (n17660, n_14878, n_15117);
  and g32475 (n17661, n17659, n17660);
  not g32476 (n_15199, n17659);
  not g32477 (n_15200, n17660);
  and g32478 (n17662, n_15199, n_15200);
  not g32479 (n_15201, n17661);
  not g32480 (n_15202, n17662);
  and g32481 (n17663, n_15201, n_15202);
  and g32482 (n17664, \b[56] , n1627);
  and g32483 (n17665, \b[54] , n1763);
  and g32484 (n17666, \b[55] , n1622);
  and g32490 (n17669, n1630, n10708);
  not g32493 (n_15207, n17670);
  and g32494 (n17671, \a[20] , n_15207);
  not g32495 (n_15208, n17671);
  and g32496 (n17672, \a[20] , n_15208);
  and g32497 (n17673, n_15207, n_15208);
  not g32498 (n_15209, n17672);
  not g32499 (n_15210, n17673);
  and g32500 (n17674, n_15209, n_15210);
  and g32501 (n17675, n_14890, n_15116);
  not g32502 (n_15211, n17674);
  not g32503 (n_15212, n17675);
  and g32504 (n17676, n_15211, n_15212);
  not g32505 (n_15213, n17676);
  and g32506 (n17677, n_15211, n_15213);
  and g32507 (n17678, n_15212, n_15213);
  not g32508 (n_15214, n17677);
  not g32509 (n_15215, n17678);
  and g32510 (n17679, n_15214, n_15215);
  and g32511 (n17680, n_15100, n_15105);
  and g32512 (n17681, \b[50] , n2539);
  and g32513 (n17682, \b[48] , n2685);
  and g32514 (n17683, \b[49] , n2534);
  not g32515 (n_15216, n17682);
  not g32516 (n_15217, n17683);
  and g32517 (n17684, n_15216, n_15217);
  not g32518 (n_15218, n17681);
  and g32519 (n17685, n_15218, n17684);
  and g32520 (n17686, n_13498, n17685);
  not g32521 (n_15219, n8949);
  and g32522 (n17687, n_15219, n17685);
  not g32523 (n_15220, n17686);
  not g32524 (n_15221, n17687);
  and g32525 (n17688, n_15220, n_15221);
  not g32526 (n_15222, n17688);
  and g32527 (n17689, \a[26] , n_15222);
  and g32528 (n17690, n_2025, n17688);
  not g32529 (n_15223, n17689);
  not g32530 (n_15224, n17690);
  and g32531 (n17691, n_15223, n_15224);
  not g32532 (n_15225, n17680);
  not g32533 (n_15226, n17691);
  and g32534 (n17692, n_15225, n_15226);
  and g32535 (n17693, n17680, n17691);
  not g32536 (n_15227, n17692);
  not g32537 (n_15228, n17693);
  and g32538 (n17694, n_15227, n_15228);
  and g32539 (n17695, \b[47] , n3050);
  and g32540 (n17696, \b[45] , n3243);
  and g32541 (n17697, \b[46] , n3045);
  and g32547 (n17700, n3053, n7703);
  not g32550 (n_15233, n17701);
  and g32551 (n17702, \a[29] , n_15233);
  not g32552 (n_15234, n17702);
  and g32553 (n17703, \a[29] , n_15234);
  and g32554 (n17704, n_15233, n_15234);
  not g32555 (n_15235, n17703);
  not g32556 (n_15236, n17704);
  and g32557 (n17705, n_15235, n_15236);
  and g32558 (n17706, n_14916, n_15087);
  and g32559 (n17707, n17705, n17706);
  not g32560 (n_15237, n17705);
  not g32561 (n_15238, n17706);
  and g32562 (n17708, n_15237, n_15238);
  not g32563 (n_15239, n17707);
  not g32564 (n_15240, n17708);
  and g32565 (n17709, n_15239, n_15240);
  and g32566 (n17710, n_15078, n_15083);
  and g32567 (n17711, \b[44] , n3638);
  and g32568 (n17712, \b[42] , n3843);
  and g32569 (n17713, \b[43] , n3633);
  not g32570 (n_15241, n17712);
  not g32571 (n_15242, n17713);
  and g32572 (n17714, n_15241, n_15242);
  not g32573 (n_15243, n17711);
  and g32574 (n17715, n_15243, n17714);
  and g32575 (n17716, n_12780, n17715);
  and g32576 (n17717, n_13499, n17715);
  not g32577 (n_15244, n17716);
  not g32578 (n_15245, n17717);
  and g32579 (n17718, n_15244, n_15245);
  not g32580 (n_15246, n17718);
  and g32581 (n17719, \a[32] , n_15246);
  and g32582 (n17720, n_2992, n17718);
  not g32583 (n_15247, n17719);
  not g32584 (n_15248, n17720);
  and g32585 (n17721, n_15247, n_15248);
  not g32586 (n_15249, n17710);
  not g32587 (n_15250, n17721);
  and g32588 (n17722, n_15249, n_15250);
  and g32589 (n17723, n17710, n17721);
  not g32590 (n_15251, n17722);
  not g32591 (n_15252, n17723);
  and g32592 (n17724, n_15251, n_15252);
  and g32593 (n17725, \b[41] , n4287);
  and g32594 (n17726, \b[39] , n4532);
  and g32595 (n17727, \b[40] , n4282);
  and g32601 (n17730, n4290, n6219);
  not g32604 (n_15257, n17731);
  and g32605 (n17732, \a[35] , n_15257);
  not g32606 (n_15258, n17732);
  and g32607 (n17733, \a[35] , n_15258);
  and g32608 (n17734, n_15257, n_15258);
  not g32609 (n_15259, n17733);
  not g32610 (n_15260, n17734);
  and g32611 (n17735, n_15259, n_15260);
  and g32612 (n17736, n_15070, n_15075);
  and g32613 (n17737, \b[35] , n5777);
  and g32614 (n17738, \b[33] , n6059);
  and g32615 (n17739, \b[34] , n5772);
  and g32621 (n17742, n4696, n5780);
  not g32624 (n_15265, n17743);
  and g32625 (n17744, \a[41] , n_15265);
  not g32626 (n_15266, n17744);
  and g32627 (n17745, \a[41] , n_15266);
  and g32628 (n17746, n_15265, n_15266);
  not g32629 (n_15267, n17745);
  not g32630 (n_15268, n17746);
  and g32631 (n17747, n_15267, n_15268);
  and g32632 (n17748, n_15016, n_15026);
  and g32633 (n17749, \b[26] , n8362);
  and g32634 (n17750, \b[24] , n8715);
  and g32635 (n17751, \b[25] , n8357);
  and g32641 (n17754, n2813, n8365);
  not g32644 (n_15273, n17755);
  and g32645 (n17756, \a[50] , n_15273);
  not g32646 (n_15274, n17756);
  and g32647 (n17757, \a[50] , n_15274);
  and g32648 (n17758, n_15273, n_15274);
  not g32649 (n_15275, n17757);
  not g32650 (n_15276, n17758);
  and g32651 (n17759, n_15275, n_15276);
  and g32652 (n17760, n_15000, n_15010);
  and g32653 (n17761, \b[23] , n9339);
  and g32654 (n17762, \b[21] , n9732);
  and g32655 (n17763, \b[22] , n9334);
  and g32661 (n17766, n2300, n9342);
  not g32664 (n_15281, n17767);
  and g32665 (n17768, \a[53] , n_15281);
  not g32666 (n_15282, n17768);
  and g32667 (n17769, \a[53] , n_15282);
  and g32668 (n17770, n_15281, n_15282);
  not g32669 (n_15283, n17769);
  not g32670 (n_15284, n17770);
  and g32671 (n17771, n_15283, n_15284);
  and g32672 (n17772, n_14984, n_14994);
  and g32673 (n17773, n_14954, n_14959);
  and g32674 (n17774, \b[10] , n13903);
  and g32675 (n17775, \b[11] , n_11555);
  not g32676 (n_15285, n17774);
  not g32677 (n_15286, n17775);
  and g32678 (n17776, n_15285, n_15286);
  not g32679 (n_15287, n17776);
  and g32680 (n17777, n17385, n_15287);
  not g32681 (n_15288, n17777);
  and g32682 (n17778, n17385, n_15288);
  and g32683 (n17779, n_15287, n_15288);
  not g32684 (n_15289, n17778);
  not g32685 (n_15290, n17779);
  and g32686 (n17780, n_15289, n_15290);
  not g32687 (n_15291, n17773);
  not g32688 (n_15292, n17780);
  and g32689 (n17781, n_15291, n_15292);
  not g32690 (n_15293, n17781);
  and g32691 (n17782, n_15291, n_15293);
  and g32692 (n17783, n_15292, n_15293);
  not g32693 (n_15294, n17782);
  not g32694 (n_15295, n17783);
  and g32695 (n17784, n_15294, n_15295);
  and g32696 (n17785, \b[14] , n12668);
  and g32697 (n17786, \b[12] , n13047);
  and g32698 (n17787, \b[13] , n12663);
  and g32704 (n17790, n1034, n12671);
  not g32707 (n_15300, n17791);
  and g32708 (n17792, \a[62] , n_15300);
  not g32709 (n_15301, n17792);
  and g32710 (n17793, \a[62] , n_15301);
  and g32711 (n17794, n_15300, n_15301);
  not g32712 (n_15302, n17793);
  not g32713 (n_15303, n17794);
  and g32714 (n17795, n_15302, n_15303);
  not g32715 (n_15304, n17784);
  not g32716 (n_15305, n17795);
  and g32717 (n17796, n_15304, n_15305);
  not g32718 (n_15306, n17796);
  and g32719 (n17797, n_15304, n_15306);
  and g32720 (n17798, n_15305, n_15306);
  not g32721 (n_15307, n17797);
  not g32722 (n_15308, n17798);
  and g32723 (n17799, n_15307, n_15308);
  and g32724 (n17800, \b[17] , n11531);
  and g32725 (n17801, \b[15] , n11896);
  and g32726 (n17802, \b[16] , n11526);
  and g32732 (n17805, n1356, n11534);
  not g32735 (n_15313, n17806);
  and g32736 (n17807, \a[59] , n_15313);
  not g32737 (n_15314, n17807);
  and g32738 (n17808, \a[59] , n_15314);
  and g32739 (n17809, n_15313, n_15314);
  not g32740 (n_15315, n17808);
  not g32741 (n_15316, n17809);
  and g32742 (n17810, n_15315, n_15316);
  not g32743 (n_15317, n17799);
  not g32744 (n_15318, n17810);
  and g32745 (n17811, n_15317, n_15318);
  not g32746 (n_15319, n17811);
  and g32747 (n17812, n_15317, n_15319);
  and g32748 (n17813, n_15318, n_15319);
  not g32749 (n_15320, n17812);
  not g32750 (n_15321, n17813);
  and g32751 (n17814, n_15320, n_15321);
  and g32752 (n17815, n_14965, n_14978);
  and g32753 (n17816, n17814, n17815);
  not g32754 (n_15322, n17814);
  not g32755 (n_15323, n17815);
  and g32756 (n17817, n_15322, n_15323);
  not g32757 (n_15324, n17816);
  not g32758 (n_15325, n17817);
  and g32759 (n17818, n_15324, n_15325);
  and g32760 (n17819, \b[20] , n10426);
  and g32761 (n17820, \b[18] , n10796);
  and g32762 (n17821, \b[19] , n10421);
  and g32768 (n17824, n1846, n10429);
  not g32771 (n_15330, n17825);
  and g32772 (n17826, \a[56] , n_15330);
  not g32773 (n_15331, n17826);
  and g32774 (n17827, \a[56] , n_15331);
  and g32775 (n17828, n_15330, n_15331);
  not g32776 (n_15332, n17827);
  not g32777 (n_15333, n17828);
  and g32778 (n17829, n_15332, n_15333);
  not g32779 (n_15334, n17818);
  and g32780 (n17830, n_15334, n17829);
  not g32781 (n_15335, n17829);
  and g32782 (n17831, n17818, n_15335);
  not g32783 (n_15336, n17830);
  not g32784 (n_15337, n17831);
  and g32785 (n17832, n_15336, n_15337);
  not g32786 (n_15338, n17772);
  and g32787 (n17833, n_15338, n17832);
  not g32788 (n_15339, n17833);
  and g32789 (n17834, n_15338, n_15339);
  and g32790 (n17835, n17832, n_15339);
  not g32791 (n_15340, n17834);
  not g32792 (n_15341, n17835);
  and g32793 (n17836, n_15340, n_15341);
  not g32794 (n_15342, n17771);
  not g32795 (n_15343, n17836);
  and g32796 (n17837, n_15342, n_15343);
  and g32797 (n17838, n17771, n_15341);
  and g32798 (n17839, n_15340, n17838);
  not g32799 (n_15344, n17837);
  not g32800 (n_15345, n17839);
  and g32801 (n17840, n_15344, n_15345);
  not g32802 (n_15346, n17760);
  and g32803 (n17841, n_15346, n17840);
  not g32804 (n_15347, n17840);
  and g32805 (n17842, n17760, n_15347);
  not g32806 (n_15348, n17841);
  not g32807 (n_15349, n17842);
  and g32808 (n17843, n_15348, n_15349);
  not g32809 (n_15350, n17759);
  and g32810 (n17844, n_15350, n17843);
  not g32811 (n_15351, n17843);
  and g32812 (n17845, n17759, n_15351);
  not g32813 (n_15352, n17844);
  not g32814 (n_15353, n17845);
  and g32815 (n17846, n_15352, n_15353);
  not g32816 (n_15354, n17748);
  and g32817 (n17847, n_15354, n17846);
  not g32818 (n_15355, n17846);
  and g32819 (n17848, n17748, n_15355);
  not g32820 (n_15356, n17847);
  not g32821 (n_15357, n17848);
  and g32822 (n17849, n_15356, n_15357);
  and g32823 (n17850, \b[29] , n7446);
  and g32824 (n17851, \b[27] , n7787);
  and g32825 (n17852, \b[28] , n7441);
  and g32831 (n17855, n3383, n7449);
  not g32834 (n_15362, n17856);
  and g32835 (n17857, \a[47] , n_15362);
  not g32836 (n_15363, n17857);
  and g32837 (n17858, \a[47] , n_15363);
  and g32838 (n17859, n_15362, n_15363);
  not g32839 (n_15364, n17858);
  not g32840 (n_15365, n17859);
  and g32841 (n17860, n_15364, n_15365);
  not g32842 (n_15366, n17860);
  and g32843 (n17861, n17849, n_15366);
  not g32844 (n_15367, n17861);
  and g32845 (n17862, n17849, n_15367);
  and g32846 (n17863, n_15366, n_15367);
  not g32847 (n_15368, n17862);
  not g32848 (n_15369, n17863);
  and g32849 (n17864, n_15368, n_15369);
  and g32850 (n17865, n_15032, n_15042);
  and g32851 (n17866, n17864, n17865);
  not g32852 (n_15370, n17864);
  not g32853 (n_15371, n17865);
  and g32854 (n17867, n_15370, n_15371);
  not g32855 (n_15372, n17866);
  not g32856 (n_15373, n17867);
  and g32857 (n17868, n_15372, n_15373);
  and g32858 (n17869, \b[32] , n6595);
  and g32859 (n17870, \b[30] , n6902);
  and g32860 (n17871, \b[31] , n6590);
  and g32866 (n17874, n4013, n6598);
  not g32869 (n_15378, n17875);
  and g32870 (n17876, \a[44] , n_15378);
  not g32871 (n_15379, n17876);
  and g32872 (n17877, \a[44] , n_15379);
  and g32873 (n17878, n_15378, n_15379);
  not g32874 (n_15380, n17877);
  not g32875 (n_15381, n17878);
  and g32876 (n17879, n_15380, n_15381);
  not g32877 (n_15382, n17868);
  and g32878 (n17880, n_15382, n17879);
  not g32879 (n_15383, n17879);
  and g32880 (n17881, n17868, n_15383);
  not g32881 (n_15384, n17880);
  not g32882 (n_15385, n17881);
  and g32883 (n17882, n_15384, n_15385);
  and g32884 (n17883, n_15048, n_15060);
  not g32885 (n_15386, n17883);
  and g32886 (n17884, n17882, n_15386);
  not g32887 (n_15387, n17882);
  and g32888 (n17885, n_15387, n17883);
  not g32889 (n_15388, n17884);
  not g32890 (n_15389, n17885);
  and g32891 (n17886, n_15388, n_15389);
  not g32892 (n_15390, n17747);
  and g32893 (n17887, n_15390, n17886);
  not g32894 (n_15391, n17887);
  and g32895 (n17888, n17886, n_15391);
  and g32896 (n17889, n_15390, n_15391);
  not g32897 (n_15392, n17888);
  not g32898 (n_15393, n17889);
  and g32899 (n17890, n_15392, n_15393);
  and g32900 (n17891, n_15063, n_15067);
  and g32901 (n17892, n17890, n17891);
  not g32902 (n_15394, n17890);
  not g32903 (n_15395, n17891);
  and g32904 (n17893, n_15394, n_15395);
  not g32905 (n_15396, n17892);
  not g32906 (n_15397, n17893);
  and g32907 (n17894, n_15396, n_15397);
  and g32908 (n17895, \b[38] , n5035);
  and g32909 (n17896, \b[36] , n5277);
  and g32910 (n17897, \b[37] , n5030);
  and g32916 (n17900, n5038, n5205);
  not g32919 (n_15402, n17901);
  and g32920 (n17902, \a[38] , n_15402);
  not g32921 (n_15403, n17902);
  and g32922 (n17903, \a[38] , n_15403);
  and g32923 (n17904, n_15402, n_15403);
  not g32924 (n_15404, n17903);
  not g32925 (n_15405, n17904);
  and g32926 (n17905, n_15404, n_15405);
  not g32927 (n_15406, n17894);
  and g32928 (n17906, n_15406, n17905);
  not g32929 (n_15407, n17905);
  and g32930 (n17907, n17894, n_15407);
  not g32931 (n_15408, n17906);
  not g32932 (n_15409, n17907);
  and g32933 (n17908, n_15408, n_15409);
  not g32934 (n_15410, n17736);
  and g32935 (n17909, n_15410, n17908);
  not g32936 (n_15411, n17908);
  and g32937 (n17910, n17736, n_15411);
  not g32938 (n_15412, n17909);
  not g32939 (n_15413, n17910);
  and g32940 (n17911, n_15412, n_15413);
  not g32941 (n_15414, n17735);
  and g32942 (n17912, n_15414, n17911);
  not g32943 (n_15415, n17912);
  and g32944 (n17913, n_15414, n_15415);
  and g32945 (n17914, n17911, n_15415);
  not g32946 (n_15416, n17913);
  not g32947 (n_15417, n17914);
  and g32948 (n17915, n_15416, n_15417);
  not g32949 (n_15418, n17915);
  and g32950 (n17916, n17724, n_15418);
  not g32951 (n_15419, n17916);
  and g32952 (n17917, n17724, n_15419);
  and g32953 (n17918, n_15418, n_15419);
  not g32954 (n_15420, n17917);
  not g32955 (n_15421, n17918);
  and g32956 (n17919, n_15420, n_15421);
  not g32957 (n_15422, n17919);
  and g32958 (n17920, n17709, n_15422);
  not g32959 (n_15423, n17709);
  and g32960 (n17921, n_15423, n17919);
  not g32961 (n_15424, n17921);
  and g32962 (n17922, n17694, n_15424);
  not g32963 (n_15425, n17920);
  and g32964 (n17923, n_15425, n17922);
  not g32965 (n_15426, n17923);
  and g32966 (n17924, n17694, n_15426);
  and g32967 (n17925, n_15424, n_15426);
  and g32968 (n17926, n_15425, n17925);
  not g32969 (n_15427, n17924);
  not g32970 (n_15428, n17926);
  and g32971 (n17927, n_15427, n_15428);
  and g32972 (n17928, n_14902, n_15110);
  and g32973 (n17929, \b[53] , n2048);
  and g32974 (n17930, \b[51] , n2198);
  and g32975 (n17931, \b[52] , n2043);
  not g32976 (n_15429, n17930);
  not g32977 (n_15430, n17931);
  and g32978 (n17932, n_15429, n_15430);
  not g32979 (n_15431, n17929);
  and g32980 (n17933, n_15431, n17932);
  not g32981 (n_15432, n2051);
  and g32982 (n17934, n_15432, n17933);
  and g32983 (n17935, n_13261, n17933);
  not g32984 (n_15433, n17934);
  not g32985 (n_15434, n17935);
  and g32986 (n17936, n_15433, n_15434);
  not g32987 (n_15435, n17936);
  and g32988 (n17937, \a[23] , n_15435);
  and g32989 (n17938, n_1590, n17936);
  not g32990 (n_15436, n17937);
  not g32991 (n_15437, n17938);
  and g32992 (n17939, n_15436, n_15437);
  not g32993 (n_15438, n17928);
  not g32994 (n_15439, n17939);
  and g32995 (n17940, n_15438, n_15439);
  not g32996 (n_15440, n17940);
  and g32997 (n17941, n_15438, n_15440);
  and g32998 (n17942, n_15439, n_15440);
  not g32999 (n_15441, n17941);
  not g33000 (n_15442, n17942);
  and g33001 (n17943, n_15441, n_15442);
  not g33002 (n_15443, n17927);
  not g33003 (n_15444, n17943);
  and g33004 (n17944, n_15443, n_15444);
  not g33005 (n_15445, n17944);
  and g33006 (n17945, n_15443, n_15445);
  and g33007 (n17946, n_15444, n_15445);
  not g33008 (n_15446, n17945);
  not g33009 (n_15447, n17946);
  and g33010 (n17947, n_15446, n_15447);
  not g33011 (n_15448, n17679);
  not g33012 (n_15449, n17947);
  and g33013 (n17948, n_15448, n_15449);
  not g33014 (n_15450, n17948);
  and g33015 (n17949, n_15448, n_15450);
  and g33016 (n17950, n_15449, n_15450);
  not g33017 (n_15451, n17949);
  not g33018 (n_15452, n17950);
  and g33019 (n17951, n_15451, n_15452);
  not g33020 (n_15453, n17951);
  and g33021 (n17952, n17663, n_15453);
  not g33022 (n_15454, n17663);
  and g33023 (n17953, n_15454, n17951);
  not g33024 (n_15455, n17953);
  and g33025 (n17954, n17648, n_15455);
  not g33026 (n_15456, n17952);
  and g33027 (n17955, n_15456, n17954);
  not g33028 (n_15457, n17955);
  and g33029 (n17956, n17648, n_15457);
  and g33030 (n17957, n_15455, n_15457);
  and g33031 (n17958, n_15456, n17957);
  not g33032 (n_15458, n17956);
  not g33033 (n_15459, n17958);
  and g33034 (n17959, n_15458, n_15459);
  not g33035 (n_15460, n17633);
  and g33036 (n17960, n_15460, n17959);
  not g33037 (n_15461, n17959);
  and g33038 (n17961, n17633, n_15461);
  not g33039 (n_15462, n17960);
  not g33040 (n_15463, n17961);
  and g33041 (n17962, n_15462, n_15463);
  not g33042 (n_15464, n17621);
  not g33043 (n_15465, n17962);
  and g33044 (n17963, n_15464, n_15465);
  not g33045 (n_15466, n17963);
  and g33046 (n17964, n_15464, n_15466);
  and g33047 (n17965, n_15465, n_15466);
  not g33048 (n_15467, n17964);
  not g33049 (n_15468, n17965);
  and g33050 (n17966, n_15467, n_15468);
  not g33051 (n_15469, n17620);
  not g33052 (n_15470, n17966);
  and g33053 (n17967, n_15469, n_15470);
  and g33054 (n17968, n17620, n_15468);
  and g33055 (n17969, n_15467, n17968);
  not g33056 (n_15471, n17967);
  not g33057 (n_15472, n17969);
  and g33058 (\f[74] , n_15471, n_15472);
  and g33059 (n17971, n_15466, n_15471);
  and g33060 (n17972, n_15460, n_15461);
  not g33061 (n_15473, n17972);
  and g33062 (n17973, n_15176, n_15473);
  and g33063 (n17974, n_15189, n_15457);
  and g33064 (n17975, \b[63] , n951);
  and g33065 (n17976, \b[61] , n1056);
  and g33066 (n17977, \b[62] , n946);
  and g33072 (n17980, n954, n13771);
  not g33075 (n_15478, n17981);
  and g33076 (n17982, \a[14] , n_15478);
  not g33077 (n_15479, n17982);
  and g33078 (n17983, \a[14] , n_15479);
  and g33079 (n17984, n_15478, n_15479);
  not g33080 (n_15480, n17983);
  not g33081 (n_15481, n17984);
  and g33082 (n17985, n_15480, n_15481);
  not g33083 (n_15482, n17974);
  not g33084 (n_15483, n17985);
  and g33085 (n17986, n_15482, n_15483);
  not g33086 (n_15484, n17986);
  and g33087 (n17987, n_15482, n_15484);
  and g33088 (n17988, n_15483, n_15484);
  not g33089 (n_15485, n17987);
  not g33090 (n_15486, n17988);
  and g33091 (n17989, n_15485, n_15486);
  and g33092 (n17990, n_15202, n_15456);
  and g33093 (n17991, \b[60] , n1302);
  and g33094 (n17992, \b[58] , n1391);
  and g33095 (n17993, \b[59] , n1297);
  and g33101 (n17996, n1305, n12211);
  not g33104 (n_15491, n17997);
  and g33105 (n17998, \a[17] , n_15491);
  not g33106 (n_15492, n17998);
  and g33107 (n17999, \a[17] , n_15492);
  and g33108 (n18000, n_15491, n_15492);
  not g33109 (n_15493, n17999);
  not g33110 (n_15494, n18000);
  and g33111 (n18001, n_15493, n_15494);
  not g33112 (n_15495, n17990);
  and g33113 (n18002, n_15495, n18001);
  not g33114 (n_15496, n18001);
  and g33115 (n18003, n17990, n_15496);
  not g33116 (n_15497, n18002);
  not g33117 (n_15498, n18003);
  and g33118 (n18004, n_15497, n_15498);
  and g33119 (n18005, \b[57] , n1627);
  and g33120 (n18006, \b[55] , n1763);
  and g33121 (n18007, \b[56] , n1622);
  and g33127 (n18010, n1630, n11410);
  not g33130 (n_15503, n18011);
  and g33131 (n18012, \a[20] , n_15503);
  not g33132 (n_15504, n18012);
  and g33133 (n18013, \a[20] , n_15504);
  and g33134 (n18014, n_15503, n_15504);
  not g33135 (n_15505, n18013);
  not g33136 (n_15506, n18014);
  and g33137 (n18015, n_15505, n_15506);
  and g33138 (n18016, n_15213, n_15450);
  and g33139 (n18017, n18015, n18016);
  not g33140 (n_15507, n18015);
  not g33141 (n_15508, n18016);
  and g33142 (n18018, n_15507, n_15508);
  not g33143 (n_15509, n18017);
  not g33144 (n_15510, n18018);
  and g33145 (n18019, n_15509, n_15510);
  and g33146 (n18020, n_15440, n_15445);
  and g33147 (n18021, \b[54] , n2048);
  and g33148 (n18022, \b[52] , n2198);
  and g33149 (n18023, \b[53] , n2043);
  and g33155 (n18026, n2051, n9998);
  not g33158 (n_15515, n18027);
  and g33159 (n18028, \a[23] , n_15515);
  not g33160 (n_15516, n18028);
  and g33161 (n18029, \a[23] , n_15516);
  and g33162 (n18030, n_15515, n_15516);
  not g33163 (n_15517, n18029);
  not g33164 (n_15518, n18030);
  and g33165 (n18031, n_15517, n_15518);
  not g33166 (n_15519, n18020);
  not g33167 (n_15520, n18031);
  and g33168 (n18032, n_15519, n_15520);
  not g33169 (n_15521, n18032);
  and g33170 (n18033, n_15519, n_15521);
  and g33171 (n18034, n_15520, n_15521);
  not g33172 (n_15522, n18033);
  not g33173 (n_15523, n18034);
  and g33174 (n18035, n_15522, n_15523);
  and g33175 (n18036, \b[51] , n2539);
  and g33176 (n18037, \b[49] , n2685);
  and g33177 (n18038, \b[50] , n2534);
  and g33183 (n18041, n2542, n8976);
  not g33186 (n_15528, n18042);
  and g33187 (n18043, \a[26] , n_15528);
  not g33188 (n_15529, n18043);
  and g33189 (n18044, \a[26] , n_15529);
  and g33190 (n18045, n_15528, n_15529);
  not g33191 (n_15530, n18044);
  not g33192 (n_15531, n18045);
  and g33193 (n18046, n_15530, n_15531);
  and g33194 (n18047, n_15227, n_15426);
  and g33195 (n18048, n18046, n18047);
  not g33196 (n_15532, n18046);
  not g33197 (n_15533, n18047);
  and g33198 (n18049, n_15532, n_15533);
  not g33199 (n_15534, n18048);
  not g33200 (n_15535, n18049);
  and g33201 (n18050, n_15534, n_15535);
  and g33202 (n18051, n_15240, n_15425);
  and g33203 (n18052, \b[48] , n3050);
  and g33204 (n18053, \b[46] , n3243);
  and g33205 (n18054, \b[47] , n3045);
  and g33211 (n18057, n3053, n8009);
  not g33214 (n_15540, n18058);
  and g33215 (n18059, \a[29] , n_15540);
  not g33216 (n_15541, n18059);
  and g33217 (n18060, \a[29] , n_15541);
  and g33218 (n18061, n_15540, n_15541);
  not g33219 (n_15542, n18060);
  not g33220 (n_15543, n18061);
  and g33221 (n18062, n_15542, n_15543);
  not g33222 (n_15544, n18051);
  and g33223 (n18063, n_15544, n18062);
  not g33224 (n_15545, n18062);
  and g33225 (n18064, n18051, n_15545);
  not g33226 (n_15546, n18063);
  not g33227 (n_15547, n18064);
  and g33228 (n18065, n_15546, n_15547);
  and g33229 (n18066, n_15412, n_15415);
  and g33230 (n18067, n_15397, n_15409);
  and g33231 (n18068, n_15388, n_15391);
  and g33232 (n18069, n_15373, n_15385);
  and g33233 (n18070, n_15356, n_15367);
  and g33234 (n18071, n_15339, n_15344);
  and g33235 (n18072, \b[24] , n9339);
  and g33236 (n18073, \b[22] , n9732);
  and g33237 (n18074, \b[23] , n9334);
  and g33243 (n18077, n2458, n9342);
  not g33246 (n_15552, n18078);
  and g33247 (n18079, \a[53] , n_15552);
  not g33248 (n_15553, n18079);
  and g33249 (n18080, \a[53] , n_15553);
  and g33250 (n18081, n_15552, n_15553);
  not g33251 (n_15554, n18080);
  not g33252 (n_15555, n18081);
  and g33253 (n18082, n_15554, n_15555);
  and g33254 (n18083, n_15288, n_15293);
  and g33255 (n18084, \b[15] , n12668);
  and g33256 (n18085, \b[13] , n13047);
  and g33257 (n18086, \b[14] , n12663);
  and g33263 (n18089, n1131, n12671);
  not g33266 (n_15560, n18090);
  and g33267 (n18091, \a[62] , n_15560);
  not g33268 (n_15561, n18091);
  and g33269 (n18092, \a[62] , n_15561);
  and g33270 (n18093, n_15560, n_15561);
  not g33271 (n_15562, n18092);
  not g33272 (n_15563, n18093);
  and g33273 (n18094, n_15562, n_15563);
  and g33274 (n18095, \b[11] , n13903);
  and g33275 (n18096, \b[12] , n_11555);
  not g33276 (n_15564, n18095);
  not g33277 (n_15565, n18096);
  and g33278 (n18097, n_15564, n_15565);
  not g33279 (n_15566, n17385);
  and g33280 (n18098, \a[11] , n_15566);
  and g33281 (n18099, n_400, n17385);
  not g33282 (n_15567, n18098);
  not g33283 (n_15568, n18099);
  and g33284 (n18100, n_15567, n_15568);
  not g33285 (n_15569, n18097);
  not g33286 (n_15570, n18100);
  and g33287 (n18101, n_15569, n_15570);
  and g33288 (n18102, n18097, n18100);
  not g33289 (n_15571, n18101);
  not g33290 (n_15572, n18102);
  and g33291 (n18103, n_15571, n_15572);
  not g33292 (n_15573, n18094);
  and g33293 (n18104, n_15573, n18103);
  not g33294 (n_15574, n18104);
  and g33295 (n18105, n_15573, n_15574);
  and g33296 (n18106, n18103, n_15574);
  not g33297 (n_15575, n18105);
  not g33298 (n_15576, n18106);
  and g33299 (n18107, n_15575, n_15576);
  not g33300 (n_15577, n18083);
  not g33301 (n_15578, n18107);
  and g33302 (n18108, n_15577, n_15578);
  not g33303 (n_15579, n18108);
  and g33304 (n18109, n_15577, n_15579);
  and g33305 (n18110, n_15578, n_15579);
  not g33306 (n_15580, n18109);
  not g33307 (n_15581, n18110);
  and g33308 (n18111, n_15580, n_15581);
  and g33309 (n18112, \b[18] , n11531);
  and g33310 (n18113, \b[16] , n11896);
  and g33311 (n18114, \b[17] , n11526);
  and g33317 (n18117, n1566, n11534);
  not g33320 (n_15586, n18118);
  and g33321 (n18119, \a[59] , n_15586);
  not g33322 (n_15587, n18119);
  and g33323 (n18120, \a[59] , n_15587);
  and g33324 (n18121, n_15586, n_15587);
  not g33325 (n_15588, n18120);
  not g33326 (n_15589, n18121);
  and g33327 (n18122, n_15588, n_15589);
  not g33328 (n_15590, n18111);
  not g33329 (n_15591, n18122);
  and g33330 (n18123, n_15590, n_15591);
  not g33331 (n_15592, n18123);
  and g33332 (n18124, n_15590, n_15592);
  and g33333 (n18125, n_15591, n_15592);
  not g33334 (n_15593, n18124);
  not g33335 (n_15594, n18125);
  and g33336 (n18126, n_15593, n_15594);
  and g33337 (n18127, n_15306, n_15319);
  and g33338 (n18128, n18126, n18127);
  not g33339 (n_15595, n18126);
  not g33340 (n_15596, n18127);
  and g33341 (n18129, n_15595, n_15596);
  not g33342 (n_15597, n18128);
  not g33343 (n_15598, n18129);
  and g33344 (n18130, n_15597, n_15598);
  and g33345 (n18131, \b[21] , n10426);
  and g33346 (n18132, \b[19] , n10796);
  and g33347 (n18133, \b[20] , n10421);
  and g33353 (n18136, n1984, n10429);
  not g33356 (n_15603, n18137);
  and g33357 (n18138, \a[56] , n_15603);
  not g33358 (n_15604, n18138);
  and g33359 (n18139, \a[56] , n_15604);
  and g33360 (n18140, n_15603, n_15604);
  not g33361 (n_15605, n18139);
  not g33362 (n_15606, n18140);
  and g33363 (n18141, n_15605, n_15606);
  not g33364 (n_15607, n18141);
  and g33365 (n18142, n18130, n_15607);
  not g33366 (n_15608, n18142);
  and g33367 (n18143, n18130, n_15608);
  and g33368 (n18144, n_15607, n_15608);
  not g33369 (n_15609, n18143);
  not g33370 (n_15610, n18144);
  and g33371 (n18145, n_15609, n_15610);
  and g33372 (n18146, n_15325, n_15337);
  not g33373 (n_15611, n18145);
  not g33374 (n_15612, n18146);
  and g33375 (n18147, n_15611, n_15612);
  and g33376 (n18148, n18145, n18146);
  not g33377 (n_15613, n18147);
  not g33378 (n_15614, n18148);
  and g33379 (n18149, n_15613, n_15614);
  not g33380 (n_15615, n18082);
  and g33381 (n18150, n_15615, n18149);
  not g33382 (n_15616, n18150);
  and g33383 (n18151, n_15615, n_15616);
  and g33384 (n18152, n18149, n_15616);
  not g33385 (n_15617, n18151);
  not g33386 (n_15618, n18152);
  and g33387 (n18153, n_15617, n_15618);
  not g33388 (n_15619, n18071);
  not g33389 (n_15620, n18153);
  and g33390 (n18154, n_15619, n_15620);
  not g33391 (n_15621, n18154);
  and g33392 (n18155, n_15619, n_15621);
  and g33393 (n18156, n_15620, n_15621);
  not g33394 (n_15622, n18155);
  not g33395 (n_15623, n18156);
  and g33396 (n18157, n_15622, n_15623);
  and g33397 (n18158, \b[27] , n8362);
  and g33398 (n18159, \b[25] , n8715);
  and g33399 (n18160, \b[26] , n8357);
  and g33405 (n18163, n2990, n8365);
  not g33408 (n_15628, n18164);
  and g33409 (n18165, \a[50] , n_15628);
  not g33410 (n_15629, n18165);
  and g33411 (n18166, \a[50] , n_15629);
  and g33412 (n18167, n_15628, n_15629);
  not g33413 (n_15630, n18166);
  not g33414 (n_15631, n18167);
  and g33415 (n18168, n_15630, n_15631);
  not g33416 (n_15632, n18157);
  not g33417 (n_15633, n18168);
  and g33418 (n18169, n_15632, n_15633);
  not g33419 (n_15634, n18169);
  and g33420 (n18170, n_15632, n_15634);
  and g33421 (n18171, n_15633, n_15634);
  not g33422 (n_15635, n18170);
  not g33423 (n_15636, n18171);
  and g33424 (n18172, n_15635, n_15636);
  and g33425 (n18173, n_15348, n_15352);
  and g33426 (n18174, n18172, n18173);
  not g33427 (n_15637, n18172);
  not g33428 (n_15638, n18173);
  and g33429 (n18175, n_15637, n_15638);
  not g33430 (n_15639, n18174);
  not g33431 (n_15640, n18175);
  and g33432 (n18176, n_15639, n_15640);
  and g33433 (n18177, \b[30] , n7446);
  and g33434 (n18178, \b[28] , n7787);
  and g33435 (n18179, \b[29] , n7441);
  and g33441 (n18182, n3577, n7449);
  not g33444 (n_15645, n18183);
  and g33445 (n18184, \a[47] , n_15645);
  not g33446 (n_15646, n18184);
  and g33447 (n18185, \a[47] , n_15646);
  and g33448 (n18186, n_15645, n_15646);
  not g33449 (n_15647, n18185);
  not g33450 (n_15648, n18186);
  and g33451 (n18187, n_15647, n_15648);
  not g33452 (n_15649, n18187);
  and g33453 (n18188, n18176, n_15649);
  not g33454 (n_15650, n18176);
  and g33455 (n18189, n_15650, n18187);
  not g33456 (n_15651, n18070);
  not g33457 (n_15652, n18189);
  and g33458 (n18190, n_15651, n_15652);
  not g33459 (n_15653, n18188);
  and g33460 (n18191, n_15653, n18190);
  not g33461 (n_15654, n18191);
  and g33462 (n18192, n_15651, n_15654);
  and g33463 (n18193, n_15653, n_15654);
  and g33464 (n18194, n_15652, n18193);
  not g33465 (n_15655, n18192);
  not g33466 (n_15656, n18194);
  and g33467 (n18195, n_15655, n_15656);
  and g33468 (n18196, \b[33] , n6595);
  and g33469 (n18197, \b[31] , n6902);
  and g33470 (n18198, \b[32] , n6590);
  and g33476 (n18201, n4223, n6598);
  not g33479 (n_15661, n18202);
  and g33480 (n18203, \a[44] , n_15661);
  not g33481 (n_15662, n18203);
  and g33482 (n18204, \a[44] , n_15662);
  and g33483 (n18205, n_15661, n_15662);
  not g33484 (n_15663, n18204);
  not g33485 (n_15664, n18205);
  and g33486 (n18206, n_15663, n_15664);
  not g33487 (n_15665, n18195);
  not g33488 (n_15666, n18206);
  and g33489 (n18207, n_15665, n_15666);
  not g33490 (n_15667, n18207);
  and g33491 (n18208, n_15665, n_15667);
  and g33492 (n18209, n_15666, n_15667);
  not g33493 (n_15668, n18208);
  not g33494 (n_15669, n18209);
  and g33495 (n18210, n_15668, n_15669);
  not g33496 (n_15670, n18069);
  and g33497 (n18211, n_15670, n18210);
  not g33498 (n_15671, n18210);
  and g33499 (n18212, n18069, n_15671);
  not g33500 (n_15672, n18211);
  not g33501 (n_15673, n18212);
  and g33502 (n18213, n_15672, n_15673);
  and g33503 (n18214, \b[36] , n5777);
  and g33504 (n18215, \b[34] , n6059);
  and g33505 (n18216, \b[35] , n5772);
  and g33511 (n18219, n4922, n5780);
  not g33514 (n_15678, n18220);
  and g33515 (n18221, \a[41] , n_15678);
  not g33516 (n_15679, n18221);
  and g33517 (n18222, \a[41] , n_15679);
  and g33518 (n18223, n_15678, n_15679);
  not g33519 (n_15680, n18222);
  not g33520 (n_15681, n18223);
  and g33521 (n18224, n_15680, n_15681);
  not g33522 (n_15682, n18213);
  not g33523 (n_15683, n18224);
  and g33524 (n18225, n_15682, n_15683);
  and g33525 (n18226, n18213, n18224);
  not g33526 (n_15684, n18225);
  not g33527 (n_15685, n18226);
  and g33528 (n18227, n_15684, n_15685);
  not g33529 (n_15686, n18227);
  and g33530 (n18228, n18068, n_15686);
  not g33531 (n_15687, n18068);
  and g33532 (n18229, n_15687, n18227);
  not g33533 (n_15688, n18228);
  not g33534 (n_15689, n18229);
  and g33535 (n18230, n_15688, n_15689);
  and g33536 (n18231, \b[39] , n5035);
  and g33537 (n18232, \b[37] , n5277);
  and g33538 (n18233, \b[38] , n5030);
  and g33544 (n18236, n5038, n5451);
  not g33547 (n_15694, n18237);
  and g33548 (n18238, \a[38] , n_15694);
  not g33549 (n_15695, n18238);
  and g33550 (n18239, \a[38] , n_15695);
  and g33551 (n18240, n_15694, n_15695);
  not g33552 (n_15696, n18239);
  not g33553 (n_15697, n18240);
  and g33554 (n18241, n_15696, n_15697);
  not g33555 (n_15698, n18241);
  and g33556 (n18242, n18230, n_15698);
  not g33557 (n_15699, n18242);
  and g33558 (n18243, n18230, n_15699);
  and g33559 (n18244, n_15698, n_15699);
  not g33560 (n_15700, n18243);
  not g33561 (n_15701, n18244);
  and g33562 (n18245, n_15700, n_15701);
  not g33563 (n_15702, n18067);
  and g33564 (n18246, n_15702, n18245);
  not g33565 (n_15703, n18245);
  and g33566 (n18247, n18067, n_15703);
  not g33567 (n_15704, n18246);
  not g33568 (n_15705, n18247);
  and g33569 (n18248, n_15704, n_15705);
  and g33570 (n18249, \b[42] , n4287);
  and g33571 (n18250, \b[40] , n4532);
  and g33572 (n18251, \b[41] , n4282);
  and g33578 (n18254, n4290, n6489);
  not g33581 (n_15710, n18255);
  and g33582 (n18256, \a[35] , n_15710);
  not g33583 (n_15711, n18256);
  and g33584 (n18257, \a[35] , n_15711);
  and g33585 (n18258, n_15710, n_15711);
  not g33586 (n_15712, n18257);
  not g33587 (n_15713, n18258);
  and g33588 (n18259, n_15712, n_15713);
  not g33589 (n_15714, n18248);
  not g33590 (n_15715, n18259);
  and g33591 (n18260, n_15714, n_15715);
  and g33592 (n18261, n18248, n18259);
  not g33593 (n_15716, n18260);
  not g33594 (n_15717, n18261);
  and g33595 (n18262, n_15716, n_15717);
  not g33596 (n_15718, n18262);
  and g33597 (n18263, n18066, n_15718);
  not g33598 (n_15719, n18066);
  and g33599 (n18264, n_15719, n18262);
  not g33600 (n_15720, n18263);
  not g33601 (n_15721, n18264);
  and g33602 (n18265, n_15720, n_15721);
  and g33603 (n18266, n_15251, n_15419);
  and g33604 (n18267, \b[45] , n3638);
  and g33605 (n18268, \b[43] , n3843);
  and g33606 (n18269, \b[44] , n3633);
  and g33612 (n18272, n3641, n7361);
  not g33615 (n_15726, n18273);
  and g33616 (n18274, \a[32] , n_15726);
  not g33617 (n_15727, n18274);
  and g33618 (n18275, \a[32] , n_15727);
  and g33619 (n18276, n_15726, n_15727);
  not g33620 (n_15728, n18275);
  not g33621 (n_15729, n18276);
  and g33622 (n18277, n_15728, n_15729);
  not g33623 (n_15730, n18266);
  not g33624 (n_15731, n18277);
  and g33625 (n18278, n_15730, n_15731);
  not g33626 (n_15732, n18278);
  and g33627 (n18279, n_15730, n_15732);
  and g33628 (n18280, n_15731, n_15732);
  not g33629 (n_15733, n18279);
  not g33630 (n_15734, n18280);
  and g33631 (n18281, n_15733, n_15734);
  not g33632 (n_15735, n18281);
  and g33633 (n18282, n18265, n_15735);
  not g33634 (n_15736, n18265);
  and g33635 (n18283, n_15736, n18281);
  not g33636 (n_15737, n18065);
  not g33637 (n_15738, n18283);
  and g33638 (n18284, n_15737, n_15738);
  not g33639 (n_15739, n18282);
  and g33640 (n18285, n_15739, n18284);
  not g33641 (n_15740, n18285);
  and g33642 (n18286, n_15737, n_15740);
  and g33643 (n18287, n_15738, n_15740);
  and g33644 (n18288, n_15739, n18287);
  not g33645 (n_15741, n18286);
  not g33646 (n_15742, n18288);
  and g33647 (n18289, n_15741, n_15742);
  not g33648 (n_15743, n18289);
  and g33649 (n18290, n18050, n_15743);
  not g33650 (n_15744, n18050);
  and g33651 (n18291, n_15744, n18289);
  not g33652 (n_15745, n18035);
  not g33653 (n_15746, n18291);
  and g33654 (n18292, n_15745, n_15746);
  not g33655 (n_15747, n18290);
  and g33656 (n18293, n_15747, n18292);
  not g33657 (n_15748, n18293);
  and g33658 (n18294, n_15745, n_15748);
  and g33659 (n18295, n_15746, n_15748);
  and g33660 (n18296, n_15747, n18295);
  not g33661 (n_15749, n18294);
  not g33662 (n_15750, n18296);
  and g33663 (n18297, n_15749, n_15750);
  not g33664 (n_15751, n18297);
  and g33665 (n18298, n18019, n_15751);
  not g33666 (n_15752, n18019);
  and g33667 (n18299, n_15752, n18297);
  not g33668 (n_15753, n18004);
  not g33669 (n_15754, n18299);
  and g33670 (n18300, n_15753, n_15754);
  not g33671 (n_15755, n18298);
  and g33672 (n18301, n_15755, n18300);
  not g33673 (n_15756, n18301);
  and g33674 (n18302, n_15753, n_15756);
  and g33675 (n18303, n_15754, n_15756);
  and g33676 (n18304, n_15755, n18303);
  not g33677 (n_15757, n18302);
  not g33678 (n_15758, n18304);
  and g33679 (n18305, n_15757, n_15758);
  not g33680 (n_15759, n17989);
  and g33681 (n18306, n_15759, n18305);
  not g33682 (n_15760, n18305);
  and g33683 (n18307, n17989, n_15760);
  not g33684 (n_15761, n18306);
  not g33685 (n_15762, n18307);
  and g33686 (n18308, n_15761, n_15762);
  not g33687 (n_15763, n17973);
  not g33688 (n_15764, n18308);
  and g33689 (n18309, n_15763, n_15764);
  not g33690 (n_15765, n18309);
  and g33691 (n18310, n_15763, n_15765);
  and g33692 (n18311, n_15764, n_15765);
  not g33693 (n_15766, n18310);
  not g33694 (n_15767, n18311);
  and g33695 (n18312, n_15766, n_15767);
  not g33696 (n_15768, n17971);
  not g33697 (n_15769, n18312);
  and g33698 (n18313, n_15768, n_15769);
  and g33699 (n18314, n17971, n_15767);
  and g33700 (n18315, n_15766, n18314);
  not g33701 (n_15770, n18313);
  not g33702 (n_15771, n18315);
  and g33703 (\f[75] , n_15770, n_15771);
  and g33704 (n18317, n_15765, n_15770);
  and g33705 (n18318, n_15759, n_15760);
  not g33706 (n_15772, n18318);
  and g33707 (n18319, n_15484, n_15772);
  and g33708 (n18320, \b[61] , n1302);
  and g33709 (n18321, \b[59] , n1391);
  and g33710 (n18322, \b[60] , n1297);
  and g33716 (n18325, n1305, n12969);
  not g33719 (n_15777, n18326);
  and g33720 (n18327, \a[17] , n_15777);
  not g33721 (n_15778, n18327);
  and g33722 (n18328, \a[17] , n_15778);
  and g33723 (n18329, n_15777, n_15778);
  not g33724 (n_15779, n18328);
  not g33725 (n_15780, n18329);
  and g33726 (n18330, n_15779, n_15780);
  and g33727 (n18331, n_15510, n_15755);
  not g33728 (n_15781, n18330);
  not g33729 (n_15782, n18331);
  and g33730 (n18332, n_15781, n_15782);
  not g33731 (n_15783, n18332);
  and g33732 (n18333, n_15781, n_15783);
  and g33733 (n18334, n_15782, n_15783);
  not g33734 (n_15784, n18333);
  not g33735 (n_15785, n18334);
  and g33736 (n18335, n_15784, n_15785);
  and g33737 (n18336, \b[55] , n2048);
  and g33738 (n18337, \b[53] , n2198);
  and g33739 (n18338, \b[54] , n2043);
  and g33745 (n18341, n2051, n10684);
  not g33748 (n_15790, n18342);
  and g33749 (n18343, \a[23] , n_15790);
  not g33750 (n_15791, n18343);
  and g33751 (n18344, \a[23] , n_15791);
  and g33752 (n18345, n_15790, n_15791);
  not g33753 (n_15792, n18344);
  not g33754 (n_15793, n18345);
  and g33755 (n18346, n_15792, n_15793);
  and g33756 (n18347, n_15535, n_15747);
  not g33757 (n_15794, n18346);
  not g33758 (n_15795, n18347);
  and g33759 (n18348, n_15794, n_15795);
  not g33760 (n_15796, n18348);
  and g33761 (n18349, n_15794, n_15796);
  and g33762 (n18350, n_15795, n_15796);
  not g33763 (n_15797, n18349);
  not g33764 (n_15798, n18350);
  and g33765 (n18351, n_15797, n_15798);
  and g33766 (n18352, \b[49] , n3050);
  and g33767 (n18353, \b[47] , n3243);
  and g33768 (n18354, \b[48] , n3045);
  and g33774 (n18357, n3053, n8625);
  not g33777 (n_15803, n18358);
  and g33778 (n18359, \a[29] , n_15803);
  not g33779 (n_15804, n18359);
  and g33780 (n18360, \a[29] , n_15804);
  and g33781 (n18361, n_15803, n_15804);
  not g33782 (n_15805, n18360);
  not g33783 (n_15806, n18361);
  and g33784 (n18362, n_15805, n_15806);
  and g33785 (n18363, n_15732, n_15739);
  not g33786 (n_15807, n18362);
  not g33787 (n_15808, n18363);
  and g33788 (n18364, n_15807, n_15808);
  not g33789 (n_15809, n18364);
  and g33790 (n18365, n_15807, n_15809);
  and g33791 (n18366, n_15808, n_15809);
  not g33792 (n_15810, n18365);
  not g33793 (n_15811, n18366);
  and g33794 (n18367, n_15810, n_15811);
  and g33795 (n18368, \b[43] , n4287);
  and g33796 (n18369, \b[41] , n4532);
  and g33797 (n18370, \b[42] , n4282);
  and g33803 (n18373, n4290, n6515);
  not g33806 (n_15816, n18374);
  and g33807 (n18375, \a[35] , n_15816);
  not g33808 (n_15817, n18375);
  and g33809 (n18376, \a[35] , n_15817);
  and g33810 (n18377, n_15816, n_15817);
  not g33811 (n_15818, n18376);
  not g33812 (n_15819, n18377);
  and g33813 (n18378, n_15818, n_15819);
  and g33814 (n18379, n_15702, n_15703);
  not g33815 (n_15820, n18379);
  and g33816 (n18380, n_15699, n_15820);
  and g33817 (n18381, \b[40] , n5035);
  and g33818 (n18382, \b[38] , n5277);
  and g33819 (n18383, \b[39] , n5030);
  and g33825 (n18386, n5038, n5955);
  not g33828 (n_15825, n18387);
  and g33829 (n18388, \a[38] , n_15825);
  not g33830 (n_15826, n18388);
  and g33831 (n18389, \a[38] , n_15826);
  and g33832 (n18390, n_15825, n_15826);
  not g33833 (n_15827, n18389);
  not g33834 (n_15828, n18390);
  and g33835 (n18391, n_15827, n_15828);
  and g33836 (n18392, n_15684, n_15689);
  and g33837 (n18393, \b[37] , n5777);
  and g33838 (n18394, \b[35] , n6059);
  and g33839 (n18395, \b[36] , n5772);
  and g33845 (n18398, n5181, n5780);
  not g33848 (n_15833, n18399);
  and g33849 (n18400, \a[41] , n_15833);
  not g33850 (n_15834, n18400);
  and g33851 (n18401, \a[41] , n_15834);
  and g33852 (n18402, n_15833, n_15834);
  not g33853 (n_15835, n18401);
  not g33854 (n_15836, n18402);
  and g33855 (n18403, n_15835, n_15836);
  and g33856 (n18404, n_15670, n_15671);
  not g33857 (n_15837, n18404);
  and g33858 (n18405, n_15667, n_15837);
  and g33859 (n18406, \b[34] , n6595);
  and g33860 (n18407, \b[32] , n6902);
  and g33861 (n18408, \b[33] , n6590);
  and g33867 (n18411, n4466, n6598);
  not g33870 (n_15842, n18412);
  and g33871 (n18413, \a[44] , n_15842);
  not g33872 (n_15843, n18413);
  and g33873 (n18414, \a[44] , n_15843);
  and g33874 (n18415, n_15842, n_15843);
  not g33875 (n_15844, n18414);
  not g33876 (n_15845, n18415);
  and g33877 (n18416, n_15844, n_15845);
  and g33878 (n18417, \b[31] , n7446);
  and g33879 (n18418, \b[29] , n7787);
  and g33880 (n18419, \b[30] , n7441);
  and g33886 (n18422, n3796, n7449);
  not g33889 (n_15850, n18423);
  and g33890 (n18424, \a[47] , n_15850);
  not g33891 (n_15851, n18424);
  and g33892 (n18425, \a[47] , n_15851);
  and g33893 (n18426, n_15850, n_15851);
  not g33894 (n_15852, n18425);
  not g33895 (n_15853, n18426);
  and g33896 (n18427, n_15852, n_15853);
  and g33897 (n18428, n_15634, n_15640);
  and g33898 (n18429, \b[12] , n13903);
  and g33899 (n18430, \b[13] , n_11555);
  not g33900 (n_15854, n18429);
  not g33901 (n_15855, n18430);
  and g33902 (n18431, n_15854, n_15855);
  and g33903 (n18432, n_400, n_15566);
  not g33904 (n_15856, n18432);
  and g33905 (n18433, n_15571, n_15856);
  not g33906 (n_15857, n18433);
  and g33907 (n18434, n18431, n_15857);
  not g33908 (n_15858, n18434);
  and g33909 (n18435, n18431, n_15858);
  and g33910 (n18436, n_15857, n_15858);
  not g33911 (n_15859, n18435);
  not g33912 (n_15860, n18436);
  and g33913 (n18437, n_15859, n_15860);
  and g33914 (n18438, \b[16] , n12668);
  and g33915 (n18439, \b[14] , n13047);
  and g33916 (n18440, \b[15] , n12663);
  and g33922 (n18443, n1237, n12671);
  not g33925 (n_15865, n18444);
  and g33926 (n18445, \a[62] , n_15865);
  not g33927 (n_15866, n18445);
  and g33928 (n18446, \a[62] , n_15866);
  and g33929 (n18447, n_15865, n_15866);
  not g33930 (n_15867, n18446);
  not g33931 (n_15868, n18447);
  and g33932 (n18448, n_15867, n_15868);
  not g33933 (n_15869, n18437);
  and g33934 (n18449, n_15869, n18448);
  not g33935 (n_15870, n18448);
  and g33936 (n18450, n18437, n_15870);
  not g33937 (n_15871, n18449);
  not g33938 (n_15872, n18450);
  and g33939 (n18451, n_15871, n_15872);
  and g33940 (n18452, n_15574, n_15579);
  and g33941 (n18453, n18451, n18452);
  not g33942 (n_15873, n18451);
  not g33943 (n_15874, n18452);
  and g33944 (n18454, n_15873, n_15874);
  not g33945 (n_15875, n18453);
  not g33946 (n_15876, n18454);
  and g33947 (n18455, n_15875, n_15876);
  and g33948 (n18456, \b[19] , n11531);
  and g33949 (n18457, \b[17] , n11896);
  and g33950 (n18458, \b[18] , n11526);
  and g33956 (n18461, n1708, n11534);
  not g33959 (n_15881, n18462);
  and g33960 (n18463, \a[59] , n_15881);
  not g33961 (n_15882, n18463);
  and g33962 (n18464, \a[59] , n_15882);
  and g33963 (n18465, n_15881, n_15882);
  not g33964 (n_15883, n18464);
  not g33965 (n_15884, n18465);
  and g33966 (n18466, n_15883, n_15884);
  not g33967 (n_15885, n18466);
  and g33968 (n18467, n18455, n_15885);
  not g33969 (n_15886, n18467);
  and g33970 (n18468, n18455, n_15886);
  and g33971 (n18469, n_15885, n_15886);
  not g33972 (n_15887, n18468);
  not g33973 (n_15888, n18469);
  and g33974 (n18470, n_15887, n_15888);
  and g33975 (n18471, n_15592, n_15598);
  and g33976 (n18472, n18470, n18471);
  not g33977 (n_15889, n18470);
  not g33978 (n_15890, n18471);
  and g33979 (n18473, n_15889, n_15890);
  not g33980 (n_15891, n18472);
  not g33981 (n_15892, n18473);
  and g33982 (n18474, n_15891, n_15892);
  and g33983 (n18475, \b[22] , n10426);
  and g33984 (n18476, \b[20] , n10796);
  and g33985 (n18477, \b[21] , n10421);
  and g33991 (n18480, n2145, n10429);
  not g33994 (n_15897, n18481);
  and g33995 (n18482, \a[56] , n_15897);
  not g33996 (n_15898, n18482);
  and g33997 (n18483, \a[56] , n_15898);
  and g33998 (n18484, n_15897, n_15898);
  not g33999 (n_15899, n18483);
  not g34000 (n_15900, n18484);
  and g34001 (n18485, n_15899, n_15900);
  not g34002 (n_15901, n18485);
  and g34003 (n18486, n18474, n_15901);
  not g34004 (n_15902, n18486);
  and g34005 (n18487, n18474, n_15902);
  and g34006 (n18488, n_15901, n_15902);
  not g34007 (n_15903, n18487);
  not g34008 (n_15904, n18488);
  and g34009 (n18489, n_15903, n_15904);
  and g34010 (n18490, n_15608, n_15613);
  and g34011 (n18491, n18489, n18490);
  not g34012 (n_15905, n18489);
  not g34013 (n_15906, n18490);
  and g34014 (n18492, n_15905, n_15906);
  not g34015 (n_15907, n18491);
  not g34016 (n_15908, n18492);
  and g34017 (n18493, n_15907, n_15908);
  and g34018 (n18494, \b[25] , n9339);
  and g34019 (n18495, \b[23] , n9732);
  and g34020 (n18496, \b[24] , n9334);
  and g34026 (n18499, n2485, n9342);
  not g34029 (n_15913, n18500);
  and g34030 (n18501, \a[53] , n_15913);
  not g34031 (n_15914, n18501);
  and g34032 (n18502, \a[53] , n_15914);
  and g34033 (n18503, n_15913, n_15914);
  not g34034 (n_15915, n18502);
  not g34035 (n_15916, n18503);
  and g34036 (n18504, n_15915, n_15916);
  not g34037 (n_15917, n18504);
  and g34038 (n18505, n18493, n_15917);
  not g34039 (n_15918, n18505);
  and g34040 (n18506, n18493, n_15918);
  and g34041 (n18507, n_15917, n_15918);
  not g34042 (n_15919, n18506);
  not g34043 (n_15920, n18507);
  and g34044 (n18508, n_15919, n_15920);
  and g34045 (n18509, n_15616, n_15621);
  and g34046 (n18510, n18508, n18509);
  not g34047 (n_15921, n18508);
  not g34048 (n_15922, n18509);
  and g34049 (n18511, n_15921, n_15922);
  not g34050 (n_15923, n18510);
  not g34051 (n_15924, n18511);
  and g34052 (n18512, n_15923, n_15924);
  and g34053 (n18513, \b[28] , n8362);
  and g34054 (n18514, \b[26] , n8715);
  and g34055 (n18515, \b[27] , n8357);
  and g34061 (n18518, n3189, n8365);
  not g34064 (n_15929, n18519);
  and g34065 (n18520, \a[50] , n_15929);
  not g34066 (n_15930, n18520);
  and g34067 (n18521, \a[50] , n_15930);
  and g34068 (n18522, n_15929, n_15930);
  not g34069 (n_15931, n18521);
  not g34070 (n_15932, n18522);
  and g34071 (n18523, n_15931, n_15932);
  not g34072 (n_15933, n18512);
  and g34073 (n18524, n_15933, n18523);
  not g34074 (n_15934, n18523);
  and g34075 (n18525, n18512, n_15934);
  not g34076 (n_15935, n18524);
  not g34077 (n_15936, n18525);
  and g34078 (n18526, n_15935, n_15936);
  not g34079 (n_15937, n18428);
  and g34080 (n18527, n_15937, n18526);
  not g34081 (n_15938, n18527);
  and g34082 (n18528, n_15937, n_15938);
  and g34083 (n18529, n18526, n_15938);
  not g34084 (n_15939, n18528);
  not g34085 (n_15940, n18529);
  and g34086 (n18530, n_15939, n_15940);
  not g34087 (n_15941, n18427);
  not g34088 (n_15942, n18530);
  and g34089 (n18531, n_15941, n_15942);
  and g34090 (n18532, n18427, n_15940);
  and g34091 (n18533, n_15939, n18532);
  not g34092 (n_15943, n18531);
  not g34093 (n_15944, n18533);
  and g34094 (n18534, n_15943, n_15944);
  not g34095 (n_15945, n18193);
  and g34096 (n18535, n_15945, n18534);
  not g34097 (n_15946, n18534);
  and g34098 (n18536, n18193, n_15946);
  not g34099 (n_15947, n18535);
  not g34100 (n_15948, n18536);
  and g34101 (n18537, n_15947, n_15948);
  not g34102 (n_15949, n18416);
  and g34103 (n18538, n_15949, n18537);
  not g34104 (n_15950, n18537);
  and g34105 (n18539, n18416, n_15950);
  not g34106 (n_15951, n18538);
  not g34107 (n_15952, n18539);
  and g34108 (n18540, n_15951, n_15952);
  not g34109 (n_15953, n18405);
  and g34110 (n18541, n_15953, n18540);
  not g34111 (n_15954, n18541);
  and g34112 (n18542, n_15953, n_15954);
  and g34113 (n18543, n18540, n_15954);
  not g34114 (n_15955, n18542);
  not g34115 (n_15956, n18543);
  and g34116 (n18544, n_15955, n_15956);
  not g34117 (n_15957, n18403);
  not g34118 (n_15958, n18544);
  and g34119 (n18545, n_15957, n_15958);
  and g34120 (n18546, n18403, n_15956);
  and g34121 (n18547, n_15955, n18546);
  not g34122 (n_15959, n18545);
  not g34123 (n_15960, n18547);
  and g34124 (n18548, n_15959, n_15960);
  not g34125 (n_15961, n18392);
  and g34126 (n18549, n_15961, n18548);
  not g34127 (n_15962, n18549);
  and g34128 (n18550, n_15961, n_15962);
  and g34129 (n18551, n18548, n_15962);
  not g34130 (n_15963, n18550);
  not g34131 (n_15964, n18551);
  and g34132 (n18552, n_15963, n_15964);
  not g34133 (n_15965, n18391);
  not g34134 (n_15966, n18552);
  and g34135 (n18553, n_15965, n_15966);
  and g34136 (n18554, n18391, n_15964);
  and g34137 (n18555, n_15963, n18554);
  not g34138 (n_15967, n18553);
  not g34139 (n_15968, n18555);
  and g34140 (n18556, n_15967, n_15968);
  not g34141 (n_15969, n18380);
  and g34142 (n18557, n_15969, n18556);
  not g34143 (n_15970, n18556);
  and g34144 (n18558, n18380, n_15970);
  not g34145 (n_15971, n18557);
  not g34146 (n_15972, n18558);
  and g34147 (n18559, n_15971, n_15972);
  not g34148 (n_15973, n18378);
  and g34149 (n18560, n_15973, n18559);
  not g34150 (n_15974, n18560);
  and g34151 (n18561, n18559, n_15974);
  and g34152 (n18562, n_15973, n_15974);
  not g34153 (n_15975, n18561);
  not g34154 (n_15976, n18562);
  and g34155 (n18563, n_15975, n_15976);
  and g34156 (n18564, n_15716, n_15721);
  and g34157 (n18565, \b[46] , n3638);
  and g34158 (n18566, \b[44] , n3843);
  and g34159 (n18567, \b[45] , n3633);
  not g34160 (n_15977, n18566);
  not g34161 (n_15978, n18567);
  and g34162 (n18568, n_15977, n_15978);
  not g34163 (n_15979, n18565);
  and g34164 (n18569, n_15979, n18568);
  and g34165 (n18570, n_12780, n18569);
  and g34166 (n18571, n_13970, n18569);
  not g34167 (n_15980, n18570);
  not g34168 (n_15981, n18571);
  and g34169 (n18572, n_15980, n_15981);
  not g34170 (n_15982, n18572);
  and g34171 (n18573, \a[32] , n_15982);
  and g34172 (n18574, n_2992, n18572);
  not g34173 (n_15983, n18573);
  not g34174 (n_15984, n18574);
  and g34175 (n18575, n_15983, n_15984);
  not g34176 (n_15985, n18564);
  not g34177 (n_15986, n18575);
  and g34178 (n18576, n_15985, n_15986);
  not g34179 (n_15987, n18576);
  and g34180 (n18577, n_15985, n_15987);
  and g34181 (n18578, n_15986, n_15987);
  not g34182 (n_15988, n18577);
  not g34183 (n_15989, n18578);
  and g34184 (n18579, n_15988, n_15989);
  not g34185 (n_15990, n18563);
  not g34186 (n_15991, n18579);
  and g34187 (n18580, n_15990, n_15991);
  not g34188 (n_15992, n18580);
  and g34189 (n18581, n_15990, n_15992);
  and g34190 (n18582, n_15991, n_15992);
  not g34191 (n_15993, n18581);
  not g34192 (n_15994, n18582);
  and g34193 (n18583, n_15993, n_15994);
  not g34194 (n_15995, n18367);
  not g34195 (n_15996, n18583);
  and g34196 (n18584, n_15995, n_15996);
  not g34197 (n_15997, n18584);
  and g34198 (n18585, n_15995, n_15997);
  and g34199 (n18586, n_15996, n_15997);
  not g34200 (n_15998, n18585);
  not g34201 (n_15999, n18586);
  and g34202 (n18587, n_15998, n_15999);
  and g34203 (n18588, n_15544, n_15545);
  not g34204 (n_16000, n18588);
  and g34205 (n18589, n_15740, n_16000);
  and g34206 (n18590, \b[52] , n2539);
  and g34207 (n18591, \b[50] , n2685);
  and g34208 (n18592, \b[51] , n2534);
  not g34209 (n_16001, n18591);
  not g34210 (n_16002, n18592);
  and g34211 (n18593, n_16001, n_16002);
  not g34212 (n_16003, n18590);
  and g34213 (n18594, n_16003, n18593);
  and g34214 (n18595, n_13498, n18594);
  not g34215 (n_16004, n9628);
  and g34216 (n18596, n_16004, n18594);
  not g34217 (n_16005, n18595);
  not g34218 (n_16006, n18596);
  and g34219 (n18597, n_16005, n_16006);
  not g34220 (n_16007, n18597);
  and g34221 (n18598, \a[26] , n_16007);
  and g34222 (n18599, n_2025, n18597);
  not g34223 (n_16008, n18598);
  not g34224 (n_16009, n18599);
  and g34225 (n18600, n_16008, n_16009);
  not g34226 (n_16010, n18589);
  not g34227 (n_16011, n18600);
  and g34228 (n18601, n_16010, n_16011);
  and g34229 (n18602, n18589, n18600);
  not g34230 (n_16012, n18601);
  not g34231 (n_16013, n18602);
  and g34232 (n18603, n_16012, n_16013);
  not g34233 (n_16014, n18587);
  and g34234 (n18604, n_16014, n18603);
  not g34235 (n_16015, n18604);
  and g34236 (n18605, n_16014, n_16015);
  and g34237 (n18606, n18603, n_16015);
  not g34238 (n_16016, n18605);
  not g34239 (n_16017, n18606);
  and g34240 (n18607, n_16016, n_16017);
  not g34241 (n_16018, n18351);
  not g34242 (n_16019, n18607);
  and g34243 (n18608, n_16018, n_16019);
  not g34244 (n_16020, n18608);
  and g34245 (n18609, n_16018, n_16020);
  and g34246 (n18610, n_16019, n_16020);
  not g34247 (n_16021, n18609);
  not g34248 (n_16022, n18610);
  and g34249 (n18611, n_16021, n_16022);
  and g34250 (n18612, n_15521, n_15748);
  and g34251 (n18613, \b[58] , n1627);
  and g34252 (n18614, \b[56] , n1763);
  and g34253 (n18615, \b[57] , n1622);
  not g34254 (n_16023, n18614);
  not g34255 (n_16024, n18615);
  and g34256 (n18616, n_16023, n_16024);
  not g34257 (n_16025, n18613);
  and g34258 (n18617, n_16025, n18616);
  and g34259 (n18618, n_14471, n18617);
  and g34260 (n18619, n_13160, n18617);
  not g34261 (n_16026, n18618);
  not g34262 (n_16027, n18619);
  and g34263 (n18620, n_16026, n_16027);
  not g34264 (n_16028, n18620);
  and g34265 (n18621, \a[20] , n_16028);
  and g34266 (n18622, n_1221, n18620);
  not g34267 (n_16029, n18621);
  not g34268 (n_16030, n18622);
  and g34269 (n18623, n_16029, n_16030);
  not g34270 (n_16031, n18612);
  not g34271 (n_16032, n18623);
  and g34272 (n18624, n_16031, n_16032);
  not g34273 (n_16033, n18624);
  and g34274 (n18625, n_16031, n_16033);
  and g34275 (n18626, n_16032, n_16033);
  not g34276 (n_16034, n18625);
  not g34277 (n_16035, n18626);
  and g34278 (n18627, n_16034, n_16035);
  not g34279 (n_16036, n18611);
  not g34280 (n_16037, n18627);
  and g34281 (n18628, n_16036, n_16037);
  not g34282 (n_16038, n18628);
  and g34283 (n18629, n_16036, n_16038);
  and g34284 (n18630, n_16037, n_16038);
  not g34285 (n_16039, n18629);
  not g34286 (n_16040, n18630);
  and g34287 (n18631, n_16039, n_16040);
  not g34288 (n_16041, n18335);
  not g34289 (n_16042, n18631);
  and g34290 (n18632, n_16041, n_16042);
  not g34291 (n_16043, n18632);
  and g34292 (n18633, n_16041, n_16043);
  and g34293 (n18634, n_16042, n_16043);
  not g34294 (n_16044, n18633);
  not g34295 (n_16045, n18634);
  and g34296 (n18635, n_16044, n_16045);
  and g34297 (n18636, n_15495, n_15496);
  not g34298 (n_16046, n18636);
  and g34299 (n18637, n_15756, n_16046);
  and g34300 (n18638, \b[62] , n1056);
  and g34301 (n18639, \b[63] , n946);
  not g34302 (n_16047, n18638);
  not g34303 (n_16048, n18639);
  and g34304 (n18640, n_16047, n_16048);
  and g34305 (n18641, n_12819, n18640);
  and g34306 (n18642, n13800, n18640);
  not g34307 (n_16049, n18641);
  not g34308 (n_16050, n18642);
  and g34309 (n18643, n_16049, n_16050);
  not g34310 (n_16051, n18643);
  and g34311 (n18644, \a[14] , n_16051);
  and g34312 (n18645, n_623, n18643);
  not g34313 (n_16052, n18644);
  not g34314 (n_16053, n18645);
  and g34315 (n18646, n_16052, n_16053);
  not g34316 (n_16054, n18637);
  not g34317 (n_16055, n18646);
  and g34318 (n18647, n_16054, n_16055);
  not g34319 (n_16056, n18647);
  and g34320 (n18648, n_16054, n_16056);
  and g34321 (n18649, n_16055, n_16056);
  not g34322 (n_16057, n18648);
  not g34323 (n_16058, n18649);
  and g34324 (n18650, n_16057, n_16058);
  not g34325 (n_16059, n18635);
  not g34326 (n_16060, n18650);
  and g34327 (n18651, n_16059, n_16060);
  and g34328 (n18652, n18635, n_16058);
  and g34329 (n18653, n_16057, n18652);
  not g34330 (n_16061, n18651);
  not g34331 (n_16062, n18653);
  and g34332 (n18654, n_16061, n_16062);
  not g34333 (n_16063, n18319);
  and g34334 (n18655, n_16063, n18654);
  not g34335 (n_16064, n18655);
  and g34336 (n18656, n_16063, n_16064);
  and g34337 (n18657, n18654, n_16064);
  not g34338 (n_16065, n18656);
  not g34339 (n_16066, n18657);
  and g34340 (n18658, n_16065, n_16066);
  not g34341 (n_16067, n18317);
  not g34342 (n_16068, n18658);
  and g34343 (n18659, n_16067, n_16068);
  and g34344 (n18660, n18317, n_16066);
  and g34345 (n18661, n_16065, n18660);
  not g34346 (n_16069, n18659);
  not g34347 (n_16070, n18661);
  and g34348 (\f[76] , n_16069, n_16070);
  and g34349 (n18663, n_16064, n_16069);
  and g34350 (n18664, n_16056, n_16061);
  and g34351 (n18665, n_15783, n_16043);
  and g34352 (n18666, \b[63] , n1056);
  and g34353 (n18667, n954, n13797);
  not g34354 (n_16071, n18666);
  not g34355 (n_16072, n18667);
  and g34356 (n18668, n_16071, n_16072);
  not g34357 (n_16073, n18668);
  and g34358 (n18669, \a[14] , n_16073);
  not g34359 (n_16074, n18669);
  and g34360 (n18670, \a[14] , n_16074);
  and g34361 (n18671, n_16073, n_16074);
  not g34362 (n_16075, n18670);
  not g34363 (n_16076, n18671);
  and g34364 (n18672, n_16075, n_16076);
  not g34365 (n_16077, n18665);
  not g34366 (n_16078, n18672);
  and g34367 (n18673, n_16077, n_16078);
  not g34368 (n_16079, n18673);
  and g34369 (n18674, n_16077, n_16079);
  and g34370 (n18675, n_16078, n_16079);
  not g34371 (n_16080, n18674);
  not g34372 (n_16081, n18675);
  and g34373 (n18676, n_16080, n_16081);
  and g34374 (n18677, \b[59] , n1627);
  and g34375 (n18678, \b[57] , n1763);
  and g34376 (n18679, \b[58] , n1622);
  and g34382 (n18682, n1630, n12179);
  not g34385 (n_16086, n18683);
  and g34386 (n18684, \a[20] , n_16086);
  not g34387 (n_16087, n18684);
  and g34388 (n18685, \a[20] , n_16087);
  and g34389 (n18686, n_16086, n_16087);
  not g34390 (n_16088, n18685);
  not g34391 (n_16089, n18686);
  and g34392 (n18687, n_16088, n_16089);
  and g34393 (n18688, n_15796, n_16020);
  and g34394 (n18689, n18687, n18688);
  not g34395 (n_16090, n18687);
  not g34396 (n_16091, n18688);
  and g34397 (n18690, n_16090, n_16091);
  not g34398 (n_16092, n18689);
  not g34399 (n_16093, n18690);
  and g34400 (n18691, n_16092, n_16093);
  and g34401 (n18692, \b[56] , n2048);
  and g34402 (n18693, \b[54] , n2198);
  and g34403 (n18694, \b[55] , n2043);
  and g34409 (n18697, n2051, n10708);
  not g34412 (n_16098, n18698);
  and g34413 (n18699, \a[23] , n_16098);
  not g34414 (n_16099, n18699);
  and g34415 (n18700, \a[23] , n_16099);
  and g34416 (n18701, n_16098, n_16099);
  not g34417 (n_16100, n18700);
  not g34418 (n_16101, n18701);
  and g34419 (n18702, n_16100, n_16101);
  and g34420 (n18703, n_16012, n_16015);
  and g34421 (n18704, n18702, n18703);
  not g34422 (n_16102, n18702);
  not g34423 (n_16103, n18703);
  and g34424 (n18705, n_16102, n_16103);
  not g34425 (n_16104, n18704);
  not g34426 (n_16105, n18705);
  and g34427 (n18706, n_16104, n_16105);
  and g34428 (n18707, \b[53] , n2539);
  and g34429 (n18708, \b[51] , n2685);
  and g34430 (n18709, \b[52] , n2534);
  and g34436 (n18712, n2542, n9972);
  not g34439 (n_16110, n18713);
  and g34440 (n18714, \a[26] , n_16110);
  not g34441 (n_16111, n18714);
  and g34442 (n18715, \a[26] , n_16111);
  and g34443 (n18716, n_16110, n_16111);
  not g34444 (n_16112, n18715);
  not g34445 (n_16113, n18716);
  and g34446 (n18717, n_16112, n_16113);
  and g34447 (n18718, n_15809, n_15997);
  and g34448 (n18719, n18717, n18718);
  not g34449 (n_16114, n18717);
  not g34450 (n_16115, n18718);
  and g34451 (n18720, n_16114, n_16115);
  not g34452 (n_16116, n18719);
  not g34453 (n_16117, n18720);
  and g34454 (n18721, n_16116, n_16117);
  and g34455 (n18722, n_15971, n_15974);
  and g34456 (n18723, \b[47] , n3638);
  and g34457 (n18724, \b[45] , n3843);
  and g34458 (n18725, \b[46] , n3633);
  not g34459 (n_16118, n18724);
  not g34460 (n_16119, n18725);
  and g34461 (n18726, n_16118, n_16119);
  not g34462 (n_16120, n18723);
  and g34463 (n18727, n_16120, n18726);
  and g34464 (n18728, n_12780, n18727);
  not g34465 (n_16121, n7703);
  and g34466 (n18729, n_16121, n18727);
  not g34467 (n_16122, n18728);
  not g34468 (n_16123, n18729);
  and g34469 (n18730, n_16122, n_16123);
  not g34470 (n_16124, n18730);
  and g34471 (n18731, \a[32] , n_16124);
  and g34472 (n18732, n_2992, n18730);
  not g34473 (n_16125, n18731);
  not g34474 (n_16126, n18732);
  and g34475 (n18733, n_16125, n_16126);
  not g34476 (n_16127, n18722);
  not g34477 (n_16128, n18733);
  and g34478 (n18734, n_16127, n_16128);
  and g34479 (n18735, n18722, n18733);
  not g34480 (n_16129, n18734);
  not g34481 (n_16130, n18735);
  and g34482 (n18736, n_16129, n_16130);
  and g34483 (n18737, \b[44] , n4287);
  and g34484 (n18738, \b[42] , n4532);
  and g34485 (n18739, \b[43] , n4282);
  and g34491 (n18742, n4290, n7072);
  not g34494 (n_16135, n18743);
  and g34495 (n18744, \a[35] , n_16135);
  not g34496 (n_16136, n18744);
  and g34497 (n18745, \a[35] , n_16136);
  and g34498 (n18746, n_16135, n_16136);
  not g34499 (n_16137, n18745);
  not g34500 (n_16138, n18746);
  and g34501 (n18747, n_16137, n_16138);
  and g34502 (n18748, n_15962, n_15967);
  and g34503 (n18749, \b[41] , n5035);
  and g34504 (n18750, \b[39] , n5277);
  and g34505 (n18751, \b[40] , n5030);
  and g34511 (n18754, n5038, n6219);
  not g34514 (n_16143, n18755);
  and g34515 (n18756, \a[38] , n_16143);
  not g34516 (n_16144, n18756);
  and g34517 (n18757, \a[38] , n_16144);
  and g34518 (n18758, n_16143, n_16144);
  not g34519 (n_16145, n18757);
  not g34520 (n_16146, n18758);
  and g34521 (n18759, n_16145, n_16146);
  and g34522 (n18760, n_15954, n_15959);
  and g34523 (n18761, n_15938, n_15943);
  and g34524 (n18762, n_15908, n_15918);
  and g34525 (n18763, \b[26] , n9339);
  and g34526 (n18764, \b[24] , n9732);
  and g34527 (n18765, \b[25] , n9334);
  and g34533 (n18768, n2813, n9342);
  not g34536 (n_16151, n18769);
  and g34537 (n18770, \a[53] , n_16151);
  not g34538 (n_16152, n18770);
  and g34539 (n18771, \a[53] , n_16152);
  and g34540 (n18772, n_16151, n_16152);
  not g34541 (n_16153, n18771);
  not g34542 (n_16154, n18772);
  and g34543 (n18773, n_16153, n_16154);
  and g34544 (n18774, n_15892, n_15902);
  and g34545 (n18775, n_15869, n_15870);
  not g34546 (n_16155, n18775);
  and g34547 (n18776, n_15858, n_16155);
  and g34548 (n18777, \b[13] , n13903);
  and g34549 (n18778, \b[14] , n_11555);
  not g34550 (n_16156, n18777);
  not g34551 (n_16157, n18778);
  and g34552 (n18779, n_16156, n_16157);
  not g34553 (n_16158, n18779);
  and g34554 (n18780, n18431, n_16158);
  not g34555 (n_16159, n18431);
  and g34556 (n18781, n_16159, n18779);
  not g34557 (n_16160, n18780);
  not g34558 (n_16161, n18781);
  and g34559 (n18782, n_16160, n_16161);
  and g34560 (n18783, \b[17] , n12668);
  and g34561 (n18784, \b[15] , n13047);
  and g34562 (n18785, \b[16] , n12663);
  not g34563 (n_16162, n18784);
  not g34564 (n_16163, n18785);
  and g34565 (n18786, n_16162, n_16163);
  not g34566 (n_16164, n18783);
  and g34567 (n18787, n_16164, n18786);
  and g34568 (n18788, n_12644, n18787);
  not g34569 (n_16165, n1356);
  and g34570 (n18789, n_16165, n18787);
  not g34571 (n_16166, n18788);
  not g34572 (n_16167, n18789);
  and g34573 (n18790, n_16166, n_16167);
  not g34574 (n_16168, n18790);
  and g34575 (n18791, \a[62] , n_16168);
  and g34576 (n18792, n_10843, n18790);
  not g34577 (n_16169, n18791);
  not g34578 (n_16170, n18792);
  and g34579 (n18793, n_16169, n_16170);
  not g34580 (n_16171, n18793);
  and g34581 (n18794, n18782, n_16171);
  not g34582 (n_16172, n18782);
  and g34583 (n18795, n_16172, n18793);
  not g34584 (n_16173, n18794);
  not g34585 (n_16174, n18795);
  and g34586 (n18796, n_16173, n_16174);
  not g34587 (n_16175, n18776);
  and g34588 (n18797, n_16175, n18796);
  not g34589 (n_16176, n18796);
  and g34590 (n18798, n18776, n_16176);
  not g34591 (n_16177, n18797);
  not g34592 (n_16178, n18798);
  and g34593 (n18799, n_16177, n_16178);
  and g34594 (n18800, \b[20] , n11531);
  and g34595 (n18801, \b[18] , n11896);
  and g34596 (n18802, \b[19] , n11526);
  and g34602 (n18805, n1846, n11534);
  not g34605 (n_16183, n18806);
  and g34606 (n18807, \a[59] , n_16183);
  not g34607 (n_16184, n18807);
  and g34608 (n18808, \a[59] , n_16184);
  and g34609 (n18809, n_16183, n_16184);
  not g34610 (n_16185, n18808);
  not g34611 (n_16186, n18809);
  and g34612 (n18810, n_16185, n_16186);
  not g34613 (n_16187, n18810);
  and g34614 (n18811, n18799, n_16187);
  not g34615 (n_16188, n18811);
  and g34616 (n18812, n18799, n_16188);
  and g34617 (n18813, n_16187, n_16188);
  not g34618 (n_16189, n18812);
  not g34619 (n_16190, n18813);
  and g34620 (n18814, n_16189, n_16190);
  and g34621 (n18815, n_15876, n_15886);
  and g34622 (n18816, n18814, n18815);
  not g34623 (n_16191, n18814);
  not g34624 (n_16192, n18815);
  and g34625 (n18817, n_16191, n_16192);
  not g34626 (n_16193, n18816);
  not g34627 (n_16194, n18817);
  and g34628 (n18818, n_16193, n_16194);
  and g34629 (n18819, \b[23] , n10426);
  and g34630 (n18820, \b[21] , n10796);
  and g34631 (n18821, \b[22] , n10421);
  and g34637 (n18824, n2300, n10429);
  not g34640 (n_16199, n18825);
  and g34641 (n18826, \a[56] , n_16199);
  not g34642 (n_16200, n18826);
  and g34643 (n18827, \a[56] , n_16200);
  and g34644 (n18828, n_16199, n_16200);
  not g34645 (n_16201, n18827);
  not g34646 (n_16202, n18828);
  and g34647 (n18829, n_16201, n_16202);
  not g34648 (n_16203, n18818);
  and g34649 (n18830, n_16203, n18829);
  not g34650 (n_16204, n18829);
  and g34651 (n18831, n18818, n_16204);
  not g34652 (n_16205, n18830);
  not g34653 (n_16206, n18831);
  and g34654 (n18832, n_16205, n_16206);
  not g34655 (n_16207, n18774);
  and g34656 (n18833, n_16207, n18832);
  not g34657 (n_16208, n18832);
  and g34658 (n18834, n18774, n_16208);
  not g34659 (n_16209, n18833);
  not g34660 (n_16210, n18834);
  and g34661 (n18835, n_16209, n_16210);
  not g34662 (n_16211, n18773);
  and g34663 (n18836, n_16211, n18835);
  not g34664 (n_16212, n18835);
  and g34665 (n18837, n18773, n_16212);
  not g34666 (n_16213, n18836);
  not g34667 (n_16214, n18837);
  and g34668 (n18838, n_16213, n_16214);
  not g34669 (n_16215, n18762);
  and g34670 (n18839, n_16215, n18838);
  not g34671 (n_16216, n18838);
  and g34672 (n18840, n18762, n_16216);
  not g34673 (n_16217, n18839);
  not g34674 (n_16218, n18840);
  and g34675 (n18841, n_16217, n_16218);
  and g34676 (n18842, \b[29] , n8362);
  and g34677 (n18843, \b[27] , n8715);
  and g34678 (n18844, \b[28] , n8357);
  and g34684 (n18847, n3383, n8365);
  not g34687 (n_16223, n18848);
  and g34688 (n18849, \a[50] , n_16223);
  not g34689 (n_16224, n18849);
  and g34690 (n18850, \a[50] , n_16224);
  and g34691 (n18851, n_16223, n_16224);
  not g34692 (n_16225, n18850);
  not g34693 (n_16226, n18851);
  and g34694 (n18852, n_16225, n_16226);
  not g34695 (n_16227, n18852);
  and g34696 (n18853, n18841, n_16227);
  not g34697 (n_16228, n18853);
  and g34698 (n18854, n18841, n_16228);
  and g34699 (n18855, n_16227, n_16228);
  not g34700 (n_16229, n18854);
  not g34701 (n_16230, n18855);
  and g34702 (n18856, n_16229, n_16230);
  and g34703 (n18857, n_15924, n_15936);
  not g34704 (n_16231, n18856);
  not g34705 (n_16232, n18857);
  and g34706 (n18858, n_16231, n_16232);
  not g34707 (n_16233, n18858);
  and g34708 (n18859, n_16231, n_16233);
  and g34709 (n18860, n_16232, n_16233);
  not g34710 (n_16234, n18859);
  not g34711 (n_16235, n18860);
  and g34712 (n18861, n_16234, n_16235);
  and g34713 (n18862, \b[32] , n7446);
  and g34714 (n18863, \b[30] , n7787);
  and g34715 (n18864, \b[31] , n7441);
  and g34721 (n18867, n4013, n7449);
  not g34724 (n_16240, n18868);
  and g34725 (n18869, \a[47] , n_16240);
  not g34726 (n_16241, n18869);
  and g34727 (n18870, \a[47] , n_16241);
  and g34728 (n18871, n_16240, n_16241);
  not g34729 (n_16242, n18870);
  not g34730 (n_16243, n18871);
  and g34731 (n18872, n_16242, n_16243);
  not g34732 (n_16244, n18861);
  and g34733 (n18873, n_16244, n18872);
  not g34734 (n_16245, n18872);
  and g34735 (n18874, n18861, n_16245);
  not g34736 (n_16246, n18873);
  not g34737 (n_16247, n18874);
  and g34738 (n18875, n_16246, n_16247);
  and g34739 (n18876, n18761, n18875);
  not g34740 (n_16248, n18761);
  not g34741 (n_16249, n18875);
  and g34742 (n18877, n_16248, n_16249);
  not g34743 (n_16250, n18876);
  not g34744 (n_16251, n18877);
  and g34745 (n18878, n_16250, n_16251);
  and g34746 (n18879, \b[35] , n6595);
  and g34747 (n18880, \b[33] , n6902);
  and g34748 (n18881, \b[34] , n6590);
  and g34754 (n18884, n4696, n6598);
  not g34757 (n_16256, n18885);
  and g34758 (n18886, \a[44] , n_16256);
  not g34759 (n_16257, n18886);
  and g34760 (n18887, \a[44] , n_16257);
  and g34761 (n18888, n_16256, n_16257);
  not g34762 (n_16258, n18887);
  not g34763 (n_16259, n18888);
  and g34764 (n18889, n_16258, n_16259);
  not g34765 (n_16260, n18889);
  and g34766 (n18890, n18878, n_16260);
  not g34767 (n_16261, n18890);
  and g34768 (n18891, n18878, n_16261);
  and g34769 (n18892, n_16260, n_16261);
  not g34770 (n_16262, n18891);
  not g34771 (n_16263, n18892);
  and g34772 (n18893, n_16262, n_16263);
  and g34773 (n18894, n_15947, n_15951);
  and g34774 (n18895, n18893, n18894);
  not g34775 (n_16264, n18893);
  not g34776 (n_16265, n18894);
  and g34777 (n18896, n_16264, n_16265);
  not g34778 (n_16266, n18895);
  not g34779 (n_16267, n18896);
  and g34780 (n18897, n_16266, n_16267);
  and g34781 (n18898, \b[38] , n5777);
  and g34782 (n18899, \b[36] , n6059);
  and g34783 (n18900, \b[37] , n5772);
  and g34789 (n18903, n5205, n5780);
  not g34792 (n_16272, n18904);
  and g34793 (n18905, \a[41] , n_16272);
  not g34794 (n_16273, n18905);
  and g34795 (n18906, \a[41] , n_16273);
  and g34796 (n18907, n_16272, n_16273);
  not g34797 (n_16274, n18906);
  not g34798 (n_16275, n18907);
  and g34799 (n18908, n_16274, n_16275);
  not g34800 (n_16276, n18897);
  and g34801 (n18909, n_16276, n18908);
  not g34802 (n_16277, n18908);
  and g34803 (n18910, n18897, n_16277);
  not g34804 (n_16278, n18909);
  not g34805 (n_16279, n18910);
  and g34806 (n18911, n_16278, n_16279);
  not g34807 (n_16280, n18760);
  and g34808 (n18912, n_16280, n18911);
  not g34809 (n_16281, n18911);
  and g34810 (n18913, n18760, n_16281);
  not g34811 (n_16282, n18912);
  not g34812 (n_16283, n18913);
  and g34813 (n18914, n_16282, n_16283);
  not g34814 (n_16284, n18759);
  and g34815 (n18915, n_16284, n18914);
  not g34816 (n_16285, n18914);
  and g34817 (n18916, n18759, n_16285);
  not g34818 (n_16286, n18915);
  not g34819 (n_16287, n18916);
  and g34820 (n18917, n_16286, n_16287);
  not g34821 (n_16288, n18748);
  and g34822 (n18918, n_16288, n18917);
  not g34823 (n_16289, n18917);
  and g34824 (n18919, n18748, n_16289);
  not g34825 (n_16290, n18918);
  not g34826 (n_16291, n18919);
  and g34827 (n18920, n_16290, n_16291);
  not g34828 (n_16292, n18747);
  and g34829 (n18921, n_16292, n18920);
  not g34830 (n_16293, n18921);
  and g34831 (n18922, n_16292, n_16293);
  and g34832 (n18923, n18920, n_16293);
  not g34833 (n_16294, n18922);
  not g34834 (n_16295, n18923);
  and g34835 (n18924, n_16294, n_16295);
  not g34836 (n_16296, n18924);
  and g34837 (n18925, n18736, n_16296);
  not g34838 (n_16297, n18925);
  and g34839 (n18926, n18736, n_16297);
  and g34840 (n18927, n_16296, n_16297);
  not g34841 (n_16298, n18926);
  not g34842 (n_16299, n18927);
  and g34843 (n18928, n_16298, n_16299);
  and g34844 (n18929, n_15987, n_15992);
  and g34845 (n18930, \b[50] , n3050);
  and g34846 (n18931, \b[48] , n3243);
  and g34847 (n18932, \b[49] , n3045);
  not g34848 (n_16300, n18931);
  not g34849 (n_16301, n18932);
  and g34850 (n18933, n_16300, n_16301);
  not g34851 (n_16302, n18930);
  and g34852 (n18934, n_16302, n18933);
  and g34853 (n18935, n_12601, n18934);
  and g34854 (n18936, n_15219, n18934);
  not g34855 (n_16303, n18935);
  not g34856 (n_16304, n18936);
  and g34857 (n18937, n_16303, n_16304);
  not g34858 (n_16305, n18937);
  and g34859 (n18938, \a[29] , n_16305);
  and g34860 (n18939, n_2476, n18937);
  not g34861 (n_16306, n18938);
  not g34862 (n_16307, n18939);
  and g34863 (n18940, n_16306, n_16307);
  not g34864 (n_16308, n18929);
  not g34865 (n_16309, n18940);
  and g34866 (n18941, n_16308, n_16309);
  and g34867 (n18942, n18929, n18940);
  not g34868 (n_16310, n18941);
  not g34869 (n_16311, n18942);
  and g34870 (n18943, n_16310, n_16311);
  not g34871 (n_16312, n18928);
  and g34872 (n18944, n_16312, n18943);
  not g34873 (n_16313, n18944);
  and g34874 (n18945, n_16312, n_16313);
  and g34875 (n18946, n18943, n_16313);
  not g34876 (n_16314, n18945);
  not g34877 (n_16315, n18946);
  and g34878 (n18947, n_16314, n_16315);
  not g34879 (n_16316, n18947);
  and g34880 (n18948, n18721, n_16316);
  not g34881 (n_16317, n18948);
  and g34882 (n18949, n18721, n_16317);
  and g34883 (n18950, n_16316, n_16317);
  not g34884 (n_16318, n18949);
  not g34885 (n_16319, n18950);
  and g34886 (n18951, n_16318, n_16319);
  not g34887 (n_16320, n18951);
  and g34888 (n18952, n18706, n_16320);
  not g34889 (n_16321, n18706);
  and g34890 (n18953, n_16321, n18951);
  not g34891 (n_16322, n18953);
  and g34892 (n18954, n18691, n_16322);
  not g34893 (n_16323, n18952);
  and g34894 (n18955, n_16323, n18954);
  not g34895 (n_16324, n18955);
  and g34896 (n18956, n18691, n_16324);
  and g34897 (n18957, n_16322, n_16324);
  and g34898 (n18958, n_16323, n18957);
  not g34899 (n_16325, n18956);
  not g34900 (n_16326, n18958);
  and g34901 (n18959, n_16325, n_16326);
  and g34902 (n18960, n_16033, n_16038);
  and g34903 (n18961, \b[62] , n1302);
  and g34904 (n18962, \b[60] , n1391);
  and g34905 (n18963, \b[61] , n1297);
  not g34906 (n_16327, n18962);
  not g34907 (n_16328, n18963);
  and g34908 (n18964, n_16327, n_16328);
  not g34909 (n_16329, n18961);
  and g34910 (n18965, n_16329, n18964);
  and g34911 (n18966, n_13260, n18965);
  and g34912 (n18967, n_13538, n18965);
  not g34913 (n_16330, n18966);
  not g34914 (n_16331, n18967);
  and g34915 (n18968, n_16330, n_16331);
  not g34916 (n_16332, n18968);
  and g34917 (n18969, \a[17] , n_16332);
  and g34918 (n18970, n_926, n18968);
  not g34919 (n_16333, n18969);
  not g34920 (n_16334, n18970);
  and g34921 (n18971, n_16333, n_16334);
  not g34922 (n_16335, n18960);
  not g34923 (n_16336, n18971);
  and g34924 (n18972, n_16335, n_16336);
  not g34925 (n_16337, n18972);
  and g34926 (n18973, n_16335, n_16337);
  and g34927 (n18974, n_16336, n_16337);
  not g34928 (n_16338, n18973);
  not g34929 (n_16339, n18974);
  and g34930 (n18975, n_16338, n_16339);
  not g34931 (n_16340, n18959);
  not g34932 (n_16341, n18975);
  and g34933 (n18976, n_16340, n_16341);
  and g34934 (n18977, n18959, n_16339);
  and g34935 (n18978, n_16338, n18977);
  not g34936 (n_16342, n18976);
  not g34937 (n_16343, n18978);
  and g34938 (n18979, n_16342, n_16343);
  not g34939 (n_16344, n18676);
  and g34940 (n18980, n_16344, n18979);
  not g34941 (n_16345, n18979);
  and g34942 (n18981, n18676, n_16345);
  not g34943 (n_16346, n18980);
  not g34944 (n_16347, n18981);
  and g34945 (n18982, n_16346, n_16347);
  not g34946 (n_16348, n18664);
  and g34947 (n18983, n_16348, n18982);
  not g34948 (n_16349, n18982);
  and g34949 (n18984, n18664, n_16349);
  not g34950 (n_16350, n18983);
  not g34951 (n_16351, n18984);
  and g34952 (n18985, n_16350, n_16351);
  not g34953 (n_16352, n18663);
  and g34954 (n18986, n_16352, n18985);
  not g34955 (n_16353, n18985);
  and g34956 (n18987, n18663, n_16353);
  not g34957 (n_16354, n18986);
  not g34958 (n_16355, n18987);
  and g34959 (\f[77] , n_16354, n_16355);
  and g34960 (n18989, n_16337, n_16342);
  and g34961 (n18990, \b[63] , n1302);
  and g34962 (n18991, \b[61] , n1391);
  and g34963 (n18992, \b[62] , n1297);
  and g34969 (n18995, n1305, n13771);
  not g34972 (n_16360, n18996);
  and g34973 (n18997, \a[17] , n_16360);
  not g34974 (n_16361, n18997);
  and g34975 (n18998, \a[17] , n_16361);
  and g34976 (n18999, n_16360, n_16361);
  not g34977 (n_16362, n18998);
  not g34978 (n_16363, n18999);
  and g34979 (n19000, n_16362, n_16363);
  not g34980 (n_16364, n18989);
  not g34981 (n_16365, n19000);
  and g34982 (n19001, n_16364, n_16365);
  not g34983 (n_16366, n19001);
  and g34984 (n19002, n_16364, n_16366);
  and g34985 (n19003, n_16365, n_16366);
  not g34986 (n_16367, n19002);
  not g34987 (n_16368, n19003);
  and g34988 (n19004, n_16367, n_16368);
  and g34989 (n19005, \b[60] , n1627);
  and g34990 (n19006, \b[58] , n1763);
  and g34991 (n19007, \b[59] , n1622);
  and g34997 (n19010, n1630, n12211);
  not g35000 (n_16373, n19011);
  and g35001 (n19012, \a[20] , n_16373);
  not g35002 (n_16374, n19012);
  and g35003 (n19013, \a[20] , n_16374);
  and g35004 (n19014, n_16373, n_16374);
  not g35005 (n_16375, n19013);
  not g35006 (n_16376, n19014);
  and g35007 (n19015, n_16375, n_16376);
  and g35008 (n19016, n_16093, n_16324);
  and g35009 (n19017, n19015, n19016);
  not g35010 (n_16377, n19015);
  not g35011 (n_16378, n19016);
  and g35012 (n19018, n_16377, n_16378);
  not g35013 (n_16379, n19017);
  not g35014 (n_16380, n19018);
  and g35015 (n19019, n_16379, n_16380);
  and g35016 (n19020, n_16105, n_16323);
  and g35017 (n19021, \b[57] , n2048);
  and g35018 (n19022, \b[55] , n2198);
  and g35019 (n19023, \b[56] , n2043);
  and g35025 (n19026, n2051, n11410);
  not g35028 (n_16385, n19027);
  and g35029 (n19028, \a[23] , n_16385);
  not g35030 (n_16386, n19028);
  and g35031 (n19029, \a[23] , n_16386);
  and g35032 (n19030, n_16385, n_16386);
  not g35033 (n_16387, n19029);
  not g35034 (n_16388, n19030);
  and g35035 (n19031, n_16387, n_16388);
  not g35036 (n_16389, n19020);
  and g35037 (n19032, n_16389, n19031);
  not g35038 (n_16390, n19031);
  and g35039 (n19033, n19020, n_16390);
  not g35040 (n_16391, n19032);
  not g35041 (n_16392, n19033);
  and g35042 (n19034, n_16391, n_16392);
  and g35043 (n19035, \b[54] , n2539);
  and g35044 (n19036, \b[52] , n2685);
  and g35045 (n19037, \b[53] , n2534);
  and g35051 (n19040, n2542, n9998);
  not g35054 (n_16397, n19041);
  and g35055 (n19042, \a[26] , n_16397);
  not g35056 (n_16398, n19042);
  and g35057 (n19043, \a[26] , n_16398);
  and g35058 (n19044, n_16397, n_16398);
  not g35059 (n_16399, n19043);
  not g35060 (n_16400, n19044);
  and g35061 (n19045, n_16399, n_16400);
  and g35062 (n19046, n_16117, n_16317);
  and g35063 (n19047, n19045, n19046);
  not g35064 (n_16401, n19045);
  not g35065 (n_16402, n19046);
  and g35066 (n19048, n_16401, n_16402);
  not g35067 (n_16403, n19047);
  not g35068 (n_16404, n19048);
  and g35069 (n19049, n_16403, n_16404);
  and g35070 (n19050, \b[51] , n3050);
  and g35071 (n19051, \b[49] , n3243);
  and g35072 (n19052, \b[50] , n3045);
  and g35078 (n19055, n3053, n8976);
  not g35081 (n_16409, n19056);
  and g35082 (n19057, \a[29] , n_16409);
  not g35083 (n_16410, n19057);
  and g35084 (n19058, \a[29] , n_16410);
  and g35085 (n19059, n_16409, n_16410);
  not g35086 (n_16411, n19058);
  not g35087 (n_16412, n19059);
  and g35088 (n19060, n_16411, n_16412);
  and g35089 (n19061, n_16310, n_16313);
  and g35090 (n19062, n19060, n19061);
  not g35091 (n_16413, n19060);
  not g35092 (n_16414, n19061);
  and g35093 (n19063, n_16413, n_16414);
  not g35094 (n_16415, n19062);
  not g35095 (n_16416, n19063);
  and g35096 (n19064, n_16415, n_16416);
  and g35097 (n19065, n_16282, n_16286);
  and g35098 (n19066, n_16267, n_16279);
  and g35099 (n19067, n_16251, n_16261);
  and g35100 (n19068, n_16244, n_16245);
  not g35101 (n_16417, n19068);
  and g35102 (n19069, n_16233, n_16417);
  and g35103 (n19070, n_16194, n_16206);
  and g35104 (n19071, \b[14] , n13903);
  and g35105 (n19072, \b[15] , n_11555);
  not g35106 (n_16418, n19071);
  not g35107 (n_16419, n19072);
  and g35108 (n19073, n_16418, n_16419);
  not g35109 (n_16420, n19073);
  and g35110 (n19074, n_623, n_16420);
  not g35111 (n_16421, n19074);
  and g35112 (n19075, n_623, n_16421);
  and g35113 (n19076, n_16420, n_16421);
  not g35114 (n_16422, n19075);
  not g35115 (n_16423, n19076);
  and g35116 (n19077, n_16422, n_16423);
  not g35117 (n_16424, n19077);
  and g35118 (n19078, n_16159, n_16424);
  not g35119 (n_16425, n19078);
  and g35120 (n19079, n_16159, n_16425);
  and g35121 (n19080, n_16424, n_16425);
  not g35122 (n_16426, n19079);
  not g35123 (n_16427, n19080);
  and g35124 (n19081, n_16426, n_16427);
  and g35125 (n19082, \b[18] , n12668);
  and g35126 (n19083, \b[16] , n13047);
  and g35127 (n19084, \b[17] , n12663);
  and g35133 (n19087, n1566, n12671);
  not g35136 (n_16432, n19088);
  and g35137 (n19089, \a[62] , n_16432);
  not g35138 (n_16433, n19089);
  and g35139 (n19090, \a[62] , n_16433);
  and g35140 (n19091, n_16432, n_16433);
  not g35141 (n_16434, n19090);
  not g35142 (n_16435, n19091);
  and g35143 (n19092, n_16434, n_16435);
  not g35144 (n_16436, n19081);
  not g35145 (n_16437, n19092);
  and g35146 (n19093, n_16436, n_16437);
  not g35147 (n_16438, n19093);
  and g35148 (n19094, n_16436, n_16438);
  and g35149 (n19095, n_16437, n_16438);
  not g35150 (n_16439, n19094);
  not g35151 (n_16440, n19095);
  and g35152 (n19096, n_16439, n_16440);
  and g35153 (n19097, n_16160, n_16173);
  and g35154 (n19098, n19096, n19097);
  not g35155 (n_16441, n19096);
  not g35156 (n_16442, n19097);
  and g35157 (n19099, n_16441, n_16442);
  not g35158 (n_16443, n19098);
  not g35159 (n_16444, n19099);
  and g35160 (n19100, n_16443, n_16444);
  and g35161 (n19101, \b[21] , n11531);
  and g35162 (n19102, \b[19] , n11896);
  and g35163 (n19103, \b[20] , n11526);
  and g35169 (n19106, n1984, n11534);
  not g35172 (n_16449, n19107);
  and g35173 (n19108, \a[59] , n_16449);
  not g35174 (n_16450, n19108);
  and g35175 (n19109, \a[59] , n_16450);
  and g35176 (n19110, n_16449, n_16450);
  not g35177 (n_16451, n19109);
  not g35178 (n_16452, n19110);
  and g35179 (n19111, n_16451, n_16452);
  not g35180 (n_16453, n19111);
  and g35181 (n19112, n19100, n_16453);
  not g35182 (n_16454, n19112);
  and g35183 (n19113, n19100, n_16454);
  and g35184 (n19114, n_16453, n_16454);
  not g35185 (n_16455, n19113);
  not g35186 (n_16456, n19114);
  and g35187 (n19115, n_16455, n_16456);
  and g35188 (n19116, n_16177, n_16188);
  and g35189 (n19117, n19115, n19116);
  not g35190 (n_16457, n19115);
  not g35191 (n_16458, n19116);
  and g35192 (n19118, n_16457, n_16458);
  not g35193 (n_16459, n19117);
  not g35194 (n_16460, n19118);
  and g35195 (n19119, n_16459, n_16460);
  and g35196 (n19120, \b[24] , n10426);
  and g35197 (n19121, \b[22] , n10796);
  and g35198 (n19122, \b[23] , n10421);
  and g35204 (n19125, n2458, n10429);
  not g35207 (n_16465, n19126);
  and g35208 (n19127, \a[56] , n_16465);
  not g35209 (n_16466, n19127);
  and g35210 (n19128, \a[56] , n_16466);
  and g35211 (n19129, n_16465, n_16466);
  not g35212 (n_16467, n19128);
  not g35213 (n_16468, n19129);
  and g35214 (n19130, n_16467, n_16468);
  not g35215 (n_16469, n19130);
  and g35216 (n19131, n19119, n_16469);
  not g35217 (n_16470, n19119);
  and g35218 (n19132, n_16470, n19130);
  not g35219 (n_16471, n19070);
  not g35220 (n_16472, n19132);
  and g35221 (n19133, n_16471, n_16472);
  not g35222 (n_16473, n19131);
  and g35223 (n19134, n_16473, n19133);
  not g35224 (n_16474, n19134);
  and g35225 (n19135, n_16471, n_16474);
  and g35226 (n19136, n_16473, n_16474);
  and g35227 (n19137, n_16472, n19136);
  not g35228 (n_16475, n19135);
  not g35229 (n_16476, n19137);
  and g35230 (n19138, n_16475, n_16476);
  and g35231 (n19139, \b[27] , n9339);
  and g35232 (n19140, \b[25] , n9732);
  and g35233 (n19141, \b[26] , n9334);
  and g35239 (n19144, n2990, n9342);
  not g35242 (n_16481, n19145);
  and g35243 (n19146, \a[53] , n_16481);
  not g35244 (n_16482, n19146);
  and g35245 (n19147, \a[53] , n_16482);
  and g35246 (n19148, n_16481, n_16482);
  not g35247 (n_16483, n19147);
  not g35248 (n_16484, n19148);
  and g35249 (n19149, n_16483, n_16484);
  not g35250 (n_16485, n19138);
  not g35251 (n_16486, n19149);
  and g35252 (n19150, n_16485, n_16486);
  not g35253 (n_16487, n19150);
  and g35254 (n19151, n_16485, n_16487);
  and g35255 (n19152, n_16486, n_16487);
  not g35256 (n_16488, n19151);
  not g35257 (n_16489, n19152);
  and g35258 (n19153, n_16488, n_16489);
  and g35259 (n19154, n_16209, n_16213);
  and g35260 (n19155, n19153, n19154);
  not g35261 (n_16490, n19153);
  not g35262 (n_16491, n19154);
  and g35263 (n19156, n_16490, n_16491);
  not g35264 (n_16492, n19155);
  not g35265 (n_16493, n19156);
  and g35266 (n19157, n_16492, n_16493);
  and g35267 (n19158, \b[30] , n8362);
  and g35268 (n19159, \b[28] , n8715);
  and g35269 (n19160, \b[29] , n8357);
  and g35275 (n19163, n3577, n8365);
  not g35278 (n_16498, n19164);
  and g35279 (n19165, \a[50] , n_16498);
  not g35280 (n_16499, n19165);
  and g35281 (n19166, \a[50] , n_16499);
  and g35282 (n19167, n_16498, n_16499);
  not g35283 (n_16500, n19166);
  not g35284 (n_16501, n19167);
  and g35285 (n19168, n_16500, n_16501);
  not g35286 (n_16502, n19168);
  and g35287 (n19169, n19157, n_16502);
  not g35288 (n_16503, n19169);
  and g35289 (n19170, n19157, n_16503);
  and g35290 (n19171, n_16502, n_16503);
  not g35291 (n_16504, n19170);
  not g35292 (n_16505, n19171);
  and g35293 (n19172, n_16504, n_16505);
  and g35294 (n19173, n_16217, n_16228);
  and g35295 (n19174, n19172, n19173);
  not g35296 (n_16506, n19172);
  not g35297 (n_16507, n19173);
  and g35298 (n19175, n_16506, n_16507);
  not g35299 (n_16508, n19174);
  not g35300 (n_16509, n19175);
  and g35301 (n19176, n_16508, n_16509);
  and g35302 (n19177, \b[33] , n7446);
  and g35303 (n19178, \b[31] , n7787);
  and g35304 (n19179, \b[32] , n7441);
  and g35310 (n19182, n4223, n7449);
  not g35313 (n_16514, n19183);
  and g35314 (n19184, \a[47] , n_16514);
  not g35315 (n_16515, n19184);
  and g35316 (n19185, \a[47] , n_16515);
  and g35317 (n19186, n_16514, n_16515);
  not g35318 (n_16516, n19185);
  not g35319 (n_16517, n19186);
  and g35320 (n19187, n_16516, n_16517);
  not g35321 (n_16518, n19187);
  and g35322 (n19188, n19176, n_16518);
  not g35323 (n_16519, n19188);
  and g35324 (n19189, n19176, n_16519);
  and g35325 (n19190, n_16518, n_16519);
  not g35326 (n_16520, n19189);
  not g35327 (n_16521, n19190);
  and g35328 (n19191, n_16520, n_16521);
  not g35329 (n_16522, n19069);
  and g35330 (n19192, n_16522, n19191);
  not g35331 (n_16523, n19191);
  and g35332 (n19193, n19069, n_16523);
  not g35333 (n_16524, n19192);
  not g35334 (n_16525, n19193);
  and g35335 (n19194, n_16524, n_16525);
  and g35336 (n19195, \b[36] , n6595);
  and g35337 (n19196, \b[34] , n6902);
  and g35338 (n19197, \b[35] , n6590);
  and g35344 (n19200, n4922, n6598);
  not g35347 (n_16530, n19201);
  and g35348 (n19202, \a[44] , n_16530);
  not g35349 (n_16531, n19202);
  and g35350 (n19203, \a[44] , n_16531);
  and g35351 (n19204, n_16530, n_16531);
  not g35352 (n_16532, n19203);
  not g35353 (n_16533, n19204);
  and g35354 (n19205, n_16532, n_16533);
  not g35355 (n_16534, n19194);
  not g35356 (n_16535, n19205);
  and g35357 (n19206, n_16534, n_16535);
  and g35358 (n19207, n19194, n19205);
  not g35359 (n_16536, n19206);
  not g35360 (n_16537, n19207);
  and g35361 (n19208, n_16536, n_16537);
  not g35362 (n_16538, n19208);
  and g35363 (n19209, n19067, n_16538);
  not g35364 (n_16539, n19067);
  and g35365 (n19210, n_16539, n19208);
  not g35366 (n_16540, n19209);
  not g35367 (n_16541, n19210);
  and g35368 (n19211, n_16540, n_16541);
  and g35369 (n19212, \b[39] , n5777);
  and g35370 (n19213, \b[37] , n6059);
  and g35371 (n19214, \b[38] , n5772);
  and g35377 (n19217, n5451, n5780);
  not g35380 (n_16546, n19218);
  and g35381 (n19219, \a[41] , n_16546);
  not g35382 (n_16547, n19219);
  and g35383 (n19220, \a[41] , n_16547);
  and g35384 (n19221, n_16546, n_16547);
  not g35385 (n_16548, n19220);
  not g35386 (n_16549, n19221);
  and g35387 (n19222, n_16548, n_16549);
  not g35388 (n_16550, n19222);
  and g35389 (n19223, n19211, n_16550);
  not g35390 (n_16551, n19223);
  and g35391 (n19224, n19211, n_16551);
  and g35392 (n19225, n_16550, n_16551);
  not g35393 (n_16552, n19224);
  not g35394 (n_16553, n19225);
  and g35395 (n19226, n_16552, n_16553);
  not g35396 (n_16554, n19066);
  and g35397 (n19227, n_16554, n19226);
  not g35398 (n_16555, n19226);
  and g35399 (n19228, n19066, n_16555);
  not g35400 (n_16556, n19227);
  not g35401 (n_16557, n19228);
  and g35402 (n19229, n_16556, n_16557);
  and g35403 (n19230, \b[42] , n5035);
  and g35404 (n19231, \b[40] , n5277);
  and g35405 (n19232, \b[41] , n5030);
  and g35411 (n19235, n5038, n6489);
  not g35414 (n_16562, n19236);
  and g35415 (n19237, \a[38] , n_16562);
  not g35416 (n_16563, n19237);
  and g35417 (n19238, \a[38] , n_16563);
  and g35418 (n19239, n_16562, n_16563);
  not g35419 (n_16564, n19238);
  not g35420 (n_16565, n19239);
  and g35421 (n19240, n_16564, n_16565);
  not g35422 (n_16566, n19229);
  not g35423 (n_16567, n19240);
  and g35424 (n19241, n_16566, n_16567);
  and g35425 (n19242, n19229, n19240);
  not g35426 (n_16568, n19241);
  not g35427 (n_16569, n19242);
  and g35428 (n19243, n_16568, n_16569);
  not g35429 (n_16570, n19243);
  and g35430 (n19244, n19065, n_16570);
  not g35431 (n_16571, n19065);
  and g35432 (n19245, n_16571, n19243);
  not g35433 (n_16572, n19244);
  not g35434 (n_16573, n19245);
  and g35435 (n19246, n_16572, n_16573);
  and g35436 (n19247, \b[45] , n4287);
  and g35437 (n19248, \b[43] , n4532);
  and g35438 (n19249, \b[44] , n4282);
  and g35444 (n19252, n4290, n7361);
  not g35447 (n_16578, n19253);
  and g35448 (n19254, \a[35] , n_16578);
  not g35449 (n_16579, n19254);
  and g35450 (n19255, \a[35] , n_16579);
  and g35451 (n19256, n_16578, n_16579);
  not g35452 (n_16580, n19255);
  not g35453 (n_16581, n19256);
  and g35454 (n19257, n_16580, n_16581);
  not g35455 (n_16582, n19257);
  and g35456 (n19258, n19246, n_16582);
  not g35457 (n_16583, n19258);
  and g35458 (n19259, n19246, n_16583);
  and g35459 (n19260, n_16582, n_16583);
  not g35460 (n_16584, n19259);
  not g35461 (n_16585, n19260);
  and g35462 (n19261, n_16584, n_16585);
  and g35463 (n19262, n_16290, n_16293);
  and g35464 (n19263, n19261, n19262);
  not g35465 (n_16586, n19261);
  not g35466 (n_16587, n19262);
  and g35467 (n19264, n_16586, n_16587);
  not g35468 (n_16588, n19263);
  not g35469 (n_16589, n19264);
  and g35470 (n19265, n_16588, n_16589);
  and g35471 (n19266, n_16129, n_16297);
  and g35472 (n19267, \b[48] , n3638);
  and g35473 (n19268, \b[46] , n3843);
  and g35474 (n19269, \b[47] , n3633);
  and g35480 (n19272, n3641, n8009);
  not g35483 (n_16594, n19273);
  and g35484 (n19274, \a[32] , n_16594);
  not g35485 (n_16595, n19274);
  and g35486 (n19275, \a[32] , n_16595);
  and g35487 (n19276, n_16594, n_16595);
  not g35488 (n_16596, n19275);
  not g35489 (n_16597, n19276);
  and g35490 (n19277, n_16596, n_16597);
  not g35491 (n_16598, n19266);
  not g35492 (n_16599, n19277);
  and g35493 (n19278, n_16598, n_16599);
  not g35494 (n_16600, n19278);
  and g35495 (n19279, n_16598, n_16600);
  and g35496 (n19280, n_16599, n_16600);
  not g35497 (n_16601, n19279);
  not g35498 (n_16602, n19280);
  and g35499 (n19281, n_16601, n_16602);
  not g35500 (n_16603, n19281);
  and g35501 (n19282, n19265, n_16603);
  not g35502 (n_16604, n19265);
  and g35503 (n19283, n_16604, n19281);
  not g35504 (n_16605, n19283);
  and g35505 (n19284, n19064, n_16605);
  not g35506 (n_16606, n19282);
  and g35507 (n19285, n_16606, n19284);
  not g35508 (n_16607, n19285);
  and g35509 (n19286, n19064, n_16607);
  and g35510 (n19287, n_16605, n_16607);
  and g35511 (n19288, n_16606, n19287);
  not g35512 (n_16608, n19286);
  not g35513 (n_16609, n19288);
  and g35514 (n19289, n_16608, n_16609);
  not g35515 (n_16610, n19289);
  and g35516 (n19290, n19049, n_16610);
  not g35517 (n_16611, n19049);
  and g35518 (n19291, n_16611, n19289);
  not g35519 (n_16612, n19034);
  not g35520 (n_16613, n19291);
  and g35521 (n19292, n_16612, n_16613);
  not g35522 (n_16614, n19290);
  and g35523 (n19293, n_16614, n19292);
  not g35524 (n_16615, n19293);
  and g35525 (n19294, n_16612, n_16615);
  and g35526 (n19295, n_16613, n_16615);
  and g35527 (n19296, n_16614, n19295);
  not g35528 (n_16616, n19294);
  not g35529 (n_16617, n19296);
  and g35530 (n19297, n_16616, n_16617);
  not g35531 (n_16618, n19297);
  and g35532 (n19298, n19019, n_16618);
  not g35533 (n_16619, n19019);
  and g35534 (n19299, n_16619, n19297);
  not g35535 (n_16620, n19004);
  not g35536 (n_16621, n19299);
  and g35537 (n19300, n_16620, n_16621);
  not g35538 (n_16622, n19298);
  and g35539 (n19301, n_16622, n19300);
  not g35540 (n_16623, n19301);
  and g35541 (n19302, n_16620, n_16623);
  and g35542 (n19303, n_16621, n_16623);
  and g35543 (n19304, n_16622, n19303);
  not g35544 (n_16624, n19302);
  not g35545 (n_16625, n19304);
  and g35546 (n19305, n_16624, n_16625);
  and g35547 (n19306, n_16079, n_16346);
  and g35548 (n19307, n19305, n19306);
  not g35549 (n_16626, n19305);
  not g35550 (n_16627, n19306);
  and g35551 (n19308, n_16626, n_16627);
  not g35552 (n_16628, n19307);
  not g35553 (n_16629, n19308);
  and g35554 (n19309, n_16628, n_16629);
  and g35555 (n19310, n_16350, n_16354);
  not g35556 (n_16630, n19310);
  and g35557 (n19311, n19309, n_16630);
  not g35558 (n_16631, n19309);
  and g35559 (n19312, n_16631, n19310);
  not g35560 (n_16632, n19311);
  not g35561 (n_16633, n19312);
  and g35562 (\f[78] , n_16632, n_16633);
  and g35563 (n19314, n_16380, n_16622);
  and g35564 (n19315, \b[62] , n1391);
  and g35565 (n19316, \b[63] , n1297);
  not g35566 (n_16634, n19315);
  not g35567 (n_16635, n19316);
  and g35568 (n19317, n_16634, n_16635);
  and g35569 (n19318, n_13260, n19317);
  and g35570 (n19319, n13800, n19317);
  not g35571 (n_16636, n19318);
  not g35572 (n_16637, n19319);
  and g35573 (n19320, n_16636, n_16637);
  not g35574 (n_16638, n19320);
  and g35575 (n19321, \a[17] , n_16638);
  and g35576 (n19322, n_926, n19320);
  not g35577 (n_16639, n19321);
  not g35578 (n_16640, n19322);
  and g35579 (n19323, n_16639, n_16640);
  not g35580 (n_16641, n19314);
  not g35581 (n_16642, n19323);
  and g35582 (n19324, n_16641, n_16642);
  and g35583 (n19325, n19314, n19323);
  not g35584 (n_16643, n19324);
  not g35585 (n_16644, n19325);
  and g35586 (n19326, n_16643, n_16644);
  and g35587 (n19327, \b[61] , n1627);
  and g35588 (n19328, \b[59] , n1763);
  and g35589 (n19329, \b[60] , n1622);
  and g35595 (n19332, n1630, n12969);
  not g35598 (n_16649, n19333);
  and g35599 (n19334, \a[20] , n_16649);
  not g35600 (n_16650, n19334);
  and g35601 (n19335, \a[20] , n_16650);
  and g35602 (n19336, n_16649, n_16650);
  not g35603 (n_16651, n19335);
  not g35604 (n_16652, n19336);
  and g35605 (n19337, n_16651, n_16652);
  and g35606 (n19338, n_16389, n_16390);
  not g35607 (n_16653, n19338);
  and g35608 (n19339, n_16615, n_16653);
  and g35609 (n19340, n19337, n19339);
  not g35610 (n_16654, n19337);
  not g35611 (n_16655, n19339);
  and g35612 (n19341, n_16654, n_16655);
  not g35613 (n_16656, n19340);
  not g35614 (n_16657, n19341);
  and g35615 (n19342, n_16656, n_16657);
  and g35616 (n19343, n_16404, n_16614);
  and g35617 (n19344, \b[58] , n2048);
  and g35618 (n19345, \b[56] , n2198);
  and g35619 (n19346, \b[57] , n2043);
  not g35620 (n_16658, n19345);
  not g35621 (n_16659, n19346);
  and g35622 (n19347, n_16658, n_16659);
  not g35623 (n_16660, n19344);
  and g35624 (n19348, n_16660, n19347);
  and g35625 (n19349, n_15432, n19348);
  and g35626 (n19350, n_13160, n19348);
  not g35627 (n_16661, n19349);
  not g35628 (n_16662, n19350);
  and g35629 (n19351, n_16661, n_16662);
  not g35630 (n_16663, n19351);
  and g35631 (n19352, \a[23] , n_16663);
  and g35632 (n19353, n_1590, n19351);
  not g35633 (n_16664, n19352);
  not g35634 (n_16665, n19353);
  and g35635 (n19354, n_16664, n_16665);
  not g35636 (n_16666, n19343);
  not g35637 (n_16667, n19354);
  and g35638 (n19355, n_16666, n_16667);
  and g35639 (n19356, n19343, n19354);
  not g35640 (n_16668, n19355);
  not g35641 (n_16669, n19356);
  and g35642 (n19357, n_16668, n_16669);
  and g35643 (n19358, \b[55] , n2539);
  and g35644 (n19359, \b[53] , n2685);
  and g35645 (n19360, \b[54] , n2534);
  and g35651 (n19363, n2542, n10684);
  not g35654 (n_16674, n19364);
  and g35655 (n19365, \a[26] , n_16674);
  not g35656 (n_16675, n19365);
  and g35657 (n19366, \a[26] , n_16675);
  and g35658 (n19367, n_16674, n_16675);
  not g35659 (n_16676, n19366);
  not g35660 (n_16677, n19367);
  and g35661 (n19368, n_16676, n_16677);
  and g35662 (n19369, n_16416, n_16607);
  and g35663 (n19370, n19368, n19369);
  not g35664 (n_16678, n19368);
  not g35665 (n_16679, n19369);
  and g35666 (n19371, n_16678, n_16679);
  not g35667 (n_16680, n19370);
  not g35668 (n_16681, n19371);
  and g35669 (n19372, n_16680, n_16681);
  and g35670 (n19373, \b[52] , n3050);
  and g35671 (n19374, \b[50] , n3243);
  and g35672 (n19375, \b[51] , n3045);
  and g35678 (n19378, n3053, n9628);
  not g35681 (n_16686, n19379);
  and g35682 (n19380, \a[29] , n_16686);
  not g35683 (n_16687, n19380);
  and g35684 (n19381, \a[29] , n_16687);
  and g35685 (n19382, n_16686, n_16687);
  not g35686 (n_16688, n19381);
  not g35687 (n_16689, n19382);
  and g35688 (n19383, n_16688, n_16689);
  and g35689 (n19384, n_16600, n_16606);
  not g35690 (n_16690, n19383);
  not g35691 (n_16691, n19384);
  and g35692 (n19385, n_16690, n_16691);
  not g35693 (n_16692, n19385);
  and g35694 (n19386, n_16690, n_16692);
  and g35695 (n19387, n_16691, n_16692);
  not g35696 (n_16693, n19386);
  not g35697 (n_16694, n19387);
  and g35698 (n19388, n_16693, n_16694);
  and g35699 (n19389, \b[49] , n3638);
  and g35700 (n19390, \b[47] , n3843);
  and g35701 (n19391, \b[48] , n3633);
  and g35707 (n19394, n3641, n8625);
  not g35710 (n_16699, n19395);
  and g35711 (n19396, \a[32] , n_16699);
  not g35712 (n_16700, n19396);
  and g35713 (n19397, \a[32] , n_16700);
  and g35714 (n19398, n_16699, n_16700);
  not g35715 (n_16701, n19397);
  not g35716 (n_16702, n19398);
  and g35717 (n19399, n_16701, n_16702);
  and g35718 (n19400, n_16583, n_16589);
  and g35719 (n19401, n19399, n19400);
  not g35720 (n_16703, n19399);
  not g35721 (n_16704, n19400);
  and g35722 (n19402, n_16703, n_16704);
  not g35723 (n_16705, n19401);
  not g35724 (n_16706, n19402);
  and g35725 (n19403, n_16705, n_16706);
  and g35726 (n19404, \b[43] , n5035);
  and g35727 (n19405, \b[41] , n5277);
  and g35728 (n19406, \b[42] , n5030);
  and g35734 (n19409, n5038, n6515);
  not g35737 (n_16711, n19410);
  and g35738 (n19411, \a[38] , n_16711);
  not g35739 (n_16712, n19411);
  and g35740 (n19412, \a[38] , n_16712);
  and g35741 (n19413, n_16711, n_16712);
  not g35742 (n_16713, n19412);
  not g35743 (n_16714, n19413);
  and g35744 (n19414, n_16713, n_16714);
  and g35745 (n19415, n_16554, n_16555);
  not g35746 (n_16715, n19415);
  and g35747 (n19416, n_16551, n_16715);
  and g35748 (n19417, \b[40] , n5777);
  and g35749 (n19418, \b[38] , n6059);
  and g35750 (n19419, \b[39] , n5772);
  and g35756 (n19422, n5780, n5955);
  not g35759 (n_16720, n19423);
  and g35760 (n19424, \a[41] , n_16720);
  not g35761 (n_16721, n19424);
  and g35762 (n19425, \a[41] , n_16721);
  and g35763 (n19426, n_16720, n_16721);
  not g35764 (n_16722, n19425);
  not g35765 (n_16723, n19426);
  and g35766 (n19427, n_16722, n_16723);
  and g35767 (n19428, n_16536, n_16541);
  and g35768 (n19429, \b[37] , n6595);
  and g35769 (n19430, \b[35] , n6902);
  and g35770 (n19431, \b[36] , n6590);
  and g35776 (n19434, n5181, n6598);
  not g35779 (n_16728, n19435);
  and g35780 (n19436, \a[44] , n_16728);
  not g35781 (n_16729, n19436);
  and g35782 (n19437, \a[44] , n_16729);
  and g35783 (n19438, n_16728, n_16729);
  not g35784 (n_16730, n19437);
  not g35785 (n_16731, n19438);
  and g35786 (n19439, n_16730, n_16731);
  and g35787 (n19440, n_16522, n_16523);
  not g35788 (n_16732, n19440);
  and g35789 (n19441, n_16519, n_16732);
  and g35790 (n19442, \b[31] , n8362);
  and g35791 (n19443, \b[29] , n8715);
  and g35792 (n19444, \b[30] , n8357);
  and g35798 (n19447, n3796, n8365);
  not g35801 (n_16737, n19448);
  and g35802 (n19449, \a[50] , n_16737);
  not g35803 (n_16738, n19449);
  and g35804 (n19450, \a[50] , n_16738);
  and g35805 (n19451, n_16737, n_16738);
  not g35806 (n_16739, n19450);
  not g35807 (n_16740, n19451);
  and g35808 (n19452, n_16739, n_16740);
  and g35809 (n19453, n_16438, n_16444);
  and g35810 (n19454, \b[15] , n13903);
  and g35811 (n19455, \b[16] , n_11555);
  not g35812 (n_16741, n19454);
  not g35813 (n_16742, n19455);
  and g35814 (n19456, n_16741, n_16742);
  and g35815 (n19457, n_16421, n_16425);
  not g35816 (n_16743, n19456);
  and g35817 (n19458, n_16743, n19457);
  not g35818 (n_16744, n19457);
  and g35819 (n19459, n19456, n_16744);
  not g35820 (n_16745, n19458);
  not g35821 (n_16746, n19459);
  and g35822 (n19460, n_16745, n_16746);
  and g35823 (n19461, \b[19] , n12668);
  and g35824 (n19462, \b[17] , n13047);
  and g35825 (n19463, \b[18] , n12663);
  not g35826 (n_16747, n19462);
  not g35827 (n_16748, n19463);
  and g35828 (n19464, n_16747, n_16748);
  not g35829 (n_16749, n19461);
  and g35830 (n19465, n_16749, n19464);
  and g35831 (n19466, n_12644, n19465);
  not g35832 (n_16750, n1708);
  and g35833 (n19467, n_16750, n19465);
  not g35834 (n_16751, n19466);
  not g35835 (n_16752, n19467);
  and g35836 (n19468, n_16751, n_16752);
  not g35837 (n_16753, n19468);
  and g35838 (n19469, \a[62] , n_16753);
  and g35839 (n19470, n_10843, n19468);
  not g35840 (n_16754, n19469);
  not g35841 (n_16755, n19470);
  and g35842 (n19471, n_16754, n_16755);
  not g35843 (n_16756, n19471);
  and g35844 (n19472, n19460, n_16756);
  not g35845 (n_16757, n19460);
  and g35846 (n19473, n_16757, n19471);
  not g35847 (n_16758, n19472);
  not g35848 (n_16759, n19473);
  and g35849 (n19474, n_16758, n_16759);
  not g35850 (n_16760, n19453);
  and g35851 (n19475, n_16760, n19474);
  not g35852 (n_16761, n19474);
  and g35853 (n19476, n19453, n_16761);
  not g35854 (n_16762, n19475);
  not g35855 (n_16763, n19476);
  and g35856 (n19477, n_16762, n_16763);
  and g35857 (n19478, \b[22] , n11531);
  and g35858 (n19479, \b[20] , n11896);
  and g35859 (n19480, \b[21] , n11526);
  and g35865 (n19483, n2145, n11534);
  not g35868 (n_16768, n19484);
  and g35869 (n19485, \a[59] , n_16768);
  not g35870 (n_16769, n19485);
  and g35871 (n19486, \a[59] , n_16769);
  and g35872 (n19487, n_16768, n_16769);
  not g35873 (n_16770, n19486);
  not g35874 (n_16771, n19487);
  and g35875 (n19488, n_16770, n_16771);
  not g35876 (n_16772, n19488);
  and g35877 (n19489, n19477, n_16772);
  not g35878 (n_16773, n19489);
  and g35879 (n19490, n19477, n_16773);
  and g35880 (n19491, n_16772, n_16773);
  not g35881 (n_16774, n19490);
  not g35882 (n_16775, n19491);
  and g35883 (n19492, n_16774, n_16775);
  and g35884 (n19493, n_16454, n_16460);
  and g35885 (n19494, n19492, n19493);
  not g35886 (n_16776, n19492);
  not g35887 (n_16777, n19493);
  and g35888 (n19495, n_16776, n_16777);
  not g35889 (n_16778, n19494);
  not g35890 (n_16779, n19495);
  and g35891 (n19496, n_16778, n_16779);
  and g35892 (n19497, \b[25] , n10426);
  and g35893 (n19498, \b[23] , n10796);
  and g35894 (n19499, \b[24] , n10421);
  and g35900 (n19502, n2485, n10429);
  not g35903 (n_16784, n19503);
  and g35904 (n19504, \a[56] , n_16784);
  not g35905 (n_16785, n19504);
  and g35906 (n19505, \a[56] , n_16785);
  and g35907 (n19506, n_16784, n_16785);
  not g35908 (n_16786, n19505);
  not g35909 (n_16787, n19506);
  and g35910 (n19507, n_16786, n_16787);
  not g35911 (n_16788, n19507);
  and g35912 (n19508, n19496, n_16788);
  not g35913 (n_16789, n19508);
  and g35914 (n19509, n19496, n_16789);
  and g35915 (n19510, n_16788, n_16789);
  not g35916 (n_16790, n19509);
  not g35917 (n_16791, n19510);
  and g35918 (n19511, n_16790, n_16791);
  not g35919 (n_16792, n19136);
  and g35920 (n19512, n_16792, n19511);
  not g35921 (n_16793, n19511);
  and g35922 (n19513, n19136, n_16793);
  not g35923 (n_16794, n19512);
  not g35924 (n_16795, n19513);
  and g35925 (n19514, n_16794, n_16795);
  and g35926 (n19515, \b[28] , n9339);
  and g35927 (n19516, \b[26] , n9732);
  and g35928 (n19517, \b[27] , n9334);
  and g35934 (n19520, n3189, n9342);
  not g35937 (n_16800, n19521);
  and g35938 (n19522, \a[53] , n_16800);
  not g35939 (n_16801, n19522);
  and g35940 (n19523, \a[53] , n_16801);
  and g35941 (n19524, n_16800, n_16801);
  not g35942 (n_16802, n19523);
  not g35943 (n_16803, n19524);
  and g35944 (n19525, n_16802, n_16803);
  and g35945 (n19526, n19514, n19525);
  not g35946 (n_16804, n19514);
  not g35947 (n_16805, n19525);
  and g35948 (n19527, n_16804, n_16805);
  not g35949 (n_16806, n19526);
  not g35950 (n_16807, n19527);
  and g35951 (n19528, n_16806, n_16807);
  and g35952 (n19529, n_16487, n_16493);
  not g35953 (n_16808, n19529);
  and g35954 (n19530, n19528, n_16808);
  not g35955 (n_16809, n19528);
  and g35956 (n19531, n_16809, n19529);
  not g35957 (n_16810, n19530);
  not g35958 (n_16811, n19531);
  and g35959 (n19532, n_16810, n_16811);
  not g35960 (n_16812, n19452);
  and g35961 (n19533, n_16812, n19532);
  not g35962 (n_16813, n19533);
  and g35963 (n19534, n19532, n_16813);
  and g35964 (n19535, n_16812, n_16813);
  not g35965 (n_16814, n19534);
  not g35966 (n_16815, n19535);
  and g35967 (n19536, n_16814, n_16815);
  and g35968 (n19537, n_16503, n_16509);
  and g35969 (n19538, n19536, n19537);
  not g35970 (n_16816, n19536);
  not g35971 (n_16817, n19537);
  and g35972 (n19539, n_16816, n_16817);
  not g35973 (n_16818, n19538);
  not g35974 (n_16819, n19539);
  and g35975 (n19540, n_16818, n_16819);
  and g35976 (n19541, \b[34] , n7446);
  and g35977 (n19542, \b[32] , n7787);
  and g35978 (n19543, \b[33] , n7441);
  and g35984 (n19546, n4466, n7449);
  not g35987 (n_16824, n19547);
  and g35988 (n19548, \a[47] , n_16824);
  not g35989 (n_16825, n19548);
  and g35990 (n19549, \a[47] , n_16825);
  and g35991 (n19550, n_16824, n_16825);
  not g35992 (n_16826, n19549);
  not g35993 (n_16827, n19550);
  and g35994 (n19551, n_16826, n_16827);
  not g35995 (n_16828, n19540);
  and g35996 (n19552, n_16828, n19551);
  not g35997 (n_16829, n19551);
  and g35998 (n19553, n19540, n_16829);
  not g35999 (n_16830, n19552);
  not g36000 (n_16831, n19553);
  and g36001 (n19554, n_16830, n_16831);
  not g36002 (n_16832, n19441);
  and g36003 (n19555, n_16832, n19554);
  not g36004 (n_16833, n19555);
  and g36005 (n19556, n_16832, n_16833);
  and g36006 (n19557, n19554, n_16833);
  not g36007 (n_16834, n19556);
  not g36008 (n_16835, n19557);
  and g36009 (n19558, n_16834, n_16835);
  not g36010 (n_16836, n19439);
  not g36011 (n_16837, n19558);
  and g36012 (n19559, n_16836, n_16837);
  and g36013 (n19560, n19439, n_16835);
  and g36014 (n19561, n_16834, n19560);
  not g36015 (n_16838, n19559);
  not g36016 (n_16839, n19561);
  and g36017 (n19562, n_16838, n_16839);
  not g36018 (n_16840, n19428);
  and g36019 (n19563, n_16840, n19562);
  not g36020 (n_16841, n19563);
  and g36021 (n19564, n_16840, n_16841);
  and g36022 (n19565, n19562, n_16841);
  not g36023 (n_16842, n19564);
  not g36024 (n_16843, n19565);
  and g36025 (n19566, n_16842, n_16843);
  not g36026 (n_16844, n19427);
  not g36027 (n_16845, n19566);
  and g36028 (n19567, n_16844, n_16845);
  and g36029 (n19568, n19427, n_16843);
  and g36030 (n19569, n_16842, n19568);
  not g36031 (n_16846, n19567);
  not g36032 (n_16847, n19569);
  and g36033 (n19570, n_16846, n_16847);
  not g36034 (n_16848, n19416);
  and g36035 (n19571, n_16848, n19570);
  not g36036 (n_16849, n19570);
  and g36037 (n19572, n19416, n_16849);
  not g36038 (n_16850, n19571);
  not g36039 (n_16851, n19572);
  and g36040 (n19573, n_16850, n_16851);
  not g36041 (n_16852, n19414);
  and g36042 (n19574, n_16852, n19573);
  not g36043 (n_16853, n19574);
  and g36044 (n19575, n19573, n_16853);
  and g36045 (n19576, n_16852, n_16853);
  not g36046 (n_16854, n19575);
  not g36047 (n_16855, n19576);
  and g36048 (n19577, n_16854, n_16855);
  and g36049 (n19578, n_16568, n_16573);
  and g36050 (n19579, n19577, n19578);
  not g36051 (n_16856, n19577);
  not g36052 (n_16857, n19578);
  and g36053 (n19580, n_16856, n_16857);
  not g36054 (n_16858, n19579);
  not g36055 (n_16859, n19580);
  and g36056 (n19581, n_16858, n_16859);
  and g36057 (n19582, \b[46] , n4287);
  and g36058 (n19583, \b[44] , n4532);
  and g36059 (n19584, \b[45] , n4282);
  and g36065 (n19587, n4290, n7677);
  not g36068 (n_16864, n19588);
  and g36069 (n19589, \a[35] , n_16864);
  not g36070 (n_16865, n19589);
  and g36071 (n19590, \a[35] , n_16865);
  and g36072 (n19591, n_16864, n_16865);
  not g36073 (n_16866, n19590);
  not g36074 (n_16867, n19591);
  and g36075 (n19592, n_16866, n_16867);
  not g36076 (n_16868, n19592);
  and g36077 (n19593, n19581, n_16868);
  not g36078 (n_16869, n19593);
  and g36079 (n19594, n19581, n_16869);
  and g36080 (n19595, n_16868, n_16869);
  not g36081 (n_16870, n19594);
  not g36082 (n_16871, n19595);
  and g36083 (n19596, n_16870, n_16871);
  not g36084 (n_16872, n19596);
  and g36085 (n19597, n19403, n_16872);
  not g36086 (n_16873, n19403);
  and g36087 (n19598, n_16873, n19596);
  not g36088 (n_16874, n19388);
  not g36089 (n_16875, n19598);
  and g36090 (n19599, n_16874, n_16875);
  not g36091 (n_16876, n19597);
  and g36092 (n19600, n_16876, n19599);
  not g36093 (n_16877, n19600);
  and g36094 (n19601, n_16874, n_16877);
  and g36095 (n19602, n_16875, n_16877);
  and g36096 (n19603, n_16876, n19602);
  not g36097 (n_16878, n19601);
  not g36098 (n_16879, n19603);
  and g36099 (n19604, n_16878, n_16879);
  not g36100 (n_16880, n19604);
  and g36101 (n19605, n19372, n_16880);
  not g36102 (n_16881, n19372);
  and g36103 (n19606, n_16881, n19604);
  not g36104 (n_16882, n19606);
  and g36105 (n19607, n19357, n_16882);
  not g36106 (n_16883, n19605);
  and g36107 (n19608, n_16883, n19607);
  not g36108 (n_16884, n19608);
  and g36109 (n19609, n19357, n_16884);
  and g36110 (n19610, n_16882, n_16884);
  and g36111 (n19611, n_16883, n19610);
  not g36112 (n_16885, n19609);
  not g36113 (n_16886, n19611);
  and g36114 (n19612, n_16885, n_16886);
  not g36115 (n_16887, n19612);
  and g36116 (n19613, n19342, n_16887);
  not g36117 (n_16888, n19342);
  and g36118 (n19614, n_16888, n19612);
  not g36119 (n_16889, n19614);
  and g36120 (n19615, n19326, n_16889);
  not g36121 (n_16890, n19613);
  and g36122 (n19616, n_16890, n19615);
  not g36123 (n_16891, n19616);
  and g36124 (n19617, n19326, n_16891);
  and g36125 (n19618, n_16889, n_16891);
  and g36126 (n19619, n_16890, n19618);
  not g36127 (n_16892, n19617);
  not g36128 (n_16893, n19619);
  and g36129 (n19620, n_16892, n_16893);
  and g36130 (n19621, n_16366, n_16623);
  and g36131 (n19622, n19620, n19621);
  not g36132 (n_16894, n19620);
  not g36133 (n_16895, n19621);
  and g36134 (n19623, n_16894, n_16895);
  not g36135 (n_16896, n19622);
  not g36136 (n_16897, n19623);
  and g36137 (n19624, n_16896, n_16897);
  and g36138 (n19625, n_16629, n_16632);
  not g36139 (n_16898, n19625);
  and g36140 (n19626, n19624, n_16898);
  not g36141 (n_16899, n19624);
  and g36142 (n19627, n_16899, n19625);
  not g36143 (n_16900, n19626);
  not g36144 (n_16901, n19627);
  and g36145 (\f[79] , n_16900, n_16901);
  and g36146 (n19629, n_16897, n_16900);
  and g36147 (n19630, n_16643, n_16891);
  and g36148 (n19631, n_16657, n_16890);
  and g36149 (n19632, \b[63] , n1391);
  and g36150 (n19633, n1305, n13797);
  not g36151 (n_16902, n19632);
  not g36152 (n_16903, n19633);
  and g36153 (n19634, n_16902, n_16903);
  not g36154 (n_16904, n19634);
  and g36155 (n19635, \a[17] , n_16904);
  not g36156 (n_16905, n19635);
  and g36157 (n19636, \a[17] , n_16905);
  and g36158 (n19637, n_16904, n_16905);
  not g36159 (n_16906, n19636);
  not g36160 (n_16907, n19637);
  and g36161 (n19638, n_16906, n_16907);
  not g36162 (n_16908, n19631);
  not g36163 (n_16909, n19638);
  and g36164 (n19639, n_16908, n_16909);
  not g36165 (n_16910, n19639);
  and g36166 (n19640, n_16908, n_16910);
  and g36167 (n19641, n_16909, n_16910);
  not g36168 (n_16911, n19640);
  not g36169 (n_16912, n19641);
  and g36170 (n19642, n_16911, n_16912);
  and g36171 (n19643, \b[62] , n1627);
  and g36172 (n19644, \b[60] , n1763);
  and g36173 (n19645, \b[61] , n1622);
  and g36179 (n19648, n1630, n13370);
  not g36182 (n_16917, n19649);
  and g36183 (n19650, \a[20] , n_16917);
  not g36184 (n_16918, n19650);
  and g36185 (n19651, \a[20] , n_16918);
  and g36186 (n19652, n_16917, n_16918);
  not g36187 (n_16919, n19651);
  not g36188 (n_16920, n19652);
  and g36189 (n19653, n_16919, n_16920);
  and g36190 (n19654, n_16668, n_16884);
  and g36191 (n19655, n19653, n19654);
  not g36192 (n_16921, n19653);
  not g36193 (n_16922, n19654);
  and g36194 (n19656, n_16921, n_16922);
  not g36195 (n_16923, n19655);
  not g36196 (n_16924, n19656);
  and g36197 (n19657, n_16923, n_16924);
  and g36198 (n19658, \b[59] , n2048);
  and g36199 (n19659, \b[57] , n2198);
  and g36200 (n19660, \b[58] , n2043);
  and g36206 (n19663, n2051, n12179);
  not g36209 (n_16929, n19664);
  and g36210 (n19665, \a[23] , n_16929);
  not g36211 (n_16930, n19665);
  and g36212 (n19666, \a[23] , n_16930);
  and g36213 (n19667, n_16929, n_16930);
  not g36214 (n_16931, n19666);
  not g36215 (n_16932, n19667);
  and g36216 (n19668, n_16931, n_16932);
  and g36217 (n19669, n_16681, n_16883);
  not g36218 (n_16933, n19668);
  not g36219 (n_16934, n19669);
  and g36220 (n19670, n_16933, n_16934);
  not g36221 (n_16935, n19670);
  and g36222 (n19671, n_16933, n_16935);
  and g36223 (n19672, n_16934, n_16935);
  not g36224 (n_16936, n19671);
  not g36225 (n_16937, n19672);
  and g36226 (n19673, n_16936, n_16937);
  and g36227 (n19674, \b[56] , n2539);
  and g36228 (n19675, \b[54] , n2685);
  and g36229 (n19676, \b[55] , n2534);
  and g36235 (n19679, n2542, n10708);
  not g36238 (n_16942, n19680);
  and g36239 (n19681, \a[26] , n_16942);
  not g36240 (n_16943, n19681);
  and g36241 (n19682, \a[26] , n_16943);
  and g36242 (n19683, n_16942, n_16943);
  not g36243 (n_16944, n19682);
  not g36244 (n_16945, n19683);
  and g36245 (n19684, n_16944, n_16945);
  and g36246 (n19685, n_16692, n_16877);
  and g36247 (n19686, n19684, n19685);
  not g36248 (n_16946, n19684);
  not g36249 (n_16947, n19685);
  and g36250 (n19687, n_16946, n_16947);
  not g36251 (n_16948, n19686);
  not g36252 (n_16949, n19687);
  and g36253 (n19688, n_16948, n_16949);
  and g36254 (n19689, \b[53] , n3050);
  and g36255 (n19690, \b[51] , n3243);
  and g36256 (n19691, \b[52] , n3045);
  and g36262 (n19694, n3053, n9972);
  not g36265 (n_16954, n19695);
  and g36266 (n19696, \a[29] , n_16954);
  not g36267 (n_16955, n19696);
  and g36268 (n19697, \a[29] , n_16955);
  and g36269 (n19698, n_16954, n_16955);
  not g36270 (n_16956, n19697);
  not g36271 (n_16957, n19698);
  and g36272 (n19699, n_16956, n_16957);
  and g36273 (n19700, n_16706, n_16876);
  not g36274 (n_16958, n19699);
  not g36275 (n_16959, n19700);
  and g36276 (n19701, n_16958, n_16959);
  not g36277 (n_16960, n19701);
  and g36278 (n19702, n_16958, n_16960);
  and g36279 (n19703, n_16959, n_16960);
  not g36280 (n_16961, n19702);
  not g36281 (n_16962, n19703);
  and g36282 (n19704, n_16961, n_16962);
  and g36283 (n19705, \b[50] , n3638);
  and g36284 (n19706, \b[48] , n3843);
  and g36285 (n19707, \b[49] , n3633);
  and g36291 (n19710, n3641, n8949);
  not g36294 (n_16967, n19711);
  and g36295 (n19712, \a[32] , n_16967);
  not g36296 (n_16968, n19712);
  and g36297 (n19713, \a[32] , n_16968);
  and g36298 (n19714, n_16967, n_16968);
  not g36299 (n_16969, n19713);
  not g36300 (n_16970, n19714);
  and g36301 (n19715, n_16969, n_16970);
  and g36302 (n19716, n_16859, n_16869);
  and g36303 (n19717, n19715, n19716);
  not g36304 (n_16971, n19715);
  not g36305 (n_16972, n19716);
  and g36306 (n19718, n_16971, n_16972);
  not g36307 (n_16973, n19717);
  not g36308 (n_16974, n19718);
  and g36309 (n19719, n_16973, n_16974);
  and g36310 (n19720, n_16850, n_16853);
  and g36311 (n19721, \b[44] , n5035);
  and g36312 (n19722, \b[42] , n5277);
  and g36313 (n19723, \b[43] , n5030);
  and g36319 (n19726, n5038, n7072);
  not g36322 (n_16979, n19727);
  and g36323 (n19728, \a[38] , n_16979);
  not g36324 (n_16980, n19728);
  and g36325 (n19729, \a[38] , n_16980);
  and g36326 (n19730, n_16979, n_16980);
  not g36327 (n_16981, n19729);
  not g36328 (n_16982, n19730);
  and g36329 (n19731, n_16981, n_16982);
  and g36330 (n19732, n_16841, n_16846);
  and g36331 (n19733, \b[41] , n5777);
  and g36332 (n19734, \b[39] , n6059);
  and g36333 (n19735, \b[40] , n5772);
  and g36339 (n19738, n5780, n6219);
  not g36342 (n_16987, n19739);
  and g36343 (n19740, \a[41] , n_16987);
  not g36344 (n_16988, n19740);
  and g36345 (n19741, \a[41] , n_16988);
  and g36346 (n19742, n_16987, n_16988);
  not g36347 (n_16989, n19741);
  not g36348 (n_16990, n19742);
  and g36349 (n19743, n_16989, n_16990);
  and g36350 (n19744, n_16833, n_16838);
  and g36351 (n19745, n_16779, n_16789);
  and g36352 (n19746, \b[26] , n10426);
  and g36353 (n19747, \b[24] , n10796);
  and g36354 (n19748, \b[25] , n10421);
  and g36360 (n19751, n2813, n10429);
  not g36363 (n_16995, n19752);
  and g36364 (n19753, \a[56] , n_16995);
  not g36365 (n_16996, n19753);
  and g36366 (n19754, \a[56] , n_16996);
  and g36367 (n19755, n_16995, n_16996);
  not g36368 (n_16997, n19754);
  not g36369 (n_16998, n19755);
  and g36370 (n19756, n_16997, n_16998);
  and g36371 (n19757, n_16762, n_16773);
  and g36372 (n19758, \b[20] , n12668);
  and g36373 (n19759, \b[18] , n13047);
  and g36374 (n19760, \b[19] , n12663);
  and g36380 (n19763, n1846, n12671);
  not g36383 (n_17003, n19764);
  and g36384 (n19765, \a[62] , n_17003);
  not g36385 (n_17004, n19765);
  and g36386 (n19766, \a[62] , n_17004);
  and g36387 (n19767, n_17003, n_17004);
  not g36388 (n_17005, n19766);
  not g36389 (n_17006, n19767);
  and g36390 (n19768, n_17005, n_17006);
  and g36391 (n19769, \b[16] , n13903);
  and g36392 (n19770, \b[17] , n_11555);
  not g36393 (n_17007, n19769);
  not g36394 (n_17008, n19770);
  and g36395 (n19771, n_17007, n_17008);
  not g36396 (n_17009, n19771);
  and g36397 (n19772, n19456, n_17009);
  and g36398 (n19773, n_16743, n19771);
  not g36399 (n_17010, n19768);
  not g36400 (n_17011, n19773);
  and g36401 (n19774, n_17010, n_17011);
  not g36402 (n_17012, n19772);
  and g36403 (n19775, n_17012, n19774);
  not g36404 (n_17013, n19775);
  and g36405 (n19776, n_17010, n_17013);
  and g36406 (n19777, n_17011, n_17013);
  and g36407 (n19778, n_17012, n19777);
  not g36408 (n_17014, n19776);
  not g36409 (n_17015, n19778);
  and g36410 (n19779, n_17014, n_17015);
  and g36411 (n19780, n_16746, n_16758);
  and g36412 (n19781, n19779, n19780);
  not g36413 (n_17016, n19779);
  not g36414 (n_17017, n19780);
  and g36415 (n19782, n_17016, n_17017);
  not g36416 (n_17018, n19781);
  not g36417 (n_17019, n19782);
  and g36418 (n19783, n_17018, n_17019);
  and g36419 (n19784, \b[23] , n11531);
  and g36420 (n19785, \b[21] , n11896);
  and g36421 (n19786, \b[22] , n11526);
  and g36427 (n19789, n2300, n11534);
  not g36430 (n_17024, n19790);
  and g36431 (n19791, \a[59] , n_17024);
  not g36432 (n_17025, n19791);
  and g36433 (n19792, \a[59] , n_17025);
  and g36434 (n19793, n_17024, n_17025);
  not g36435 (n_17026, n19792);
  not g36436 (n_17027, n19793);
  and g36437 (n19794, n_17026, n_17027);
  not g36438 (n_17028, n19783);
  and g36439 (n19795, n_17028, n19794);
  not g36440 (n_17029, n19794);
  and g36441 (n19796, n19783, n_17029);
  not g36442 (n_17030, n19795);
  not g36443 (n_17031, n19796);
  and g36444 (n19797, n_17030, n_17031);
  not g36445 (n_17032, n19757);
  and g36446 (n19798, n_17032, n19797);
  not g36447 (n_17033, n19797);
  and g36448 (n19799, n19757, n_17033);
  not g36449 (n_17034, n19798);
  not g36450 (n_17035, n19799);
  and g36451 (n19800, n_17034, n_17035);
  not g36452 (n_17036, n19756);
  and g36453 (n19801, n_17036, n19800);
  not g36454 (n_17037, n19800);
  and g36455 (n19802, n19756, n_17037);
  not g36456 (n_17038, n19801);
  not g36457 (n_17039, n19802);
  and g36458 (n19803, n_17038, n_17039);
  not g36459 (n_17040, n19745);
  and g36460 (n19804, n_17040, n19803);
  not g36461 (n_17041, n19803);
  and g36462 (n19805, n19745, n_17041);
  not g36463 (n_17042, n19804);
  not g36464 (n_17043, n19805);
  and g36465 (n19806, n_17042, n_17043);
  and g36466 (n19807, \b[29] , n9339);
  and g36467 (n19808, \b[27] , n9732);
  and g36468 (n19809, \b[28] , n9334);
  and g36474 (n19812, n3383, n9342);
  not g36477 (n_17048, n19813);
  and g36478 (n19814, \a[53] , n_17048);
  not g36479 (n_17049, n19814);
  and g36480 (n19815, \a[53] , n_17049);
  and g36481 (n19816, n_17048, n_17049);
  not g36482 (n_17050, n19815);
  not g36483 (n_17051, n19816);
  and g36484 (n19817, n_17050, n_17051);
  not g36485 (n_17052, n19817);
  and g36486 (n19818, n19806, n_17052);
  not g36487 (n_17053, n19818);
  and g36488 (n19819, n19806, n_17053);
  and g36489 (n19820, n_17052, n_17053);
  not g36490 (n_17054, n19819);
  not g36491 (n_17055, n19820);
  and g36492 (n19821, n_17054, n_17055);
  and g36493 (n19822, n_16792, n_16793);
  not g36494 (n_17056, n19822);
  and g36495 (n19823, n_16807, n_17056);
  not g36496 (n_17057, n19821);
  not g36497 (n_17058, n19823);
  and g36498 (n19824, n_17057, n_17058);
  not g36499 (n_17059, n19824);
  and g36500 (n19825, n_17057, n_17059);
  and g36501 (n19826, n_17058, n_17059);
  not g36502 (n_17060, n19825);
  not g36503 (n_17061, n19826);
  and g36504 (n19827, n_17060, n_17061);
  and g36505 (n19828, \b[32] , n8362);
  and g36506 (n19829, \b[30] , n8715);
  and g36507 (n19830, \b[31] , n8357);
  and g36513 (n19833, n4013, n8365);
  not g36516 (n_17066, n19834);
  and g36517 (n19835, \a[50] , n_17066);
  not g36518 (n_17067, n19835);
  and g36519 (n19836, \a[50] , n_17067);
  and g36520 (n19837, n_17066, n_17067);
  not g36521 (n_17068, n19836);
  not g36522 (n_17069, n19837);
  and g36523 (n19838, n_17068, n_17069);
  not g36524 (n_17070, n19827);
  and g36525 (n19839, n_17070, n19838);
  not g36526 (n_17071, n19838);
  and g36527 (n19840, n19827, n_17071);
  not g36528 (n_17072, n19839);
  not g36529 (n_17073, n19840);
  and g36530 (n19841, n_17072, n_17073);
  and g36531 (n19842, n_16810, n_16813);
  and g36532 (n19843, n19841, n19842);
  not g36533 (n_17074, n19841);
  not g36534 (n_17075, n19842);
  and g36535 (n19844, n_17074, n_17075);
  not g36536 (n_17076, n19843);
  not g36537 (n_17077, n19844);
  and g36538 (n19845, n_17076, n_17077);
  and g36539 (n19846, \b[35] , n7446);
  and g36540 (n19847, \b[33] , n7787);
  and g36541 (n19848, \b[34] , n7441);
  and g36547 (n19851, n4696, n7449);
  not g36550 (n_17082, n19852);
  and g36551 (n19853, \a[47] , n_17082);
  not g36552 (n_17083, n19853);
  and g36553 (n19854, \a[47] , n_17083);
  and g36554 (n19855, n_17082, n_17083);
  not g36555 (n_17084, n19854);
  not g36556 (n_17085, n19855);
  and g36557 (n19856, n_17084, n_17085);
  not g36558 (n_17086, n19856);
  and g36559 (n19857, n19845, n_17086);
  not g36560 (n_17087, n19857);
  and g36561 (n19858, n19845, n_17087);
  and g36562 (n19859, n_17086, n_17087);
  not g36563 (n_17088, n19858);
  not g36564 (n_17089, n19859);
  and g36565 (n19860, n_17088, n_17089);
  and g36566 (n19861, n_16819, n_16831);
  not g36567 (n_17090, n19860);
  not g36568 (n_17091, n19861);
  and g36569 (n19862, n_17090, n_17091);
  not g36570 (n_17092, n19862);
  and g36571 (n19863, n_17090, n_17092);
  and g36572 (n19864, n_17091, n_17092);
  not g36573 (n_17093, n19863);
  not g36574 (n_17094, n19864);
  and g36575 (n19865, n_17093, n_17094);
  and g36576 (n19866, \b[38] , n6595);
  and g36577 (n19867, \b[36] , n6902);
  and g36578 (n19868, \b[37] , n6590);
  and g36584 (n19871, n5205, n6598);
  not g36587 (n_17099, n19872);
  and g36588 (n19873, \a[44] , n_17099);
  not g36589 (n_17100, n19873);
  and g36590 (n19874, \a[44] , n_17100);
  and g36591 (n19875, n_17099, n_17100);
  not g36592 (n_17101, n19874);
  not g36593 (n_17102, n19875);
  and g36594 (n19876, n_17101, n_17102);
  not g36595 (n_17103, n19865);
  and g36596 (n19877, n_17103, n19876);
  not g36597 (n_17104, n19876);
  and g36598 (n19878, n19865, n_17104);
  not g36599 (n_17105, n19877);
  not g36600 (n_17106, n19878);
  and g36601 (n19879, n_17105, n_17106);
  not g36602 (n_17107, n19744);
  not g36603 (n_17108, n19879);
  and g36604 (n19880, n_17107, n_17108);
  and g36605 (n19881, n19744, n19879);
  not g36606 (n_17109, n19880);
  not g36607 (n_17110, n19881);
  and g36608 (n19882, n_17109, n_17110);
  not g36609 (n_17111, n19743);
  and g36610 (n19883, n_17111, n19882);
  not g36611 (n_17112, n19882);
  and g36612 (n19884, n19743, n_17112);
  not g36613 (n_17113, n19883);
  not g36614 (n_17114, n19884);
  and g36615 (n19885, n_17113, n_17114);
  not g36616 (n_17115, n19732);
  and g36617 (n19886, n_17115, n19885);
  not g36618 (n_17116, n19885);
  and g36619 (n19887, n19732, n_17116);
  not g36620 (n_17117, n19886);
  not g36621 (n_17118, n19887);
  and g36622 (n19888, n_17117, n_17118);
  not g36623 (n_17119, n19731);
  and g36624 (n19889, n_17119, n19888);
  not g36625 (n_17120, n19888);
  and g36626 (n19890, n19731, n_17120);
  not g36627 (n_17121, n19889);
  not g36628 (n_17122, n19890);
  and g36629 (n19891, n_17121, n_17122);
  not g36630 (n_17123, n19720);
  and g36631 (n19892, n_17123, n19891);
  not g36632 (n_17124, n19891);
  and g36633 (n19893, n19720, n_17124);
  not g36634 (n_17125, n19892);
  not g36635 (n_17126, n19893);
  and g36636 (n19894, n_17125, n_17126);
  and g36637 (n19895, \b[47] , n4287);
  and g36638 (n19896, \b[45] , n4532);
  and g36639 (n19897, \b[46] , n4282);
  and g36645 (n19900, n4290, n7703);
  not g36648 (n_17131, n19901);
  and g36649 (n19902, \a[35] , n_17131);
  not g36650 (n_17132, n19902);
  and g36651 (n19903, \a[35] , n_17132);
  and g36652 (n19904, n_17131, n_17132);
  not g36653 (n_17133, n19903);
  not g36654 (n_17134, n19904);
  and g36655 (n19905, n_17133, n_17134);
  not g36656 (n_17135, n19905);
  and g36657 (n19906, n19894, n_17135);
  not g36658 (n_17136, n19906);
  and g36659 (n19907, n19894, n_17136);
  and g36660 (n19908, n_17135, n_17136);
  not g36661 (n_17137, n19907);
  not g36662 (n_17138, n19908);
  and g36663 (n19909, n_17137, n_17138);
  not g36664 (n_17139, n19909);
  and g36665 (n19910, n19719, n_17139);
  not g36666 (n_17140, n19719);
  and g36667 (n19911, n_17140, n19909);
  not g36668 (n_17141, n19704);
  not g36669 (n_17142, n19911);
  and g36670 (n19912, n_17141, n_17142);
  not g36671 (n_17143, n19910);
  and g36672 (n19913, n_17143, n19912);
  not g36673 (n_17144, n19913);
  and g36674 (n19914, n_17141, n_17144);
  and g36675 (n19915, n_17142, n_17144);
  and g36676 (n19916, n_17143, n19915);
  not g36677 (n_17145, n19914);
  not g36678 (n_17146, n19916);
  and g36679 (n19917, n_17145, n_17146);
  not g36680 (n_17147, n19917);
  and g36681 (n19918, n19688, n_17147);
  not g36682 (n_17148, n19688);
  and g36683 (n19919, n_17148, n19917);
  not g36684 (n_17149, n19673);
  not g36685 (n_17150, n19919);
  and g36686 (n19920, n_17149, n_17150);
  not g36687 (n_17151, n19918);
  and g36688 (n19921, n_17151, n19920);
  not g36689 (n_17152, n19921);
  and g36690 (n19922, n_17149, n_17152);
  and g36691 (n19923, n_17150, n_17152);
  and g36692 (n19924, n_17151, n19923);
  not g36693 (n_17153, n19922);
  not g36694 (n_17154, n19924);
  and g36695 (n19925, n_17153, n_17154);
  not g36696 (n_17155, n19657);
  and g36697 (n19926, n_17155, n19925);
  not g36698 (n_17156, n19925);
  and g36699 (n19927, n19657, n_17156);
  not g36700 (n_17157, n19926);
  not g36701 (n_17158, n19927);
  and g36702 (n19928, n_17157, n_17158);
  not g36703 (n_17159, n19642);
  and g36704 (n19929, n_17159, n19928);
  not g36705 (n_17160, n19928);
  and g36706 (n19930, n19642, n_17160);
  not g36707 (n_17161, n19929);
  not g36708 (n_17162, n19930);
  and g36709 (n19931, n_17161, n_17162);
  not g36710 (n_17163, n19630);
  and g36711 (n19932, n_17163, n19931);
  not g36712 (n_17164, n19932);
  and g36713 (n19933, n_17163, n_17164);
  and g36714 (n19934, n19931, n_17164);
  not g36715 (n_17165, n19933);
  not g36716 (n_17166, n19934);
  and g36717 (n19935, n_17165, n_17166);
  not g36718 (n_17167, n19629);
  not g36719 (n_17168, n19935);
  and g36720 (n19936, n_17167, n_17168);
  and g36721 (n19937, n19629, n_17166);
  and g36722 (n19938, n_17165, n19937);
  not g36723 (n_17169, n19936);
  not g36724 (n_17170, n19938);
  and g36725 (\f[80] , n_17169, n_17170);
  and g36726 (n19940, n_17164, n_17169);
  and g36727 (n19941, n_16910, n_17161);
  and g36728 (n19942, n_16924, n_17158);
  and g36729 (n19943, \b[63] , n1627);
  and g36730 (n19944, \b[61] , n1763);
  and g36731 (n19945, \b[62] , n1622);
  and g36737 (n19948, n1630, n13771);
  not g36740 (n_17175, n19949);
  and g36741 (n19950, \a[20] , n_17175);
  not g36742 (n_17176, n19950);
  and g36743 (n19951, \a[20] , n_17176);
  and g36744 (n19952, n_17175, n_17176);
  not g36745 (n_17177, n19951);
  not g36746 (n_17178, n19952);
  and g36747 (n19953, n_17177, n_17178);
  not g36748 (n_17179, n19942);
  not g36749 (n_17180, n19953);
  and g36750 (n19954, n_17179, n_17180);
  not g36751 (n_17181, n19954);
  and g36752 (n19955, n_17179, n_17181);
  and g36753 (n19956, n_17180, n_17181);
  not g36754 (n_17182, n19955);
  not g36755 (n_17183, n19956);
  and g36756 (n19957, n_17182, n_17183);
  and g36757 (n19958, \b[60] , n2048);
  and g36758 (n19959, \b[58] , n2198);
  and g36759 (n19960, \b[59] , n2043);
  and g36765 (n19963, n2051, n12211);
  not g36768 (n_17188, n19964);
  and g36769 (n19965, \a[23] , n_17188);
  not g36770 (n_17189, n19965);
  and g36771 (n19966, \a[23] , n_17189);
  and g36772 (n19967, n_17188, n_17189);
  not g36773 (n_17190, n19966);
  not g36774 (n_17191, n19967);
  and g36775 (n19968, n_17190, n_17191);
  and g36776 (n19969, n_16935, n_17152);
  and g36777 (n19970, n19968, n19969);
  not g36778 (n_17192, n19968);
  not g36779 (n_17193, n19969);
  and g36780 (n19971, n_17192, n_17193);
  not g36781 (n_17194, n19970);
  not g36782 (n_17195, n19971);
  and g36783 (n19972, n_17194, n_17195);
  and g36784 (n19973, \b[54] , n3050);
  and g36785 (n19974, \b[52] , n3243);
  and g36786 (n19975, \b[53] , n3045);
  and g36792 (n19978, n3053, n9998);
  not g36795 (n_17200, n19979);
  and g36796 (n19980, \a[29] , n_17200);
  not g36797 (n_17201, n19980);
  and g36798 (n19981, \a[29] , n_17201);
  and g36799 (n19982, n_17200, n_17201);
  not g36800 (n_17202, n19981);
  not g36801 (n_17203, n19982);
  and g36802 (n19983, n_17202, n_17203);
  and g36803 (n19984, n_16960, n_17144);
  and g36804 (n19985, n19983, n19984);
  not g36805 (n_17204, n19983);
  not g36806 (n_17205, n19984);
  and g36807 (n19986, n_17204, n_17205);
  not g36808 (n_17206, n19985);
  not g36809 (n_17207, n19986);
  and g36810 (n19987, n_17206, n_17207);
  and g36811 (n19988, n_17109, n_17113);
  and g36812 (n19989, n_17103, n_17104);
  not g36813 (n_17208, n19989);
  and g36814 (n19990, n_17092, n_17208);
  and g36815 (n19991, n_17077, n_17087);
  and g36816 (n19992, \b[27] , n10426);
  and g36817 (n19993, \b[25] , n10796);
  and g36818 (n19994, \b[26] , n10421);
  and g36824 (n19997, n2990, n10429);
  not g36827 (n_17213, n19998);
  and g36828 (n19999, \a[56] , n_17213);
  not g36829 (n_17214, n19999);
  and g36830 (n20000, \a[56] , n_17214);
  and g36831 (n20001, n_17213, n_17214);
  not g36832 (n_17215, n20000);
  not g36833 (n_17216, n20001);
  and g36834 (n20002, n_17215, n_17216);
  and g36835 (n20003, n_17019, n_17031);
  and g36836 (n20004, \b[21] , n12668);
  and g36837 (n20005, \b[19] , n13047);
  and g36838 (n20006, \b[20] , n12663);
  and g36844 (n20009, n1984, n12671);
  not g36847 (n_17221, n20010);
  and g36848 (n20011, \a[62] , n_17221);
  not g36849 (n_17222, n20011);
  and g36850 (n20012, \a[62] , n_17222);
  and g36851 (n20013, n_17221, n_17222);
  not g36852 (n_17223, n20012);
  not g36853 (n_17224, n20013);
  and g36854 (n20014, n_17223, n_17224);
  and g36855 (n20015, \b[17] , n13903);
  and g36856 (n20016, \b[18] , n_11555);
  not g36857 (n_17225, n20015);
  not g36858 (n_17226, n20016);
  and g36859 (n20017, n_17225, n_17226);
  not g36860 (n_17227, n20017);
  and g36861 (n20018, n_926, n_17227);
  and g36862 (n20019, \a[17] , n20017);
  not g36863 (n_17228, n20018);
  not g36864 (n_17229, n20019);
  and g36865 (n20020, n_17228, n_17229);
  and g36866 (n20021, n_17009, n20020);
  not g36867 (n_17230, n20020);
  and g36868 (n20022, n19771, n_17230);
  not g36869 (n_17231, n20021);
  not g36870 (n_17232, n20022);
  and g36871 (n20023, n_17231, n_17232);
  not g36872 (n_17233, n20014);
  and g36873 (n20024, n_17233, n20023);
  not g36874 (n_17234, n20024);
  and g36875 (n20025, n_17233, n_17234);
  and g36876 (n20026, n20023, n_17234);
  not g36877 (n_17235, n20025);
  not g36878 (n_17236, n20026);
  and g36879 (n20027, n_17235, n_17236);
  not g36880 (n_17237, n19777);
  not g36881 (n_17238, n20027);
  and g36882 (n20028, n_17237, n_17238);
  not g36883 (n_17239, n20028);
  and g36884 (n20029, n_17237, n_17239);
  and g36885 (n20030, n_17238, n_17239);
  not g36886 (n_17240, n20029);
  not g36887 (n_17241, n20030);
  and g36888 (n20031, n_17240, n_17241);
  and g36889 (n20032, \b[24] , n11531);
  and g36890 (n20033, \b[22] , n11896);
  and g36891 (n20034, \b[23] , n11526);
  and g36897 (n20037, n2458, n11534);
  not g36900 (n_17246, n20038);
  and g36901 (n20039, \a[59] , n_17246);
  not g36902 (n_17247, n20039);
  and g36903 (n20040, \a[59] , n_17247);
  and g36904 (n20041, n_17246, n_17247);
  not g36905 (n_17248, n20040);
  not g36906 (n_17249, n20041);
  and g36907 (n20042, n_17248, n_17249);
  and g36908 (n20043, n20031, n20042);
  not g36909 (n_17250, n20031);
  not g36910 (n_17251, n20042);
  and g36911 (n20044, n_17250, n_17251);
  not g36912 (n_17252, n20043);
  not g36913 (n_17253, n20044);
  and g36914 (n20045, n_17252, n_17253);
  not g36915 (n_17254, n20003);
  and g36916 (n20046, n_17254, n20045);
  not g36917 (n_17255, n20045);
  and g36918 (n20047, n20003, n_17255);
  not g36919 (n_17256, n20046);
  not g36920 (n_17257, n20047);
  and g36921 (n20048, n_17256, n_17257);
  not g36922 (n_17258, n20002);
  and g36923 (n20049, n_17258, n20048);
  not g36924 (n_17259, n20049);
  and g36925 (n20050, n20048, n_17259);
  and g36926 (n20051, n_17258, n_17259);
  not g36927 (n_17260, n20050);
  not g36928 (n_17261, n20051);
  and g36929 (n20052, n_17260, n_17261);
  and g36930 (n20053, n_17034, n_17038);
  and g36931 (n20054, n20052, n20053);
  not g36932 (n_17262, n20052);
  not g36933 (n_17263, n20053);
  and g36934 (n20055, n_17262, n_17263);
  not g36935 (n_17264, n20054);
  not g36936 (n_17265, n20055);
  and g36937 (n20056, n_17264, n_17265);
  and g36938 (n20057, \b[30] , n9339);
  and g36939 (n20058, \b[28] , n9732);
  and g36940 (n20059, \b[29] , n9334);
  and g36946 (n20062, n3577, n9342);
  not g36949 (n_17270, n20063);
  and g36950 (n20064, \a[53] , n_17270);
  not g36951 (n_17271, n20064);
  and g36952 (n20065, \a[53] , n_17271);
  and g36953 (n20066, n_17270, n_17271);
  not g36954 (n_17272, n20065);
  not g36955 (n_17273, n20066);
  and g36956 (n20067, n_17272, n_17273);
  not g36957 (n_17274, n20067);
  and g36958 (n20068, n20056, n_17274);
  not g36959 (n_17275, n20068);
  and g36960 (n20069, n20056, n_17275);
  and g36961 (n20070, n_17274, n_17275);
  not g36962 (n_17276, n20069);
  not g36963 (n_17277, n20070);
  and g36964 (n20071, n_17276, n_17277);
  and g36965 (n20072, n_17042, n_17053);
  and g36966 (n20073, n20071, n20072);
  not g36967 (n_17278, n20071);
  not g36968 (n_17279, n20072);
  and g36969 (n20074, n_17278, n_17279);
  not g36970 (n_17280, n20073);
  not g36971 (n_17281, n20074);
  and g36972 (n20075, n_17280, n_17281);
  and g36973 (n20076, \b[33] , n8362);
  and g36974 (n20077, \b[31] , n8715);
  and g36975 (n20078, \b[32] , n8357);
  and g36981 (n20081, n4223, n8365);
  not g36984 (n_17286, n20082);
  and g36985 (n20083, \a[50] , n_17286);
  not g36986 (n_17287, n20083);
  and g36987 (n20084, \a[50] , n_17287);
  and g36988 (n20085, n_17286, n_17287);
  not g36989 (n_17288, n20084);
  not g36990 (n_17289, n20085);
  and g36991 (n20086, n_17288, n_17289);
  and g36992 (n20087, n_17070, n_17071);
  not g36993 (n_17290, n20087);
  and g36994 (n20088, n_17059, n_17290);
  not g36995 (n_17291, n20086);
  not g36996 (n_17292, n20088);
  and g36997 (n20089, n_17291, n_17292);
  and g36998 (n20090, n20086, n20088);
  not g36999 (n_17293, n20089);
  not g37000 (n_17294, n20090);
  and g37001 (n20091, n_17293, n_17294);
  not g37002 (n_17295, n20075);
  and g37003 (n20092, n_17295, n20091);
  not g37004 (n_17296, n20091);
  and g37005 (n20093, n20075, n_17296);
  not g37006 (n_17297, n20092);
  not g37007 (n_17298, n20093);
  and g37008 (n20094, n_17297, n_17298);
  and g37009 (n20095, \b[36] , n7446);
  and g37010 (n20096, \b[34] , n7787);
  and g37011 (n20097, \b[35] , n7441);
  and g37017 (n20100, n4922, n7449);
  not g37020 (n_17303, n20101);
  and g37021 (n20102, \a[47] , n_17303);
  not g37022 (n_17304, n20102);
  and g37023 (n20103, \a[47] , n_17304);
  and g37024 (n20104, n_17303, n_17304);
  not g37025 (n_17305, n20103);
  not g37026 (n_17306, n20104);
  and g37027 (n20105, n_17305, n_17306);
  not g37028 (n_17307, n20094);
  not g37029 (n_17308, n20105);
  and g37030 (n20106, n_17307, n_17308);
  and g37031 (n20107, n20094, n20105);
  not g37032 (n_17309, n20106);
  not g37033 (n_17310, n20107);
  and g37034 (n20108, n_17309, n_17310);
  not g37035 (n_17311, n20108);
  and g37036 (n20109, n19991, n_17311);
  not g37037 (n_17312, n19991);
  and g37038 (n20110, n_17312, n20108);
  not g37039 (n_17313, n20109);
  not g37040 (n_17314, n20110);
  and g37041 (n20111, n_17313, n_17314);
  and g37042 (n20112, \b[39] , n6595);
  and g37043 (n20113, \b[37] , n6902);
  and g37044 (n20114, \b[38] , n6590);
  and g37050 (n20117, n5451, n6598);
  not g37053 (n_17319, n20118);
  and g37054 (n20119, \a[44] , n_17319);
  not g37055 (n_17320, n20119);
  and g37056 (n20120, \a[44] , n_17320);
  and g37057 (n20121, n_17319, n_17320);
  not g37058 (n_17321, n20120);
  not g37059 (n_17322, n20121);
  and g37060 (n20122, n_17321, n_17322);
  not g37061 (n_17323, n20122);
  and g37062 (n20123, n20111, n_17323);
  not g37063 (n_17324, n20123);
  and g37064 (n20124, n20111, n_17324);
  and g37065 (n20125, n_17323, n_17324);
  not g37066 (n_17325, n20124);
  not g37067 (n_17326, n20125);
  and g37068 (n20126, n_17325, n_17326);
  not g37069 (n_17327, n19990);
  and g37070 (n20127, n_17327, n20126);
  not g37071 (n_17328, n20126);
  and g37072 (n20128, n19990, n_17328);
  not g37073 (n_17329, n20127);
  not g37074 (n_17330, n20128);
  and g37075 (n20129, n_17329, n_17330);
  and g37076 (n20130, \b[42] , n5777);
  and g37077 (n20131, \b[40] , n6059);
  and g37078 (n20132, \b[41] , n5772);
  and g37084 (n20135, n5780, n6489);
  not g37087 (n_17335, n20136);
  and g37088 (n20137, \a[41] , n_17335);
  not g37089 (n_17336, n20137);
  and g37090 (n20138, \a[41] , n_17336);
  and g37091 (n20139, n_17335, n_17336);
  not g37092 (n_17337, n20138);
  not g37093 (n_17338, n20139);
  and g37094 (n20140, n_17337, n_17338);
  not g37095 (n_17339, n20129);
  not g37096 (n_17340, n20140);
  and g37097 (n20141, n_17339, n_17340);
  and g37098 (n20142, n20129, n20140);
  not g37099 (n_17341, n20141);
  not g37100 (n_17342, n20142);
  and g37101 (n20143, n_17341, n_17342);
  not g37102 (n_17343, n20143);
  and g37103 (n20144, n19988, n_17343);
  not g37104 (n_17344, n19988);
  and g37105 (n20145, n_17344, n20143);
  not g37106 (n_17345, n20144);
  not g37107 (n_17346, n20145);
  and g37108 (n20146, n_17345, n_17346);
  and g37109 (n20147, \b[45] , n5035);
  and g37110 (n20148, \b[43] , n5277);
  and g37111 (n20149, \b[44] , n5030);
  and g37117 (n20152, n5038, n7361);
  not g37120 (n_17351, n20153);
  and g37121 (n20154, \a[38] , n_17351);
  not g37122 (n_17352, n20154);
  and g37123 (n20155, \a[38] , n_17352);
  and g37124 (n20156, n_17351, n_17352);
  not g37125 (n_17353, n20155);
  not g37126 (n_17354, n20156);
  and g37127 (n20157, n_17353, n_17354);
  not g37128 (n_17355, n20157);
  and g37129 (n20158, n20146, n_17355);
  not g37130 (n_17356, n20158);
  and g37131 (n20159, n20146, n_17356);
  and g37132 (n20160, n_17355, n_17356);
  not g37133 (n_17357, n20159);
  not g37134 (n_17358, n20160);
  and g37135 (n20161, n_17357, n_17358);
  and g37136 (n20162, n_17117, n_17121);
  and g37137 (n20163, n20161, n20162);
  not g37138 (n_17359, n20161);
  not g37139 (n_17360, n20162);
  and g37140 (n20164, n_17359, n_17360);
  not g37141 (n_17361, n20163);
  not g37142 (n_17362, n20164);
  and g37143 (n20165, n_17361, n_17362);
  and g37144 (n20166, \b[48] , n4287);
  and g37145 (n20167, \b[46] , n4532);
  and g37146 (n20168, \b[47] , n4282);
  and g37152 (n20171, n4290, n8009);
  not g37155 (n_17367, n20172);
  and g37156 (n20173, \a[35] , n_17367);
  not g37157 (n_17368, n20173);
  and g37158 (n20174, \a[35] , n_17368);
  and g37159 (n20175, n_17367, n_17368);
  not g37160 (n_17369, n20174);
  not g37161 (n_17370, n20175);
  and g37162 (n20176, n_17369, n_17370);
  not g37163 (n_17371, n20176);
  and g37164 (n20177, n20165, n_17371);
  not g37165 (n_17372, n20177);
  and g37166 (n20178, n20165, n_17372);
  and g37167 (n20179, n_17371, n_17372);
  not g37168 (n_17373, n20178);
  not g37169 (n_17374, n20179);
  and g37170 (n20180, n_17373, n_17374);
  and g37171 (n20181, n_17125, n_17136);
  and g37172 (n20182, n20180, n20181);
  not g37173 (n_17375, n20180);
  not g37174 (n_17376, n20181);
  and g37175 (n20183, n_17375, n_17376);
  not g37176 (n_17377, n20182);
  not g37177 (n_17378, n20183);
  and g37178 (n20184, n_17377, n_17378);
  and g37179 (n20185, \b[51] , n3638);
  and g37180 (n20186, \b[49] , n3843);
  and g37181 (n20187, \b[50] , n3633);
  and g37187 (n20190, n3641, n8976);
  not g37190 (n_17383, n20191);
  and g37191 (n20192, \a[32] , n_17383);
  not g37192 (n_17384, n20192);
  and g37193 (n20193, \a[32] , n_17384);
  and g37194 (n20194, n_17383, n_17384);
  not g37195 (n_17385, n20193);
  not g37196 (n_17386, n20194);
  and g37197 (n20195, n_17385, n_17386);
  and g37198 (n20196, n_16974, n_17143);
  not g37199 (n_17387, n20195);
  not g37200 (n_17388, n20196);
  and g37201 (n20197, n_17387, n_17388);
  and g37202 (n20198, n20195, n20196);
  not g37203 (n_17389, n20197);
  not g37204 (n_17390, n20198);
  and g37205 (n20199, n_17389, n_17390);
  and g37206 (n20200, n20184, n20199);
  not g37207 (n_17391, n20200);
  and g37208 (n20201, n20184, n_17391);
  and g37209 (n20202, n20199, n_17391);
  not g37210 (n_17392, n20201);
  not g37211 (n_17393, n20202);
  and g37212 (n20203, n_17392, n_17393);
  not g37213 (n_17394, n20203);
  and g37214 (n20204, n19987, n_17394);
  not g37215 (n_17395, n20204);
  and g37216 (n20205, n19987, n_17395);
  and g37217 (n20206, n_17394, n_17395);
  not g37218 (n_17396, n20205);
  not g37219 (n_17397, n20206);
  and g37220 (n20207, n_17396, n_17397);
  and g37221 (n20208, \b[57] , n2539);
  and g37222 (n20209, \b[55] , n2685);
  and g37223 (n20210, \b[56] , n2534);
  and g37229 (n20213, n2542, n11410);
  not g37232 (n_17402, n20214);
  and g37233 (n20215, \a[26] , n_17402);
  not g37234 (n_17403, n20215);
  and g37235 (n20216, \a[26] , n_17403);
  and g37236 (n20217, n_17402, n_17403);
  not g37237 (n_17404, n20216);
  not g37238 (n_17405, n20217);
  and g37239 (n20218, n_17404, n_17405);
  and g37240 (n20219, n_16949, n_17151);
  not g37241 (n_17406, n20218);
  not g37242 (n_17407, n20219);
  and g37243 (n20220, n_17406, n_17407);
  and g37244 (n20221, n20218, n20219);
  not g37245 (n_17408, n20220);
  not g37246 (n_17409, n20221);
  and g37247 (n20222, n_17408, n_17409);
  not g37248 (n_17410, n20207);
  and g37249 (n20223, n_17410, n20222);
  not g37250 (n_17411, n20223);
  and g37251 (n20224, n_17410, n_17411);
  and g37252 (n20225, n20222, n_17411);
  not g37253 (n_17412, n20224);
  not g37254 (n_17413, n20225);
  and g37255 (n20226, n_17412, n_17413);
  not g37256 (n_17414, n20226);
  and g37257 (n20227, n19972, n_17414);
  not g37258 (n_17415, n20227);
  and g37259 (n20228, n19972, n_17415);
  and g37260 (n20229, n_17414, n_17415);
  not g37261 (n_17416, n20228);
  not g37262 (n_17417, n20229);
  and g37263 (n20230, n_17416, n_17417);
  not g37264 (n_17418, n19957);
  and g37265 (n20231, n_17418, n20230);
  not g37266 (n_17419, n20230);
  and g37267 (n20232, n19957, n_17419);
  not g37268 (n_17420, n20231);
  not g37269 (n_17421, n20232);
  and g37270 (n20233, n_17420, n_17421);
  not g37271 (n_17422, n19941);
  not g37272 (n_17423, n20233);
  and g37273 (n20234, n_17422, n_17423);
  not g37274 (n_17424, n20234);
  and g37275 (n20235, n_17422, n_17424);
  and g37276 (n20236, n_17423, n_17424);
  not g37277 (n_17425, n20235);
  not g37278 (n_17426, n20236);
  and g37279 (n20237, n_17425, n_17426);
  not g37280 (n_17427, n19940);
  not g37281 (n_17428, n20237);
  and g37282 (n20238, n_17427, n_17428);
  and g37283 (n20239, n19940, n_17426);
  and g37284 (n20240, n_17425, n20239);
  not g37285 (n_17429, n20238);
  not g37286 (n_17430, n20240);
  and g37287 (\f[81] , n_17429, n_17430);
  and g37288 (n20242, n_17424, n_17429);
  and g37289 (n20243, n_17418, n_17419);
  not g37290 (n_17431, n20243);
  and g37291 (n20244, n_17181, n_17431);
  and g37292 (n20245, \b[61] , n2048);
  and g37293 (n20246, \b[59] , n2198);
  and g37294 (n20247, \b[60] , n2043);
  and g37300 (n20250, n2051, n12969);
  not g37303 (n_17436, n20251);
  and g37304 (n20252, \a[23] , n_17436);
  not g37305 (n_17437, n20252);
  and g37306 (n20253, \a[23] , n_17437);
  and g37307 (n20254, n_17436, n_17437);
  not g37308 (n_17438, n20253);
  not g37309 (n_17439, n20254);
  and g37310 (n20255, n_17438, n_17439);
  and g37311 (n20256, n_17408, n_17411);
  and g37312 (n20257, n20255, n20256);
  not g37313 (n_17440, n20255);
  not g37314 (n_17441, n20256);
  and g37315 (n20258, n_17440, n_17441);
  not g37316 (n_17442, n20257);
  not g37317 (n_17443, n20258);
  and g37318 (n20259, n_17442, n_17443);
  and g37319 (n20260, \b[58] , n2539);
  and g37320 (n20261, \b[56] , n2685);
  and g37321 (n20262, \b[57] , n2534);
  and g37327 (n20265, n2542, n11436);
  not g37330 (n_17448, n20266);
  and g37331 (n20267, \a[26] , n_17448);
  not g37332 (n_17449, n20267);
  and g37333 (n20268, \a[26] , n_17449);
  and g37334 (n20269, n_17448, n_17449);
  not g37335 (n_17450, n20268);
  not g37336 (n_17451, n20269);
  and g37337 (n20270, n_17450, n_17451);
  and g37338 (n20271, n_17207, n_17395);
  and g37339 (n20272, n20270, n20271);
  not g37340 (n_17452, n20270);
  not g37341 (n_17453, n20271);
  and g37342 (n20273, n_17452, n_17453);
  not g37343 (n_17454, n20272);
  not g37344 (n_17455, n20273);
  and g37345 (n20274, n_17454, n_17455);
  and g37346 (n20275, \b[55] , n3050);
  and g37347 (n20276, \b[53] , n3243);
  and g37348 (n20277, \b[54] , n3045);
  and g37354 (n20280, n3053, n10684);
  not g37357 (n_17460, n20281);
  and g37358 (n20282, \a[29] , n_17460);
  not g37359 (n_17461, n20282);
  and g37360 (n20283, \a[29] , n_17461);
  and g37361 (n20284, n_17460, n_17461);
  not g37362 (n_17462, n20283);
  not g37363 (n_17463, n20284);
  and g37364 (n20285, n_17462, n_17463);
  and g37365 (n20286, n_17389, n_17391);
  and g37366 (n20287, n20285, n20286);
  not g37367 (n_17464, n20285);
  not g37368 (n_17465, n20286);
  and g37369 (n20288, n_17464, n_17465);
  not g37370 (n_17466, n20287);
  not g37371 (n_17467, n20288);
  and g37372 (n20289, n_17466, n_17467);
  and g37373 (n20290, \b[52] , n3638);
  and g37374 (n20291, \b[50] , n3843);
  and g37375 (n20292, \b[51] , n3633);
  and g37381 (n20295, n3641, n9628);
  not g37384 (n_17472, n20296);
  and g37385 (n20297, \a[32] , n_17472);
  not g37386 (n_17473, n20297);
  and g37387 (n20298, \a[32] , n_17473);
  and g37388 (n20299, n_17472, n_17473);
  not g37389 (n_17474, n20298);
  not g37390 (n_17475, n20299);
  and g37391 (n20300, n_17474, n_17475);
  and g37392 (n20301, n_17372, n_17378);
  and g37393 (n20302, n20300, n20301);
  not g37394 (n_17476, n20300);
  not g37395 (n_17477, n20301);
  and g37396 (n20303, n_17476, n_17477);
  not g37397 (n_17478, n20302);
  not g37398 (n_17479, n20303);
  and g37399 (n20304, n_17478, n_17479);
  and g37400 (n20305, \b[43] , n5777);
  and g37401 (n20306, \b[41] , n6059);
  and g37402 (n20307, \b[42] , n5772);
  and g37408 (n20310, n5780, n6515);
  not g37411 (n_17484, n20311);
  and g37412 (n20312, \a[41] , n_17484);
  not g37413 (n_17485, n20312);
  and g37414 (n20313, \a[41] , n_17485);
  and g37415 (n20314, n_17484, n_17485);
  not g37416 (n_17486, n20313);
  not g37417 (n_17487, n20314);
  and g37418 (n20315, n_17486, n_17487);
  and g37419 (n20316, n_17327, n_17328);
  not g37420 (n_17488, n20316);
  and g37421 (n20317, n_17324, n_17488);
  and g37422 (n20318, \b[40] , n6595);
  and g37423 (n20319, \b[38] , n6902);
  and g37424 (n20320, \b[39] , n6590);
  and g37430 (n20323, n5955, n6598);
  not g37433 (n_17493, n20324);
  and g37434 (n20325, \a[44] , n_17493);
  not g37435 (n_17494, n20325);
  and g37436 (n20326, \a[44] , n_17494);
  and g37437 (n20327, n_17493, n_17494);
  not g37438 (n_17495, n20326);
  not g37439 (n_17496, n20327);
  and g37440 (n20328, n_17495, n_17496);
  and g37441 (n20329, n_17309, n_17314);
  and g37442 (n20330, \b[31] , n9339);
  and g37443 (n20331, \b[29] , n9732);
  and g37444 (n20332, \b[30] , n9334);
  and g37450 (n20335, n3796, n9342);
  not g37453 (n_17501, n20336);
  and g37454 (n20337, \a[53] , n_17501);
  not g37455 (n_17502, n20337);
  and g37456 (n20338, \a[53] , n_17502);
  and g37457 (n20339, n_17501, n_17502);
  not g37458 (n_17503, n20338);
  not g37459 (n_17504, n20339);
  and g37460 (n20340, n_17503, n_17504);
  and g37461 (n20341, n_17253, n_17256);
  and g37462 (n20342, \b[25] , n11531);
  and g37463 (n20343, \b[23] , n11896);
  and g37464 (n20344, \b[24] , n11526);
  and g37470 (n20347, n2485, n11534);
  not g37473 (n_17509, n20348);
  and g37474 (n20349, \a[59] , n_17509);
  not g37475 (n_17510, n20349);
  and g37476 (n20350, \a[59] , n_17510);
  and g37477 (n20351, n_17509, n_17510);
  not g37478 (n_17511, n20350);
  not g37479 (n_17512, n20351);
  and g37480 (n20352, n_17511, n_17512);
  and g37481 (n20353, \b[18] , n13903);
  and g37482 (n20354, \b[19] , n_11555);
  not g37483 (n_17513, n20353);
  not g37484 (n_17514, n20354);
  and g37485 (n20355, n_17513, n_17514);
  and g37486 (n20356, n_17228, n_17231);
  not g37487 (n_17515, n20355);
  and g37488 (n20357, n_17515, n20356);
  not g37489 (n_17516, n20356);
  and g37490 (n20358, n20355, n_17516);
  not g37491 (n_17517, n20357);
  not g37492 (n_17518, n20358);
  and g37493 (n20359, n_17517, n_17518);
  and g37494 (n20360, \b[22] , n12668);
  and g37495 (n20361, \b[20] , n13047);
  and g37496 (n20362, \b[21] , n12663);
  and g37502 (n20365, n2145, n12671);
  not g37505 (n_17523, n20366);
  and g37506 (n20367, \a[62] , n_17523);
  not g37507 (n_17524, n20367);
  and g37508 (n20368, \a[62] , n_17524);
  and g37509 (n20369, n_17523, n_17524);
  not g37510 (n_17525, n20368);
  not g37511 (n_17526, n20369);
  and g37512 (n20370, n_17525, n_17526);
  not g37513 (n_17527, n20359);
  and g37514 (n20371, n_17527, n20370);
  not g37515 (n_17528, n20370);
  and g37516 (n20372, n20359, n_17528);
  not g37517 (n_17529, n20371);
  not g37518 (n_17530, n20372);
  and g37519 (n20373, n_17529, n_17530);
  and g37520 (n20374, n_17234, n_17239);
  not g37521 (n_17531, n20374);
  and g37522 (n20375, n20373, n_17531);
  not g37523 (n_17532, n20373);
  and g37524 (n20376, n_17532, n20374);
  not g37525 (n_17533, n20375);
  not g37526 (n_17534, n20376);
  and g37527 (n20377, n_17533, n_17534);
  not g37528 (n_17535, n20352);
  and g37529 (n20378, n_17535, n20377);
  not g37530 (n_17536, n20378);
  and g37531 (n20379, n20377, n_17536);
  and g37532 (n20380, n_17535, n_17536);
  not g37533 (n_17537, n20379);
  not g37534 (n_17538, n20380);
  and g37535 (n20381, n_17537, n_17538);
  not g37536 (n_17539, n20341);
  and g37537 (n20382, n_17539, n20381);
  not g37538 (n_17540, n20381);
  and g37539 (n20383, n20341, n_17540);
  not g37540 (n_17541, n20382);
  not g37541 (n_17542, n20383);
  and g37542 (n20384, n_17541, n_17542);
  and g37543 (n20385, \b[28] , n10426);
  and g37544 (n20386, \b[26] , n10796);
  and g37545 (n20387, \b[27] , n10421);
  and g37551 (n20390, n3189, n10429);
  not g37554 (n_17547, n20391);
  and g37555 (n20392, \a[56] , n_17547);
  not g37556 (n_17548, n20392);
  and g37557 (n20393, \a[56] , n_17548);
  and g37558 (n20394, n_17547, n_17548);
  not g37559 (n_17549, n20393);
  not g37560 (n_17550, n20394);
  and g37561 (n20395, n_17549, n_17550);
  and g37562 (n20396, n20384, n20395);
  not g37563 (n_17551, n20384);
  not g37564 (n_17552, n20395);
  and g37565 (n20397, n_17551, n_17552);
  not g37566 (n_17553, n20396);
  not g37567 (n_17554, n20397);
  and g37568 (n20398, n_17553, n_17554);
  and g37569 (n20399, n_17259, n_17265);
  not g37570 (n_17555, n20399);
  and g37571 (n20400, n20398, n_17555);
  not g37572 (n_17556, n20398);
  and g37573 (n20401, n_17556, n20399);
  not g37574 (n_17557, n20400);
  not g37575 (n_17558, n20401);
  and g37576 (n20402, n_17557, n_17558);
  not g37577 (n_17559, n20340);
  and g37578 (n20403, n_17559, n20402);
  not g37579 (n_17560, n20403);
  and g37580 (n20404, n20402, n_17560);
  and g37581 (n20405, n_17559, n_17560);
  not g37582 (n_17561, n20404);
  not g37583 (n_17562, n20405);
  and g37584 (n20406, n_17561, n_17562);
  and g37585 (n20407, n_17275, n_17281);
  and g37586 (n20408, n20406, n20407);
  not g37587 (n_17563, n20406);
  not g37588 (n_17564, n20407);
  and g37589 (n20409, n_17563, n_17564);
  not g37590 (n_17565, n20408);
  not g37591 (n_17566, n20409);
  and g37592 (n20410, n_17565, n_17566);
  and g37593 (n20411, \b[34] , n8362);
  and g37594 (n20412, \b[32] , n8715);
  and g37595 (n20413, \b[33] , n8357);
  and g37601 (n20416, n4466, n8365);
  not g37604 (n_17571, n20417);
  and g37605 (n20418, \a[50] , n_17571);
  not g37606 (n_17572, n20418);
  and g37607 (n20419, \a[50] , n_17572);
  and g37608 (n20420, n_17571, n_17572);
  not g37609 (n_17573, n20419);
  not g37610 (n_17574, n20420);
  and g37611 (n20421, n_17573, n_17574);
  not g37612 (n_17575, n20421);
  and g37613 (n20422, n20410, n_17575);
  not g37614 (n_17576, n20422);
  and g37615 (n20423, n20410, n_17576);
  and g37616 (n20424, n_17575, n_17576);
  not g37617 (n_17577, n20423);
  not g37618 (n_17578, n20424);
  and g37619 (n20425, n_17577, n_17578);
  and g37620 (n20426, n20075, n20091);
  not g37621 (n_17579, n20426);
  and g37622 (n20427, n_17293, n_17579);
  and g37623 (n20428, n20425, n20427);
  not g37624 (n_17580, n20425);
  not g37625 (n_17581, n20427);
  and g37626 (n20429, n_17580, n_17581);
  not g37627 (n_17582, n20428);
  not g37628 (n_17583, n20429);
  and g37629 (n20430, n_17582, n_17583);
  and g37630 (n20431, \b[37] , n7446);
  and g37631 (n20432, \b[35] , n7787);
  and g37632 (n20433, \b[36] , n7441);
  and g37638 (n20436, n5181, n7449);
  not g37641 (n_17588, n20437);
  and g37642 (n20438, \a[47] , n_17588);
  not g37643 (n_17589, n20438);
  and g37644 (n20439, \a[47] , n_17589);
  and g37645 (n20440, n_17588, n_17589);
  not g37646 (n_17590, n20439);
  not g37647 (n_17591, n20440);
  and g37648 (n20441, n_17590, n_17591);
  not g37649 (n_17592, n20430);
  and g37650 (n20442, n_17592, n20441);
  not g37651 (n_17593, n20441);
  and g37652 (n20443, n20430, n_17593);
  not g37653 (n_17594, n20442);
  not g37654 (n_17595, n20443);
  and g37655 (n20444, n_17594, n_17595);
  not g37656 (n_17596, n20329);
  and g37657 (n20445, n_17596, n20444);
  not g37658 (n_17597, n20445);
  and g37659 (n20446, n_17596, n_17597);
  and g37660 (n20447, n20444, n_17597);
  not g37661 (n_17598, n20446);
  not g37662 (n_17599, n20447);
  and g37663 (n20448, n_17598, n_17599);
  not g37664 (n_17600, n20328);
  not g37665 (n_17601, n20448);
  and g37666 (n20449, n_17600, n_17601);
  and g37667 (n20450, n20328, n_17599);
  and g37668 (n20451, n_17598, n20450);
  not g37669 (n_17602, n20449);
  not g37670 (n_17603, n20451);
  and g37671 (n20452, n_17602, n_17603);
  not g37672 (n_17604, n20317);
  and g37673 (n20453, n_17604, n20452);
  not g37674 (n_17605, n20452);
  and g37675 (n20454, n20317, n_17605);
  not g37676 (n_17606, n20453);
  not g37677 (n_17607, n20454);
  and g37678 (n20455, n_17606, n_17607);
  not g37679 (n_17608, n20315);
  and g37680 (n20456, n_17608, n20455);
  not g37681 (n_17609, n20456);
  and g37682 (n20457, n20455, n_17609);
  and g37683 (n20458, n_17608, n_17609);
  not g37684 (n_17610, n20457);
  not g37685 (n_17611, n20458);
  and g37686 (n20459, n_17610, n_17611);
  and g37687 (n20460, n_17341, n_17346);
  and g37688 (n20461, n20459, n20460);
  not g37689 (n_17612, n20459);
  not g37690 (n_17613, n20460);
  and g37691 (n20462, n_17612, n_17613);
  not g37692 (n_17614, n20461);
  not g37693 (n_17615, n20462);
  and g37694 (n20463, n_17614, n_17615);
  and g37695 (n20464, \b[46] , n5035);
  and g37696 (n20465, \b[44] , n5277);
  and g37697 (n20466, \b[45] , n5030);
  and g37703 (n20469, n5038, n7677);
  not g37706 (n_17620, n20470);
  and g37707 (n20471, \a[38] , n_17620);
  not g37708 (n_17621, n20471);
  and g37709 (n20472, \a[38] , n_17621);
  and g37710 (n20473, n_17620, n_17621);
  not g37711 (n_17622, n20472);
  not g37712 (n_17623, n20473);
  and g37713 (n20474, n_17622, n_17623);
  not g37714 (n_17624, n20474);
  and g37715 (n20475, n20463, n_17624);
  not g37716 (n_17625, n20475);
  and g37717 (n20476, n20463, n_17625);
  and g37718 (n20477, n_17624, n_17625);
  not g37719 (n_17626, n20476);
  not g37720 (n_17627, n20477);
  and g37721 (n20478, n_17626, n_17627);
  and g37722 (n20479, n_17356, n_17362);
  and g37723 (n20480, n20478, n20479);
  not g37724 (n_17628, n20478);
  not g37725 (n_17629, n20479);
  and g37726 (n20481, n_17628, n_17629);
  not g37727 (n_17630, n20480);
  not g37728 (n_17631, n20481);
  and g37729 (n20482, n_17630, n_17631);
  and g37730 (n20483, \b[49] , n4287);
  and g37731 (n20484, \b[47] , n4532);
  and g37732 (n20485, \b[48] , n4282);
  and g37738 (n20488, n4290, n8625);
  not g37741 (n_17636, n20489);
  and g37742 (n20490, \a[35] , n_17636);
  not g37743 (n_17637, n20490);
  and g37744 (n20491, \a[35] , n_17637);
  and g37745 (n20492, n_17636, n_17637);
  not g37746 (n_17638, n20491);
  not g37747 (n_17639, n20492);
  and g37748 (n20493, n_17638, n_17639);
  not g37749 (n_17640, n20493);
  and g37750 (n20494, n20482, n_17640);
  not g37751 (n_17641, n20494);
  and g37752 (n20495, n20482, n_17641);
  and g37753 (n20496, n_17640, n_17641);
  not g37754 (n_17642, n20495);
  not g37755 (n_17643, n20496);
  and g37756 (n20497, n_17642, n_17643);
  not g37757 (n_17644, n20497);
  and g37758 (n20498, n20304, n_17644);
  not g37759 (n_17645, n20304);
  and g37760 (n20499, n_17645, n20497);
  not g37761 (n_17646, n20499);
  and g37762 (n20500, n20289, n_17646);
  not g37763 (n_17647, n20498);
  and g37764 (n20501, n_17647, n20500);
  not g37765 (n_17648, n20501);
  and g37766 (n20502, n20289, n_17648);
  and g37767 (n20503, n_17646, n_17648);
  and g37768 (n20504, n_17647, n20503);
  not g37769 (n_17649, n20502);
  not g37770 (n_17650, n20504);
  and g37771 (n20505, n_17649, n_17650);
  not g37772 (n_17651, n20505);
  and g37773 (n20506, n20274, n_17651);
  not g37774 (n_17652, n20274);
  and g37775 (n20507, n_17652, n20505);
  not g37776 (n_17653, n20507);
  and g37777 (n20508, n20259, n_17653);
  not g37778 (n_17654, n20506);
  and g37779 (n20509, n_17654, n20508);
  not g37780 (n_17655, n20509);
  and g37781 (n20510, n20259, n_17655);
  and g37782 (n20511, n_17653, n_17655);
  and g37783 (n20512, n_17654, n20511);
  not g37784 (n_17656, n20510);
  not g37785 (n_17657, n20512);
  and g37786 (n20513, n_17656, n_17657);
  and g37787 (n20514, n_17195, n_17415);
  and g37788 (n20515, \b[62] , n1763);
  and g37789 (n20516, \b[63] , n1622);
  not g37790 (n_17658, n20515);
  not g37791 (n_17659, n20516);
  and g37792 (n20517, n_17658, n_17659);
  and g37793 (n20518, n_14471, n20517);
  and g37794 (n20519, n13800, n20517);
  not g37795 (n_17660, n20518);
  not g37796 (n_17661, n20519);
  and g37797 (n20520, n_17660, n_17661);
  not g37798 (n_17662, n20520);
  and g37799 (n20521, \a[20] , n_17662);
  and g37800 (n20522, n_1221, n20520);
  not g37801 (n_17663, n20521);
  not g37802 (n_17664, n20522);
  and g37803 (n20523, n_17663, n_17664);
  not g37804 (n_17665, n20514);
  not g37805 (n_17666, n20523);
  and g37806 (n20524, n_17665, n_17666);
  not g37807 (n_17667, n20524);
  and g37808 (n20525, n_17665, n_17667);
  and g37809 (n20526, n_17666, n_17667);
  not g37810 (n_17668, n20525);
  not g37811 (n_17669, n20526);
  and g37812 (n20527, n_17668, n_17669);
  not g37813 (n_17670, n20513);
  not g37814 (n_17671, n20527);
  and g37815 (n20528, n_17670, n_17671);
  and g37816 (n20529, n20513, n_17669);
  and g37817 (n20530, n_17668, n20529);
  not g37818 (n_17672, n20528);
  not g37819 (n_17673, n20530);
  and g37820 (n20531, n_17672, n_17673);
  not g37821 (n_17674, n20244);
  and g37822 (n20532, n_17674, n20531);
  not g37823 (n_17675, n20532);
  and g37824 (n20533, n_17674, n_17675);
  and g37825 (n20534, n20531, n_17675);
  not g37826 (n_17676, n20533);
  not g37827 (n_17677, n20534);
  and g37828 (n20535, n_17676, n_17677);
  not g37829 (n_17678, n20242);
  not g37830 (n_17679, n20535);
  and g37831 (n20536, n_17678, n_17679);
  and g37832 (n20537, n20242, n_17677);
  and g37833 (n20538, n_17676, n20537);
  not g37834 (n_17680, n20536);
  not g37835 (n_17681, n20538);
  and g37836 (\f[82] , n_17680, n_17681);
  and g37837 (n20540, n_17675, n_17680);
  and g37838 (n20541, n_17667, n_17672);
  and g37839 (n20542, n_17443, n_17655);
  and g37840 (n20543, \b[63] , n1763);
  and g37841 (n20544, n1630, n13797);
  not g37842 (n_17682, n20543);
  not g37843 (n_17683, n20544);
  and g37844 (n20545, n_17682, n_17683);
  not g37845 (n_17684, n20545);
  and g37846 (n20546, \a[20] , n_17684);
  not g37847 (n_17685, n20546);
  and g37848 (n20547, \a[20] , n_17685);
  and g37849 (n20548, n_17684, n_17685);
  not g37850 (n_17686, n20547);
  not g37851 (n_17687, n20548);
  and g37852 (n20549, n_17686, n_17687);
  not g37853 (n_17688, n20542);
  not g37854 (n_17689, n20549);
  and g37855 (n20550, n_17688, n_17689);
  not g37856 (n_17690, n20550);
  and g37857 (n20551, n_17688, n_17690);
  and g37858 (n20552, n_17689, n_17690);
  not g37859 (n_17691, n20551);
  not g37860 (n_17692, n20552);
  and g37861 (n20553, n_17691, n_17692);
  and g37862 (n20554, \b[62] , n2048);
  and g37863 (n20555, \b[60] , n2198);
  and g37864 (n20556, \b[61] , n2043);
  and g37870 (n20559, n2051, n13370);
  not g37873 (n_17697, n20560);
  and g37874 (n20561, \a[23] , n_17697);
  not g37875 (n_17698, n20561);
  and g37876 (n20562, \a[23] , n_17698);
  and g37877 (n20563, n_17697, n_17698);
  not g37878 (n_17699, n20562);
  not g37879 (n_17700, n20563);
  and g37880 (n20564, n_17699, n_17700);
  and g37881 (n20565, n_17455, n_17654);
  not g37882 (n_17701, n20564);
  not g37883 (n_17702, n20565);
  and g37884 (n20566, n_17701, n_17702);
  not g37885 (n_17703, n20566);
  and g37886 (n20567, n_17701, n_17703);
  and g37887 (n20568, n_17702, n_17703);
  not g37888 (n_17704, n20567);
  not g37889 (n_17705, n20568);
  and g37890 (n20569, n_17704, n_17705);
  and g37891 (n20570, \b[59] , n2539);
  and g37892 (n20571, \b[57] , n2685);
  and g37893 (n20572, \b[58] , n2534);
  and g37899 (n20575, n2542, n12179);
  not g37902 (n_17710, n20576);
  and g37903 (n20577, \a[26] , n_17710);
  not g37904 (n_17711, n20577);
  and g37905 (n20578, \a[26] , n_17711);
  and g37906 (n20579, n_17710, n_17711);
  not g37907 (n_17712, n20578);
  not g37908 (n_17713, n20579);
  and g37909 (n20580, n_17712, n_17713);
  and g37910 (n20581, n_17467, n_17648);
  and g37911 (n20582, n20580, n20581);
  not g37912 (n_17714, n20580);
  not g37913 (n_17715, n20581);
  and g37914 (n20583, n_17714, n_17715);
  not g37915 (n_17716, n20582);
  not g37916 (n_17717, n20583);
  and g37917 (n20584, n_17716, n_17717);
  and g37918 (n20585, \b[56] , n3050);
  and g37919 (n20586, \b[54] , n3243);
  and g37920 (n20587, \b[55] , n3045);
  and g37926 (n20590, n3053, n10708);
  not g37929 (n_17722, n20591);
  and g37930 (n20592, \a[29] , n_17722);
  not g37931 (n_17723, n20592);
  and g37932 (n20593, \a[29] , n_17723);
  and g37933 (n20594, n_17722, n_17723);
  not g37934 (n_17724, n20593);
  not g37935 (n_17725, n20594);
  and g37936 (n20595, n_17724, n_17725);
  and g37937 (n20596, n_17479, n_17647);
  not g37938 (n_17726, n20595);
  not g37939 (n_17727, n20596);
  and g37940 (n20597, n_17726, n_17727);
  not g37941 (n_17728, n20597);
  and g37942 (n20598, n_17726, n_17728);
  and g37943 (n20599, n_17727, n_17728);
  not g37944 (n_17729, n20598);
  not g37945 (n_17730, n20599);
  and g37946 (n20600, n_17729, n_17730);
  and g37947 (n20601, \b[53] , n3638);
  and g37948 (n20602, \b[51] , n3843);
  and g37949 (n20603, \b[52] , n3633);
  and g37955 (n20606, n3641, n9972);
  not g37958 (n_17735, n20607);
  and g37959 (n20608, \a[32] , n_17735);
  not g37960 (n_17736, n20608);
  and g37961 (n20609, \a[32] , n_17736);
  and g37962 (n20610, n_17735, n_17736);
  not g37963 (n_17737, n20609);
  not g37964 (n_17738, n20610);
  and g37965 (n20611, n_17737, n_17738);
  and g37966 (n20612, n_17631, n_17641);
  and g37967 (n20613, n20611, n20612);
  not g37968 (n_17739, n20611);
  not g37969 (n_17740, n20612);
  and g37970 (n20614, n_17739, n_17740);
  not g37971 (n_17741, n20613);
  not g37972 (n_17742, n20614);
  and g37973 (n20615, n_17741, n_17742);
  and g37974 (n20616, n_17606, n_17609);
  and g37975 (n20617, \b[44] , n5777);
  and g37976 (n20618, \b[42] , n6059);
  and g37977 (n20619, \b[43] , n5772);
  and g37983 (n20622, n5780, n7072);
  not g37986 (n_17747, n20623);
  and g37987 (n20624, \a[41] , n_17747);
  not g37988 (n_17748, n20624);
  and g37989 (n20625, \a[41] , n_17748);
  and g37990 (n20626, n_17747, n_17748);
  not g37991 (n_17749, n20625);
  not g37992 (n_17750, n20626);
  and g37993 (n20627, n_17749, n_17750);
  and g37994 (n20628, n_17597, n_17602);
  and g37995 (n20629, \b[41] , n6595);
  and g37996 (n20630, \b[39] , n6902);
  and g37997 (n20631, \b[40] , n6590);
  and g38003 (n20634, n6219, n6598);
  not g38006 (n_17755, n20635);
  and g38007 (n20636, \a[44] , n_17755);
  not g38008 (n_17756, n20636);
  and g38009 (n20637, \a[44] , n_17756);
  and g38010 (n20638, n_17755, n_17756);
  not g38011 (n_17757, n20637);
  not g38012 (n_17758, n20638);
  and g38013 (n20639, n_17757, n_17758);
  and g38014 (n20640, n_17583, n_17595);
  and g38015 (n20641, \b[38] , n7446);
  and g38016 (n20642, \b[36] , n7787);
  and g38017 (n20643, \b[37] , n7441);
  and g38023 (n20646, n5205, n7449);
  not g38026 (n_17763, n20647);
  and g38027 (n20648, \a[47] , n_17763);
  not g38028 (n_17764, n20648);
  and g38029 (n20649, \a[47] , n_17764);
  and g38030 (n20650, n_17763, n_17764);
  not g38031 (n_17765, n20649);
  not g38032 (n_17766, n20650);
  and g38033 (n20651, n_17765, n_17766);
  and g38034 (n20652, n_17566, n_17576);
  and g38035 (n20653, \b[35] , n8362);
  and g38036 (n20654, \b[33] , n8715);
  and g38037 (n20655, \b[34] , n8357);
  and g38043 (n20658, n4696, n8365);
  not g38046 (n_17771, n20659);
  and g38047 (n20660, \a[50] , n_17771);
  not g38048 (n_17772, n20660);
  and g38049 (n20661, \a[50] , n_17772);
  and g38050 (n20662, n_17771, n_17772);
  not g38051 (n_17773, n20661);
  not g38052 (n_17774, n20662);
  and g38053 (n20663, n_17773, n_17774);
  and g38054 (n20664, n_17557, n_17560);
  and g38055 (n20665, n_17533, n_17536);
  and g38056 (n20666, \b[26] , n11531);
  and g38057 (n20667, \b[24] , n11896);
  and g38058 (n20668, \b[25] , n11526);
  and g38064 (n20671, n2813, n11534);
  not g38067 (n_17779, n20672);
  and g38068 (n20673, \a[59] , n_17779);
  not g38069 (n_17780, n20673);
  and g38070 (n20674, \a[59] , n_17780);
  and g38071 (n20675, n_17779, n_17780);
  not g38072 (n_17781, n20674);
  not g38073 (n_17782, n20675);
  and g38074 (n20676, n_17781, n_17782);
  and g38075 (n20677, n_17518, n_17530);
  and g38076 (n20678, \b[19] , n13903);
  and g38077 (n20679, \b[20] , n_11555);
  not g38078 (n_17783, n20678);
  not g38079 (n_17784, n20679);
  and g38080 (n20680, n_17783, n_17784);
  and g38081 (n20681, n_17515, n20680);
  not g38082 (n_17785, n20680);
  and g38083 (n20682, n20355, n_17785);
  not g38084 (n_17786, n20681);
  not g38085 (n_17787, n20682);
  and g38086 (n20683, n_17786, n_17787);
  and g38087 (n20684, \b[23] , n12668);
  and g38088 (n20685, \b[21] , n13047);
  and g38089 (n20686, \b[22] , n12663);
  not g38090 (n_17788, n20685);
  not g38091 (n_17789, n20686);
  and g38092 (n20687, n_17788, n_17789);
  not g38093 (n_17790, n20684);
  and g38094 (n20688, n_17790, n20687);
  and g38095 (n20689, n_12644, n20688);
  not g38096 (n_17791, n2300);
  and g38097 (n20690, n_17791, n20688);
  not g38098 (n_17792, n20689);
  not g38099 (n_17793, n20690);
  and g38100 (n20691, n_17792, n_17793);
  not g38101 (n_17794, n20691);
  and g38102 (n20692, \a[62] , n_17794);
  and g38103 (n20693, n_10843, n20691);
  not g38104 (n_17795, n20692);
  not g38105 (n_17796, n20693);
  and g38106 (n20694, n_17795, n_17796);
  not g38107 (n_17797, n20694);
  and g38108 (n20695, n20683, n_17797);
  not g38109 (n_17798, n20683);
  and g38110 (n20696, n_17798, n20694);
  not g38111 (n_17799, n20695);
  not g38112 (n_17800, n20696);
  and g38113 (n20697, n_17799, n_17800);
  not g38114 (n_17801, n20677);
  and g38115 (n20698, n_17801, n20697);
  not g38116 (n_17802, n20697);
  and g38117 (n20699, n20677, n_17802);
  not g38118 (n_17803, n20698);
  not g38119 (n_17804, n20699);
  and g38120 (n20700, n_17803, n_17804);
  not g38121 (n_17805, n20676);
  and g38122 (n20701, n_17805, n20700);
  not g38123 (n_17806, n20700);
  and g38124 (n20702, n20676, n_17806);
  not g38125 (n_17807, n20701);
  not g38126 (n_17808, n20702);
  and g38127 (n20703, n_17807, n_17808);
  not g38128 (n_17809, n20665);
  and g38129 (n20704, n_17809, n20703);
  not g38130 (n_17810, n20703);
  and g38131 (n20705, n20665, n_17810);
  not g38132 (n_17811, n20704);
  not g38133 (n_17812, n20705);
  and g38134 (n20706, n_17811, n_17812);
  and g38135 (n20707, \b[29] , n10426);
  and g38136 (n20708, \b[27] , n10796);
  and g38137 (n20709, \b[28] , n10421);
  and g38143 (n20712, n3383, n10429);
  not g38146 (n_17817, n20713);
  and g38147 (n20714, \a[56] , n_17817);
  not g38148 (n_17818, n20714);
  and g38149 (n20715, \a[56] , n_17818);
  and g38150 (n20716, n_17817, n_17818);
  not g38151 (n_17819, n20715);
  not g38152 (n_17820, n20716);
  and g38153 (n20717, n_17819, n_17820);
  not g38154 (n_17821, n20717);
  and g38155 (n20718, n20706, n_17821);
  not g38156 (n_17822, n20718);
  and g38157 (n20719, n20706, n_17822);
  and g38158 (n20720, n_17821, n_17822);
  not g38159 (n_17823, n20719);
  not g38160 (n_17824, n20720);
  and g38161 (n20721, n_17823, n_17824);
  and g38162 (n20722, n_17539, n_17540);
  not g38163 (n_17825, n20722);
  and g38164 (n20723, n_17554, n_17825);
  not g38165 (n_17826, n20721);
  not g38166 (n_17827, n20723);
  and g38167 (n20724, n_17826, n_17827);
  not g38168 (n_17828, n20724);
  and g38169 (n20725, n_17826, n_17828);
  and g38170 (n20726, n_17827, n_17828);
  not g38171 (n_17829, n20725);
  not g38172 (n_17830, n20726);
  and g38173 (n20727, n_17829, n_17830);
  and g38174 (n20728, \b[32] , n9339);
  and g38175 (n20729, \b[30] , n9732);
  and g38176 (n20730, \b[31] , n9334);
  and g38182 (n20733, n4013, n9342);
  not g38185 (n_17835, n20734);
  and g38186 (n20735, \a[53] , n_17835);
  not g38187 (n_17836, n20735);
  and g38188 (n20736, \a[53] , n_17836);
  and g38189 (n20737, n_17835, n_17836);
  not g38190 (n_17837, n20736);
  not g38191 (n_17838, n20737);
  and g38192 (n20738, n_17837, n_17838);
  not g38193 (n_17839, n20727);
  and g38194 (n20739, n_17839, n20738);
  not g38195 (n_17840, n20738);
  and g38196 (n20740, n20727, n_17840);
  not g38197 (n_17841, n20739);
  not g38198 (n_17842, n20740);
  and g38199 (n20741, n_17841, n_17842);
  not g38200 (n_17843, n20664);
  not g38201 (n_17844, n20741);
  and g38202 (n20742, n_17843, n_17844);
  and g38203 (n20743, n20664, n20741);
  not g38204 (n_17845, n20742);
  not g38205 (n_17846, n20743);
  and g38206 (n20744, n_17845, n_17846);
  not g38207 (n_17847, n20663);
  and g38208 (n20745, n_17847, n20744);
  not g38209 (n_17848, n20744);
  and g38210 (n20746, n20663, n_17848);
  not g38211 (n_17849, n20745);
  not g38212 (n_17850, n20746);
  and g38213 (n20747, n_17849, n_17850);
  not g38214 (n_17851, n20652);
  and g38215 (n20748, n_17851, n20747);
  not g38216 (n_17852, n20747);
  and g38217 (n20749, n20652, n_17852);
  not g38218 (n_17853, n20748);
  not g38219 (n_17854, n20749);
  and g38220 (n20750, n_17853, n_17854);
  not g38221 (n_17855, n20651);
  and g38222 (n20751, n_17855, n20750);
  not g38223 (n_17856, n20750);
  and g38224 (n20752, n20651, n_17856);
  not g38225 (n_17857, n20751);
  not g38226 (n_17858, n20752);
  and g38227 (n20753, n_17857, n_17858);
  not g38228 (n_17859, n20640);
  and g38229 (n20754, n_17859, n20753);
  not g38230 (n_17860, n20753);
  and g38231 (n20755, n20640, n_17860);
  not g38232 (n_17861, n20754);
  not g38233 (n_17862, n20755);
  and g38234 (n20756, n_17861, n_17862);
  not g38235 (n_17863, n20639);
  and g38236 (n20757, n_17863, n20756);
  not g38237 (n_17864, n20756);
  and g38238 (n20758, n20639, n_17864);
  not g38239 (n_17865, n20757);
  not g38240 (n_17866, n20758);
  and g38241 (n20759, n_17865, n_17866);
  not g38242 (n_17867, n20628);
  and g38243 (n20760, n_17867, n20759);
  not g38244 (n_17868, n20759);
  and g38245 (n20761, n20628, n_17868);
  not g38246 (n_17869, n20760);
  not g38247 (n_17870, n20761);
  and g38248 (n20762, n_17869, n_17870);
  not g38249 (n_17871, n20627);
  and g38250 (n20763, n_17871, n20762);
  not g38251 (n_17872, n20762);
  and g38252 (n20764, n20627, n_17872);
  not g38253 (n_17873, n20763);
  not g38254 (n_17874, n20764);
  and g38255 (n20765, n_17873, n_17874);
  not g38256 (n_17875, n20616);
  and g38257 (n20766, n_17875, n20765);
  not g38258 (n_17876, n20765);
  and g38259 (n20767, n20616, n_17876);
  not g38260 (n_17877, n20766);
  not g38261 (n_17878, n20767);
  and g38262 (n20768, n_17877, n_17878);
  and g38263 (n20769, \b[47] , n5035);
  and g38264 (n20770, \b[45] , n5277);
  and g38265 (n20771, \b[46] , n5030);
  and g38271 (n20774, n5038, n7703);
  not g38274 (n_17883, n20775);
  and g38275 (n20776, \a[38] , n_17883);
  not g38276 (n_17884, n20776);
  and g38277 (n20777, \a[38] , n_17884);
  and g38278 (n20778, n_17883, n_17884);
  not g38279 (n_17885, n20777);
  not g38280 (n_17886, n20778);
  and g38281 (n20779, n_17885, n_17886);
  not g38282 (n_17887, n20779);
  and g38283 (n20780, n20768, n_17887);
  not g38284 (n_17888, n20780);
  and g38285 (n20781, n20768, n_17888);
  and g38286 (n20782, n_17887, n_17888);
  not g38287 (n_17889, n20781);
  not g38288 (n_17890, n20782);
  and g38289 (n20783, n_17889, n_17890);
  and g38290 (n20784, n_17615, n_17625);
  and g38291 (n20785, n20783, n20784);
  not g38292 (n_17891, n20783);
  not g38293 (n_17892, n20784);
  and g38294 (n20786, n_17891, n_17892);
  not g38295 (n_17893, n20785);
  not g38296 (n_17894, n20786);
  and g38297 (n20787, n_17893, n_17894);
  and g38298 (n20788, \b[50] , n4287);
  and g38299 (n20789, \b[48] , n4532);
  and g38300 (n20790, \b[49] , n4282);
  and g38306 (n20793, n4290, n8949);
  not g38309 (n_17899, n20794);
  and g38310 (n20795, \a[35] , n_17899);
  not g38311 (n_17900, n20795);
  and g38312 (n20796, \a[35] , n_17900);
  and g38313 (n20797, n_17899, n_17900);
  not g38314 (n_17901, n20796);
  not g38315 (n_17902, n20797);
  and g38316 (n20798, n_17901, n_17902);
  not g38317 (n_17903, n20798);
  and g38318 (n20799, n20787, n_17903);
  not g38319 (n_17904, n20787);
  and g38320 (n20800, n_17904, n20798);
  not g38321 (n_17905, n20800);
  and g38322 (n20801, n20615, n_17905);
  not g38323 (n_17906, n20799);
  and g38324 (n20802, n_17906, n20801);
  not g38325 (n_17907, n20802);
  and g38326 (n20803, n20615, n_17907);
  and g38327 (n20804, n_17905, n_17907);
  and g38328 (n20805, n_17906, n20804);
  not g38329 (n_17908, n20803);
  not g38330 (n_17909, n20805);
  and g38331 (n20806, n_17908, n_17909);
  not g38332 (n_17910, n20600);
  and g38333 (n20807, n_17910, n20806);
  not g38334 (n_17911, n20806);
  and g38335 (n20808, n20600, n_17911);
  not g38336 (n_17912, n20807);
  not g38337 (n_17913, n20808);
  and g38338 (n20809, n_17912, n_17913);
  not g38339 (n_17914, n20809);
  and g38340 (n20810, n20584, n_17914);
  not g38341 (n_17915, n20810);
  and g38342 (n20811, n20584, n_17915);
  and g38343 (n20812, n_17914, n_17915);
  not g38344 (n_17916, n20811);
  not g38345 (n_17917, n20812);
  and g38346 (n20813, n_17916, n_17917);
  not g38347 (n_17918, n20569);
  and g38348 (n20814, n_17918, n20813);
  not g38349 (n_17919, n20813);
  and g38350 (n20815, n20569, n_17919);
  not g38351 (n_17920, n20814);
  not g38352 (n_17921, n20815);
  and g38353 (n20816, n_17920, n_17921);
  not g38354 (n_17922, n20553);
  not g38355 (n_17923, n20816);
  and g38356 (n20817, n_17922, n_17923);
  and g38357 (n20818, n20553, n20816);
  not g38358 (n_17924, n20817);
  not g38359 (n_17925, n20818);
  and g38360 (n20819, n_17924, n_17925);
  not g38361 (n_17926, n20541);
  and g38362 (n20820, n_17926, n20819);
  not g38363 (n_17927, n20819);
  and g38364 (n20821, n20541, n_17927);
  not g38365 (n_17928, n20820);
  not g38366 (n_17929, n20821);
  and g38367 (n20822, n_17928, n_17929);
  not g38368 (n_17930, n20540);
  and g38369 (n20823, n_17930, n20822);
  not g38370 (n_17931, n20822);
  and g38371 (n20824, n20540, n_17931);
  not g38372 (n_17932, n20823);
  not g38373 (n_17933, n20824);
  and g38374 (\f[83] , n_17932, n_17933);
  and g38375 (n20826, n_17918, n_17919);
  not g38376 (n_17934, n20826);
  and g38377 (n20827, n_17703, n_17934);
  and g38378 (n20828, \b[63] , n2048);
  and g38379 (n20829, \b[61] , n2198);
  and g38380 (n20830, \b[62] , n2043);
  and g38386 (n20833, n2051, n13771);
  not g38389 (n_17939, n20834);
  and g38390 (n20835, \a[23] , n_17939);
  not g38391 (n_17940, n20835);
  and g38392 (n20836, \a[23] , n_17940);
  and g38393 (n20837, n_17939, n_17940);
  not g38394 (n_17941, n20836);
  not g38395 (n_17942, n20837);
  and g38396 (n20838, n_17941, n_17942);
  not g38397 (n_17943, n20827);
  not g38398 (n_17944, n20838);
  and g38399 (n20839, n_17943, n_17944);
  not g38400 (n_17945, n20839);
  and g38401 (n20840, n_17943, n_17945);
  and g38402 (n20841, n_17944, n_17945);
  not g38403 (n_17946, n20840);
  not g38404 (n_17947, n20841);
  and g38405 (n20842, n_17946, n_17947);
  and g38406 (n20843, \b[60] , n2539);
  and g38407 (n20844, \b[58] , n2685);
  and g38408 (n20845, \b[59] , n2534);
  and g38414 (n20848, n2542, n12211);
  not g38417 (n_17952, n20849);
  and g38418 (n20850, \a[26] , n_17952);
  not g38419 (n_17953, n20850);
  and g38420 (n20851, \a[26] , n_17953);
  and g38421 (n20852, n_17952, n_17953);
  not g38422 (n_17954, n20851);
  not g38423 (n_17955, n20852);
  and g38424 (n20853, n_17954, n_17955);
  and g38425 (n20854, n_17717, n_17915);
  and g38426 (n20855, n20853, n20854);
  not g38427 (n_17956, n20853);
  not g38428 (n_17957, n20854);
  and g38429 (n20856, n_17956, n_17957);
  not g38430 (n_17958, n20855);
  not g38431 (n_17959, n20856);
  and g38432 (n20857, n_17958, n_17959);
  and g38433 (n20858, n_17910, n_17911);
  not g38434 (n_17960, n20858);
  and g38435 (n20859, n_17728, n_17960);
  and g38436 (n20860, \b[57] , n3050);
  and g38437 (n20861, \b[55] , n3243);
  and g38438 (n20862, \b[56] , n3045);
  and g38444 (n20865, n3053, n11410);
  not g38447 (n_17965, n20866);
  and g38448 (n20867, \a[29] , n_17965);
  not g38449 (n_17966, n20867);
  and g38450 (n20868, \a[29] , n_17966);
  and g38451 (n20869, n_17965, n_17966);
  not g38452 (n_17967, n20868);
  not g38453 (n_17968, n20869);
  and g38454 (n20870, n_17967, n_17968);
  not g38455 (n_17969, n20859);
  and g38456 (n20871, n_17969, n20870);
  not g38457 (n_17970, n20870);
  and g38458 (n20872, n20859, n_17970);
  not g38459 (n_17971, n20871);
  not g38460 (n_17972, n20872);
  and g38461 (n20873, n_17971, n_17972);
  and g38462 (n20874, \b[54] , n3638);
  and g38463 (n20875, \b[52] , n3843);
  and g38464 (n20876, \b[53] , n3633);
  and g38470 (n20879, n3641, n9998);
  not g38473 (n_17977, n20880);
  and g38474 (n20881, \a[32] , n_17977);
  not g38475 (n_17978, n20881);
  and g38476 (n20882, \a[32] , n_17978);
  and g38477 (n20883, n_17977, n_17978);
  not g38478 (n_17979, n20882);
  not g38479 (n_17980, n20883);
  and g38480 (n20884, n_17979, n_17980);
  and g38481 (n20885, n_17742, n_17907);
  and g38482 (n20886, n20884, n20885);
  not g38483 (n_17981, n20884);
  not g38484 (n_17982, n20885);
  and g38485 (n20887, n_17981, n_17982);
  not g38486 (n_17983, n20886);
  not g38487 (n_17984, n20887);
  and g38488 (n20888, n_17983, n_17984);
  and g38489 (n20889, n_17894, n_17906);
  and g38490 (n20890, n_17845, n_17849);
  and g38491 (n20891, \b[20] , n13903);
  and g38492 (n20892, \b[21] , n_11555);
  not g38493 (n_17985, n20891);
  not g38494 (n_17986, n20892);
  and g38495 (n20893, n_17985, n_17986);
  not g38496 (n_17987, n20893);
  and g38497 (n20894, n_1221, n_17987);
  and g38498 (n20895, \a[20] , n20893);
  not g38499 (n_17988, n20894);
  not g38500 (n_17989, n20895);
  and g38501 (n20896, n_17988, n_17989);
  and g38502 (n20897, n_17785, n20896);
  not g38503 (n_17990, n20896);
  and g38504 (n20898, n20680, n_17990);
  not g38505 (n_17991, n20897);
  not g38506 (n_17992, n20898);
  and g38507 (n20899, n_17991, n_17992);
  and g38508 (n20900, \b[24] , n12668);
  and g38509 (n20901, \b[22] , n13047);
  and g38510 (n20902, \b[23] , n12663);
  and g38516 (n20905, n2458, n12671);
  not g38519 (n_17997, n20906);
  and g38520 (n20907, \a[62] , n_17997);
  not g38521 (n_17998, n20907);
  and g38522 (n20908, \a[62] , n_17998);
  and g38523 (n20909, n_17997, n_17998);
  not g38524 (n_17999, n20908);
  not g38525 (n_18000, n20909);
  and g38526 (n20910, n_17999, n_18000);
  not g38527 (n_18001, n20910);
  and g38528 (n20911, n20899, n_18001);
  not g38529 (n_18002, n20911);
  and g38530 (n20912, n20899, n_18002);
  and g38531 (n20913, n_18001, n_18002);
  not g38532 (n_18003, n20912);
  not g38533 (n_18004, n20913);
  and g38534 (n20914, n_18003, n_18004);
  and g38535 (n20915, n_17786, n_17799);
  not g38536 (n_18005, n20914);
  not g38537 (n_18006, n20915);
  and g38538 (n20916, n_18005, n_18006);
  not g38539 (n_18007, n20916);
  and g38540 (n20917, n_18005, n_18007);
  and g38541 (n20918, n_18006, n_18007);
  not g38542 (n_18008, n20917);
  not g38543 (n_18009, n20918);
  and g38544 (n20919, n_18008, n_18009);
  and g38545 (n20920, \b[27] , n11531);
  and g38546 (n20921, \b[25] , n11896);
  and g38547 (n20922, \b[26] , n11526);
  and g38553 (n20925, n2990, n11534);
  not g38556 (n_18014, n20926);
  and g38557 (n20927, \a[59] , n_18014);
  not g38558 (n_18015, n20927);
  and g38559 (n20928, \a[59] , n_18015);
  and g38560 (n20929, n_18014, n_18015);
  not g38561 (n_18016, n20928);
  not g38562 (n_18017, n20929);
  and g38563 (n20930, n_18016, n_18017);
  not g38564 (n_18018, n20919);
  not g38565 (n_18019, n20930);
  and g38566 (n20931, n_18018, n_18019);
  not g38567 (n_18020, n20931);
  and g38568 (n20932, n_18018, n_18020);
  and g38569 (n20933, n_18019, n_18020);
  not g38570 (n_18021, n20932);
  not g38571 (n_18022, n20933);
  and g38572 (n20934, n_18021, n_18022);
  and g38573 (n20935, n_17803, n_17807);
  and g38574 (n20936, n20934, n20935);
  not g38575 (n_18023, n20934);
  not g38576 (n_18024, n20935);
  and g38577 (n20937, n_18023, n_18024);
  not g38578 (n_18025, n20936);
  not g38579 (n_18026, n20937);
  and g38580 (n20938, n_18025, n_18026);
  and g38581 (n20939, \b[30] , n10426);
  and g38582 (n20940, \b[28] , n10796);
  and g38583 (n20941, \b[29] , n10421);
  and g38589 (n20944, n3577, n10429);
  not g38592 (n_18031, n20945);
  and g38593 (n20946, \a[56] , n_18031);
  not g38594 (n_18032, n20946);
  and g38595 (n20947, \a[56] , n_18032);
  and g38596 (n20948, n_18031, n_18032);
  not g38597 (n_18033, n20947);
  not g38598 (n_18034, n20948);
  and g38599 (n20949, n_18033, n_18034);
  not g38600 (n_18035, n20949);
  and g38601 (n20950, n20938, n_18035);
  not g38602 (n_18036, n20950);
  and g38603 (n20951, n20938, n_18036);
  and g38604 (n20952, n_18035, n_18036);
  not g38605 (n_18037, n20951);
  not g38606 (n_18038, n20952);
  and g38607 (n20953, n_18037, n_18038);
  and g38608 (n20954, n_17811, n_17822);
  and g38609 (n20955, n20953, n20954);
  not g38610 (n_18039, n20953);
  not g38611 (n_18040, n20954);
  and g38612 (n20956, n_18039, n_18040);
  not g38613 (n_18041, n20955);
  not g38614 (n_18042, n20956);
  and g38615 (n20957, n_18041, n_18042);
  and g38616 (n20958, \b[33] , n9339);
  and g38617 (n20959, \b[31] , n9732);
  and g38618 (n20960, \b[32] , n9334);
  and g38624 (n20963, n4223, n9342);
  not g38627 (n_18047, n20964);
  and g38628 (n20965, \a[53] , n_18047);
  not g38629 (n_18048, n20965);
  and g38630 (n20966, \a[53] , n_18048);
  and g38631 (n20967, n_18047, n_18048);
  not g38632 (n_18049, n20966);
  not g38633 (n_18050, n20967);
  and g38634 (n20968, n_18049, n_18050);
  and g38635 (n20969, n_17839, n_17840);
  not g38636 (n_18051, n20969);
  and g38637 (n20970, n_17828, n_18051);
  not g38638 (n_18052, n20968);
  not g38639 (n_18053, n20970);
  and g38640 (n20971, n_18052, n_18053);
  and g38641 (n20972, n20968, n20970);
  not g38642 (n_18054, n20971);
  not g38643 (n_18055, n20972);
  and g38644 (n20973, n_18054, n_18055);
  not g38645 (n_18056, n20957);
  and g38646 (n20974, n_18056, n20973);
  not g38647 (n_18057, n20973);
  and g38648 (n20975, n20957, n_18057);
  not g38649 (n_18058, n20974);
  not g38650 (n_18059, n20975);
  and g38651 (n20976, n_18058, n_18059);
  and g38652 (n20977, \b[36] , n8362);
  and g38653 (n20978, \b[34] , n8715);
  and g38654 (n20979, \b[35] , n8357);
  and g38660 (n20982, n4922, n8365);
  not g38663 (n_18064, n20983);
  and g38664 (n20984, \a[50] , n_18064);
  not g38665 (n_18065, n20984);
  and g38666 (n20985, \a[50] , n_18065);
  and g38667 (n20986, n_18064, n_18065);
  not g38668 (n_18066, n20985);
  not g38669 (n_18067, n20986);
  and g38670 (n20987, n_18066, n_18067);
  not g38671 (n_18068, n20976);
  not g38672 (n_18069, n20987);
  and g38673 (n20988, n_18068, n_18069);
  and g38674 (n20989, n20976, n20987);
  not g38675 (n_18070, n20988);
  not g38676 (n_18071, n20989);
  and g38677 (n20990, n_18070, n_18071);
  not g38678 (n_18072, n20990);
  and g38679 (n20991, n20890, n_18072);
  not g38680 (n_18073, n20890);
  and g38681 (n20992, n_18073, n20990);
  not g38682 (n_18074, n20991);
  not g38683 (n_18075, n20992);
  and g38684 (n20993, n_18074, n_18075);
  and g38685 (n20994, \b[39] , n7446);
  and g38686 (n20995, \b[37] , n7787);
  and g38687 (n20996, \b[38] , n7441);
  and g38693 (n20999, n5451, n7449);
  not g38696 (n_18080, n21000);
  and g38697 (n21001, \a[47] , n_18080);
  not g38698 (n_18081, n21001);
  and g38699 (n21002, \a[47] , n_18081);
  and g38700 (n21003, n_18080, n_18081);
  not g38701 (n_18082, n21002);
  not g38702 (n_18083, n21003);
  and g38703 (n21004, n_18082, n_18083);
  not g38704 (n_18084, n21004);
  and g38705 (n21005, n20993, n_18084);
  not g38706 (n_18085, n21005);
  and g38707 (n21006, n20993, n_18085);
  and g38708 (n21007, n_18084, n_18085);
  not g38709 (n_18086, n21006);
  not g38710 (n_18087, n21007);
  and g38711 (n21008, n_18086, n_18087);
  and g38712 (n21009, n_17853, n_17857);
  and g38713 (n21010, n21008, n21009);
  not g38714 (n_18088, n21008);
  not g38715 (n_18089, n21009);
  and g38716 (n21011, n_18088, n_18089);
  not g38717 (n_18090, n21010);
  not g38718 (n_18091, n21011);
  and g38719 (n21012, n_18090, n_18091);
  and g38720 (n21013, \b[42] , n6595);
  and g38721 (n21014, \b[40] , n6902);
  and g38722 (n21015, \b[41] , n6590);
  and g38728 (n21018, n6489, n6598);
  not g38731 (n_18096, n21019);
  and g38732 (n21020, \a[44] , n_18096);
  not g38733 (n_18097, n21020);
  and g38734 (n21021, \a[44] , n_18097);
  and g38735 (n21022, n_18096, n_18097);
  not g38736 (n_18098, n21021);
  not g38737 (n_18099, n21022);
  and g38738 (n21023, n_18098, n_18099);
  not g38739 (n_18100, n21023);
  and g38740 (n21024, n21012, n_18100);
  not g38741 (n_18101, n21024);
  and g38742 (n21025, n21012, n_18101);
  and g38743 (n21026, n_18100, n_18101);
  not g38744 (n_18102, n21025);
  not g38745 (n_18103, n21026);
  and g38746 (n21027, n_18102, n_18103);
  and g38747 (n21028, n_17861, n_17865);
  and g38748 (n21029, n21027, n21028);
  not g38749 (n_18104, n21027);
  not g38750 (n_18105, n21028);
  and g38751 (n21030, n_18104, n_18105);
  not g38752 (n_18106, n21029);
  not g38753 (n_18107, n21030);
  and g38754 (n21031, n_18106, n_18107);
  and g38755 (n21032, \b[45] , n5777);
  and g38756 (n21033, \b[43] , n6059);
  and g38757 (n21034, \b[44] , n5772);
  and g38763 (n21037, n5780, n7361);
  not g38766 (n_18112, n21038);
  and g38767 (n21039, \a[41] , n_18112);
  not g38768 (n_18113, n21039);
  and g38769 (n21040, \a[41] , n_18113);
  and g38770 (n21041, n_18112, n_18113);
  not g38771 (n_18114, n21040);
  not g38772 (n_18115, n21041);
  and g38773 (n21042, n_18114, n_18115);
  not g38774 (n_18116, n21042);
  and g38775 (n21043, n21031, n_18116);
  not g38776 (n_18117, n21043);
  and g38777 (n21044, n21031, n_18117);
  and g38778 (n21045, n_18116, n_18117);
  not g38779 (n_18118, n21044);
  not g38780 (n_18119, n21045);
  and g38781 (n21046, n_18118, n_18119);
  and g38782 (n21047, n_17869, n_17873);
  and g38783 (n21048, n21046, n21047);
  not g38784 (n_18120, n21046);
  not g38785 (n_18121, n21047);
  and g38786 (n21049, n_18120, n_18121);
  not g38787 (n_18122, n21048);
  not g38788 (n_18123, n21049);
  and g38789 (n21050, n_18122, n_18123);
  and g38790 (n21051, \b[48] , n5035);
  and g38791 (n21052, \b[46] , n5277);
  and g38792 (n21053, \b[47] , n5030);
  and g38798 (n21056, n5038, n8009);
  not g38801 (n_18128, n21057);
  and g38802 (n21058, \a[38] , n_18128);
  not g38803 (n_18129, n21058);
  and g38804 (n21059, \a[38] , n_18129);
  and g38805 (n21060, n_18128, n_18129);
  not g38806 (n_18130, n21059);
  not g38807 (n_18131, n21060);
  and g38808 (n21061, n_18130, n_18131);
  not g38809 (n_18132, n21061);
  and g38810 (n21062, n21050, n_18132);
  not g38811 (n_18133, n21062);
  and g38812 (n21063, n21050, n_18133);
  and g38813 (n21064, n_18132, n_18133);
  not g38814 (n_18134, n21063);
  not g38815 (n_18135, n21064);
  and g38816 (n21065, n_18134, n_18135);
  and g38817 (n21066, n_17877, n_17888);
  and g38818 (n21067, n21065, n21066);
  not g38819 (n_18136, n21065);
  not g38820 (n_18137, n21066);
  and g38821 (n21068, n_18136, n_18137);
  not g38822 (n_18138, n21067);
  not g38823 (n_18139, n21068);
  and g38824 (n21069, n_18138, n_18139);
  and g38825 (n21070, \b[51] , n4287);
  and g38826 (n21071, \b[49] , n4532);
  and g38827 (n21072, \b[50] , n4282);
  and g38833 (n21075, n4290, n8976);
  not g38836 (n_18144, n21076);
  and g38837 (n21077, \a[35] , n_18144);
  not g38838 (n_18145, n21077);
  and g38839 (n21078, \a[35] , n_18145);
  and g38840 (n21079, n_18144, n_18145);
  not g38841 (n_18146, n21078);
  not g38842 (n_18147, n21079);
  and g38843 (n21080, n_18146, n_18147);
  not g38844 (n_18148, n21080);
  and g38845 (n21081, n21069, n_18148);
  not g38846 (n_18149, n21069);
  and g38847 (n21082, n_18149, n21080);
  not g38848 (n_18150, n20889);
  not g38849 (n_18151, n21082);
  and g38850 (n21083, n_18150, n_18151);
  not g38851 (n_18152, n21081);
  and g38852 (n21084, n_18152, n21083);
  not g38853 (n_18153, n21084);
  and g38854 (n21085, n_18150, n_18153);
  and g38855 (n21086, n_18152, n_18153);
  and g38856 (n21087, n_18151, n21086);
  not g38857 (n_18154, n21085);
  not g38858 (n_18155, n21087);
  and g38859 (n21088, n_18154, n_18155);
  not g38860 (n_18156, n21088);
  and g38861 (n21089, n20888, n_18156);
  not g38862 (n_18157, n20888);
  and g38863 (n21090, n_18157, n21088);
  not g38864 (n_18158, n20873);
  not g38865 (n_18159, n21090);
  and g38866 (n21091, n_18158, n_18159);
  not g38867 (n_18160, n21089);
  and g38868 (n21092, n_18160, n21091);
  not g38869 (n_18161, n21092);
  and g38870 (n21093, n_18158, n_18161);
  and g38871 (n21094, n_18159, n_18161);
  and g38872 (n21095, n_18160, n21094);
  not g38873 (n_18162, n21093);
  not g38874 (n_18163, n21095);
  and g38875 (n21096, n_18162, n_18163);
  not g38876 (n_18164, n21096);
  and g38877 (n21097, n20857, n_18164);
  not g38878 (n_18165, n20857);
  and g38879 (n21098, n_18165, n21096);
  not g38880 (n_18166, n20842);
  not g38881 (n_18167, n21098);
  and g38882 (n21099, n_18166, n_18167);
  not g38883 (n_18168, n21097);
  and g38884 (n21100, n_18168, n21099);
  not g38885 (n_18169, n21100);
  and g38886 (n21101, n_18166, n_18169);
  and g38887 (n21102, n_18167, n_18169);
  and g38888 (n21103, n_18168, n21102);
  not g38889 (n_18170, n21101);
  not g38890 (n_18171, n21103);
  and g38891 (n21104, n_18170, n_18171);
  and g38892 (n21105, n_17690, n_17924);
  and g38893 (n21106, n21104, n21105);
  not g38894 (n_18172, n21104);
  not g38895 (n_18173, n21105);
  and g38896 (n21107, n_18172, n_18173);
  not g38897 (n_18174, n21106);
  not g38898 (n_18175, n21107);
  and g38899 (n21108, n_18174, n_18175);
  and g38900 (n21109, n_17928, n_17932);
  not g38901 (n_18176, n21109);
  and g38902 (n21110, n21108, n_18176);
  not g38903 (n_18177, n21108);
  and g38904 (n21111, n_18177, n21109);
  not g38905 (n_18178, n21110);
  not g38906 (n_18179, n21111);
  and g38907 (\f[84] , n_18178, n_18179);
  and g38908 (n21113, n_17959, n_18168);
  and g38909 (n21114, \b[62] , n2198);
  and g38910 (n21115, \b[63] , n2043);
  not g38911 (n_18180, n21114);
  not g38912 (n_18181, n21115);
  and g38913 (n21116, n_18180, n_18181);
  and g38914 (n21117, n_15432, n21116);
  and g38915 (n21118, n13800, n21116);
  not g38916 (n_18182, n21117);
  not g38917 (n_18183, n21118);
  and g38918 (n21119, n_18182, n_18183);
  not g38919 (n_18184, n21119);
  and g38920 (n21120, \a[23] , n_18184);
  and g38921 (n21121, n_1590, n21119);
  not g38922 (n_18185, n21120);
  not g38923 (n_18186, n21121);
  and g38924 (n21122, n_18185, n_18186);
  not g38925 (n_18187, n21113);
  not g38926 (n_18188, n21122);
  and g38927 (n21123, n_18187, n_18188);
  and g38928 (n21124, n21113, n21122);
  not g38929 (n_18189, n21123);
  not g38930 (n_18190, n21124);
  and g38931 (n21125, n_18189, n_18190);
  and g38932 (n21126, \b[61] , n2539);
  and g38933 (n21127, \b[59] , n2685);
  and g38934 (n21128, \b[60] , n2534);
  and g38940 (n21131, n2542, n12969);
  not g38943 (n_18195, n21132);
  and g38944 (n21133, \a[26] , n_18195);
  not g38945 (n_18196, n21133);
  and g38946 (n21134, \a[26] , n_18196);
  and g38947 (n21135, n_18195, n_18196);
  not g38948 (n_18197, n21134);
  not g38949 (n_18198, n21135);
  and g38950 (n21136, n_18197, n_18198);
  and g38951 (n21137, n_17969, n_17970);
  not g38952 (n_18199, n21137);
  and g38953 (n21138, n_18161, n_18199);
  and g38954 (n21139, n21136, n21138);
  not g38955 (n_18200, n21136);
  not g38956 (n_18201, n21138);
  and g38957 (n21140, n_18200, n_18201);
  not g38958 (n_18202, n21139);
  not g38959 (n_18203, n21140);
  and g38960 (n21141, n_18202, n_18203);
  and g38961 (n21142, n_17984, n_18160);
  and g38962 (n21143, \b[58] , n3050);
  and g38963 (n21144, \b[56] , n3243);
  and g38964 (n21145, \b[57] , n3045);
  not g38965 (n_18204, n21144);
  not g38966 (n_18205, n21145);
  and g38967 (n21146, n_18204, n_18205);
  not g38968 (n_18206, n21143);
  and g38969 (n21147, n_18206, n21146);
  and g38970 (n21148, n_12601, n21147);
  and g38971 (n21149, n_13160, n21147);
  not g38972 (n_18207, n21148);
  not g38973 (n_18208, n21149);
  and g38974 (n21150, n_18207, n_18208);
  not g38975 (n_18209, n21150);
  and g38976 (n21151, \a[29] , n_18209);
  and g38977 (n21152, n_2476, n21150);
  not g38978 (n_18210, n21151);
  not g38979 (n_18211, n21152);
  and g38980 (n21153, n_18210, n_18211);
  not g38981 (n_18212, n21142);
  not g38982 (n_18213, n21153);
  and g38983 (n21154, n_18212, n_18213);
  and g38984 (n21155, n21142, n21153);
  not g38985 (n_18214, n21154);
  not g38986 (n_18215, n21155);
  and g38987 (n21156, n_18214, n_18215);
  and g38988 (n21157, \b[55] , n3638);
  and g38989 (n21158, \b[53] , n3843);
  and g38990 (n21159, \b[54] , n3633);
  and g38996 (n21162, n3641, n10684);
  not g38999 (n_18220, n21163);
  and g39000 (n21164, \a[32] , n_18220);
  not g39001 (n_18221, n21164);
  and g39002 (n21165, \a[32] , n_18221);
  and g39003 (n21166, n_18220, n_18221);
  not g39004 (n_18222, n21165);
  not g39005 (n_18223, n21166);
  and g39006 (n21167, n_18222, n_18223);
  not g39007 (n_18224, n21086);
  and g39008 (n21168, n_18224, n21167);
  not g39009 (n_18225, n21167);
  and g39010 (n21169, n21086, n_18225);
  not g39011 (n_18226, n21168);
  not g39012 (n_18227, n21169);
  and g39013 (n21170, n_18226, n_18227);
  and g39014 (n21171, \b[43] , n6595);
  and g39015 (n21172, \b[41] , n6902);
  and g39016 (n21173, \b[42] , n6590);
  and g39022 (n21176, n6515, n6598);
  not g39025 (n_18232, n21177);
  and g39026 (n21178, \a[44] , n_18232);
  not g39027 (n_18233, n21178);
  and g39028 (n21179, \a[44] , n_18233);
  and g39029 (n21180, n_18232, n_18233);
  not g39030 (n_18234, n21179);
  not g39031 (n_18235, n21180);
  and g39032 (n21181, n_18234, n_18235);
  and g39033 (n21182, n_18085, n_18091);
  and g39034 (n21183, \b[40] , n7446);
  and g39035 (n21184, \b[38] , n7787);
  and g39036 (n21185, \b[39] , n7441);
  and g39042 (n21188, n5955, n7449);
  not g39045 (n_18240, n21189);
  and g39046 (n21190, \a[47] , n_18240);
  not g39047 (n_18241, n21190);
  and g39048 (n21191, \a[47] , n_18241);
  and g39049 (n21192, n_18240, n_18241);
  not g39050 (n_18242, n21191);
  not g39051 (n_18243, n21192);
  and g39052 (n21193, n_18242, n_18243);
  and g39053 (n21194, n_18070, n_18075);
  and g39054 (n21195, n_18020, n_18026);
  and g39055 (n21196, \b[28] , n11531);
  and g39056 (n21197, \b[26] , n11896);
  and g39057 (n21198, \b[27] , n11526);
  and g39063 (n21201, n3189, n11534);
  not g39066 (n_18248, n21202);
  and g39067 (n21203, \a[59] , n_18248);
  not g39068 (n_18249, n21203);
  and g39069 (n21204, \a[59] , n_18249);
  and g39070 (n21205, n_18248, n_18249);
  not g39071 (n_18250, n21204);
  not g39072 (n_18251, n21205);
  and g39073 (n21206, n_18250, n_18251);
  and g39074 (n21207, n_18002, n_18007);
  and g39075 (n21208, \b[21] , n13903);
  and g39076 (n21209, \b[22] , n_11555);
  not g39077 (n_18252, n21208);
  not g39078 (n_18253, n21209);
  and g39079 (n21210, n_18252, n_18253);
  and g39080 (n21211, n_17988, n_17991);
  not g39081 (n_18254, n21210);
  and g39082 (n21212, n_18254, n21211);
  not g39083 (n_18255, n21211);
  and g39084 (n21213, n21210, n_18255);
  not g39085 (n_18256, n21212);
  not g39086 (n_18257, n21213);
  and g39087 (n21214, n_18256, n_18257);
  and g39088 (n21215, \b[25] , n12668);
  and g39089 (n21216, \b[23] , n13047);
  and g39090 (n21217, \b[24] , n12663);
  not g39091 (n_18258, n21216);
  not g39092 (n_18259, n21217);
  and g39093 (n21218, n_18258, n_18259);
  not g39094 (n_18260, n21215);
  and g39095 (n21219, n_18260, n21218);
  and g39096 (n21220, n_12644, n21219);
  not g39097 (n_18261, n2485);
  and g39098 (n21221, n_18261, n21219);
  not g39099 (n_18262, n21220);
  not g39100 (n_18263, n21221);
  and g39101 (n21222, n_18262, n_18263);
  not g39102 (n_18264, n21222);
  and g39103 (n21223, \a[62] , n_18264);
  and g39104 (n21224, n_10843, n21222);
  not g39105 (n_18265, n21223);
  not g39106 (n_18266, n21224);
  and g39107 (n21225, n_18265, n_18266);
  not g39108 (n_18267, n21225);
  and g39109 (n21226, n21214, n_18267);
  not g39110 (n_18268, n21214);
  and g39111 (n21227, n_18268, n21225);
  not g39112 (n_18269, n21226);
  not g39113 (n_18270, n21227);
  and g39114 (n21228, n_18269, n_18270);
  not g39115 (n_18271, n21207);
  and g39116 (n21229, n_18271, n21228);
  not g39117 (n_18272, n21228);
  and g39118 (n21230, n21207, n_18272);
  not g39119 (n_18273, n21229);
  not g39120 (n_18274, n21230);
  and g39121 (n21231, n_18273, n_18274);
  not g39122 (n_18275, n21206);
  and g39123 (n21232, n_18275, n21231);
  not g39124 (n_18276, n21231);
  and g39125 (n21233, n21206, n_18276);
  not g39126 (n_18277, n21232);
  not g39127 (n_18278, n21233);
  and g39128 (n21234, n_18277, n_18278);
  not g39129 (n_18279, n21195);
  and g39130 (n21235, n_18279, n21234);
  not g39131 (n_18280, n21234);
  and g39132 (n21236, n21195, n_18280);
  not g39133 (n_18281, n21235);
  not g39134 (n_18282, n21236);
  and g39135 (n21237, n_18281, n_18282);
  and g39136 (n21238, \b[31] , n10426);
  and g39137 (n21239, \b[29] , n10796);
  and g39138 (n21240, \b[30] , n10421);
  and g39144 (n21243, n3796, n10429);
  not g39147 (n_18287, n21244);
  and g39148 (n21245, \a[56] , n_18287);
  not g39149 (n_18288, n21245);
  and g39150 (n21246, \a[56] , n_18288);
  and g39151 (n21247, n_18287, n_18288);
  not g39152 (n_18289, n21246);
  not g39153 (n_18290, n21247);
  and g39154 (n21248, n_18289, n_18290);
  not g39155 (n_18291, n21248);
  and g39156 (n21249, n21237, n_18291);
  not g39157 (n_18292, n21249);
  and g39158 (n21250, n21237, n_18292);
  and g39159 (n21251, n_18291, n_18292);
  not g39160 (n_18293, n21250);
  not g39161 (n_18294, n21251);
  and g39162 (n21252, n_18293, n_18294);
  and g39163 (n21253, n_18036, n_18042);
  and g39164 (n21254, n21252, n21253);
  not g39165 (n_18295, n21252);
  not g39166 (n_18296, n21253);
  and g39167 (n21255, n_18295, n_18296);
  not g39168 (n_18297, n21254);
  not g39169 (n_18298, n21255);
  and g39170 (n21256, n_18297, n_18298);
  and g39171 (n21257, \b[34] , n9339);
  and g39172 (n21258, \b[32] , n9732);
  and g39173 (n21259, \b[33] , n9334);
  and g39179 (n21262, n4466, n9342);
  not g39182 (n_18303, n21263);
  and g39183 (n21264, \a[53] , n_18303);
  not g39184 (n_18304, n21264);
  and g39185 (n21265, \a[53] , n_18304);
  and g39186 (n21266, n_18303, n_18304);
  not g39187 (n_18305, n21265);
  not g39188 (n_18306, n21266);
  and g39189 (n21267, n_18305, n_18306);
  not g39190 (n_18307, n21267);
  and g39191 (n21268, n21256, n_18307);
  not g39192 (n_18308, n21268);
  and g39193 (n21269, n21256, n_18308);
  and g39194 (n21270, n_18307, n_18308);
  not g39195 (n_18309, n21269);
  not g39196 (n_18310, n21270);
  and g39197 (n21271, n_18309, n_18310);
  and g39198 (n21272, n20957, n20973);
  not g39199 (n_18311, n21272);
  and g39200 (n21273, n_18054, n_18311);
  and g39201 (n21274, n21271, n21273);
  not g39202 (n_18312, n21271);
  not g39203 (n_18313, n21273);
  and g39204 (n21275, n_18312, n_18313);
  not g39205 (n_18314, n21274);
  not g39206 (n_18315, n21275);
  and g39207 (n21276, n_18314, n_18315);
  and g39208 (n21277, \b[37] , n8362);
  and g39209 (n21278, \b[35] , n8715);
  and g39210 (n21279, \b[36] , n8357);
  and g39216 (n21282, n5181, n8365);
  not g39219 (n_18320, n21283);
  and g39220 (n21284, \a[50] , n_18320);
  not g39221 (n_18321, n21284);
  and g39222 (n21285, \a[50] , n_18321);
  and g39223 (n21286, n_18320, n_18321);
  not g39224 (n_18322, n21285);
  not g39225 (n_18323, n21286);
  and g39226 (n21287, n_18322, n_18323);
  not g39227 (n_18324, n21276);
  and g39228 (n21288, n_18324, n21287);
  not g39229 (n_18325, n21287);
  and g39230 (n21289, n21276, n_18325);
  not g39231 (n_18326, n21288);
  not g39232 (n_18327, n21289);
  and g39233 (n21290, n_18326, n_18327);
  not g39234 (n_18328, n21194);
  and g39235 (n21291, n_18328, n21290);
  not g39236 (n_18329, n21291);
  and g39237 (n21292, n_18328, n_18329);
  and g39238 (n21293, n21290, n_18329);
  not g39239 (n_18330, n21292);
  not g39240 (n_18331, n21293);
  and g39241 (n21294, n_18330, n_18331);
  not g39242 (n_18332, n21193);
  not g39243 (n_18333, n21294);
  and g39244 (n21295, n_18332, n_18333);
  and g39245 (n21296, n21193, n_18331);
  and g39246 (n21297, n_18330, n21296);
  not g39247 (n_18334, n21295);
  not g39248 (n_18335, n21297);
  and g39249 (n21298, n_18334, n_18335);
  not g39250 (n_18336, n21182);
  and g39251 (n21299, n_18336, n21298);
  not g39252 (n_18337, n21298);
  and g39253 (n21300, n21182, n_18337);
  not g39254 (n_18338, n21299);
  not g39255 (n_18339, n21300);
  and g39256 (n21301, n_18338, n_18339);
  not g39257 (n_18340, n21181);
  and g39258 (n21302, n_18340, n21301);
  not g39259 (n_18341, n21302);
  and g39260 (n21303, n21301, n_18341);
  and g39261 (n21304, n_18340, n_18341);
  not g39262 (n_18342, n21303);
  not g39263 (n_18343, n21304);
  and g39264 (n21305, n_18342, n_18343);
  and g39265 (n21306, n_18101, n_18107);
  and g39266 (n21307, n21305, n21306);
  not g39267 (n_18344, n21305);
  not g39268 (n_18345, n21306);
  and g39269 (n21308, n_18344, n_18345);
  not g39270 (n_18346, n21307);
  not g39271 (n_18347, n21308);
  and g39272 (n21309, n_18346, n_18347);
  and g39273 (n21310, \b[46] , n5777);
  and g39274 (n21311, \b[44] , n6059);
  and g39275 (n21312, \b[45] , n5772);
  and g39281 (n21315, n5780, n7677);
  not g39284 (n_18352, n21316);
  and g39285 (n21317, \a[41] , n_18352);
  not g39286 (n_18353, n21317);
  and g39287 (n21318, \a[41] , n_18353);
  and g39288 (n21319, n_18352, n_18353);
  not g39289 (n_18354, n21318);
  not g39290 (n_18355, n21319);
  and g39291 (n21320, n_18354, n_18355);
  not g39292 (n_18356, n21320);
  and g39293 (n21321, n21309, n_18356);
  not g39294 (n_18357, n21321);
  and g39295 (n21322, n21309, n_18357);
  and g39296 (n21323, n_18356, n_18357);
  not g39297 (n_18358, n21322);
  not g39298 (n_18359, n21323);
  and g39299 (n21324, n_18358, n_18359);
  and g39300 (n21325, n_18117, n_18123);
  and g39301 (n21326, n21324, n21325);
  not g39302 (n_18360, n21324);
  not g39303 (n_18361, n21325);
  and g39304 (n21327, n_18360, n_18361);
  not g39305 (n_18362, n21326);
  not g39306 (n_18363, n21327);
  and g39307 (n21328, n_18362, n_18363);
  and g39308 (n21329, \b[49] , n5035);
  and g39309 (n21330, \b[47] , n5277);
  and g39310 (n21331, \b[48] , n5030);
  and g39316 (n21334, n5038, n8625);
  not g39319 (n_18368, n21335);
  and g39320 (n21336, \a[38] , n_18368);
  not g39321 (n_18369, n21336);
  and g39322 (n21337, \a[38] , n_18369);
  and g39323 (n21338, n_18368, n_18369);
  not g39324 (n_18370, n21337);
  not g39325 (n_18371, n21338);
  and g39326 (n21339, n_18370, n_18371);
  not g39327 (n_18372, n21339);
  and g39328 (n21340, n21328, n_18372);
  not g39329 (n_18373, n21340);
  and g39330 (n21341, n21328, n_18373);
  and g39331 (n21342, n_18372, n_18373);
  not g39332 (n_18374, n21341);
  not g39333 (n_18375, n21342);
  and g39334 (n21343, n_18374, n_18375);
  and g39335 (n21344, n_18133, n_18139);
  and g39336 (n21345, n21343, n21344);
  not g39337 (n_18376, n21343);
  not g39338 (n_18377, n21344);
  and g39339 (n21346, n_18376, n_18377);
  not g39340 (n_18378, n21345);
  not g39341 (n_18379, n21346);
  and g39342 (n21347, n_18378, n_18379);
  and g39343 (n21348, \b[52] , n4287);
  and g39344 (n21349, \b[50] , n4532);
  and g39345 (n21350, \b[51] , n4282);
  and g39351 (n21353, n4290, n9628);
  not g39354 (n_18384, n21354);
  and g39355 (n21355, \a[35] , n_18384);
  not g39356 (n_18385, n21355);
  and g39357 (n21356, \a[35] , n_18385);
  and g39358 (n21357, n_18384, n_18385);
  not g39359 (n_18386, n21356);
  not g39360 (n_18387, n21357);
  and g39361 (n21358, n_18386, n_18387);
  not g39362 (n_18388, n21358);
  and g39363 (n21359, n21347, n_18388);
  not g39364 (n_18389, n21359);
  and g39365 (n21360, n21347, n_18389);
  and g39366 (n21361, n_18388, n_18389);
  not g39367 (n_18390, n21360);
  not g39368 (n_18391, n21361);
  and g39369 (n21362, n_18390, n_18391);
  not g39370 (n_18392, n21170);
  not g39371 (n_18393, n21362);
  and g39372 (n21363, n_18392, n_18393);
  and g39373 (n21364, n21170, n21362);
  not g39374 (n_18394, n21364);
  and g39375 (n21365, n21156, n_18394);
  not g39376 (n_18395, n21363);
  and g39377 (n21366, n_18395, n21365);
  not g39378 (n_18396, n21366);
  and g39379 (n21367, n21156, n_18396);
  and g39380 (n21368, n_18394, n_18396);
  and g39381 (n21369, n_18395, n21368);
  not g39382 (n_18397, n21367);
  not g39383 (n_18398, n21369);
  and g39384 (n21370, n_18397, n_18398);
  not g39385 (n_18399, n21370);
  and g39386 (n21371, n21141, n_18399);
  not g39387 (n_18400, n21141);
  and g39388 (n21372, n_18400, n21370);
  not g39389 (n_18401, n21372);
  and g39390 (n21373, n21125, n_18401);
  not g39391 (n_18402, n21371);
  and g39392 (n21374, n_18402, n21373);
  not g39393 (n_18403, n21374);
  and g39394 (n21375, n21125, n_18403);
  and g39395 (n21376, n_18401, n_18403);
  and g39396 (n21377, n_18402, n21376);
  not g39397 (n_18404, n21375);
  not g39398 (n_18405, n21377);
  and g39399 (n21378, n_18404, n_18405);
  and g39400 (n21379, n_17945, n_18169);
  and g39401 (n21380, n21378, n21379);
  not g39402 (n_18406, n21378);
  not g39403 (n_18407, n21379);
  and g39404 (n21381, n_18406, n_18407);
  not g39405 (n_18408, n21380);
  not g39406 (n_18409, n21381);
  and g39407 (n21382, n_18408, n_18409);
  and g39408 (n21383, n_18175, n_18178);
  not g39409 (n_18410, n21383);
  and g39410 (n21384, n21382, n_18410);
  not g39411 (n_18411, n21382);
  and g39412 (n21385, n_18411, n21383);
  not g39413 (n_18412, n21384);
  not g39414 (n_18413, n21385);
  and g39415 (\f[85] , n_18412, n_18413);
  and g39416 (n21387, n_18409, n_18412);
  and g39417 (n21388, n_18189, n_18403);
  and g39418 (n21389, n_18203, n_18402);
  and g39419 (n21390, \b[63] , n2198);
  and g39420 (n21391, n2051, n13797);
  not g39421 (n_18414, n21390);
  not g39422 (n_18415, n21391);
  and g39423 (n21392, n_18414, n_18415);
  not g39424 (n_18416, n21392);
  and g39425 (n21393, \a[23] , n_18416);
  not g39426 (n_18417, n21393);
  and g39427 (n21394, \a[23] , n_18417);
  and g39428 (n21395, n_18416, n_18417);
  not g39429 (n_18418, n21394);
  not g39430 (n_18419, n21395);
  and g39431 (n21396, n_18418, n_18419);
  not g39432 (n_18420, n21389);
  not g39433 (n_18421, n21396);
  and g39434 (n21397, n_18420, n_18421);
  not g39435 (n_18422, n21397);
  and g39436 (n21398, n_18420, n_18422);
  and g39437 (n21399, n_18421, n_18422);
  not g39438 (n_18423, n21398);
  not g39439 (n_18424, n21399);
  and g39440 (n21400, n_18423, n_18424);
  and g39441 (n21401, \b[62] , n2539);
  and g39442 (n21402, \b[60] , n2685);
  and g39443 (n21403, \b[61] , n2534);
  and g39449 (n21406, n2542, n13370);
  not g39452 (n_18429, n21407);
  and g39453 (n21408, \a[26] , n_18429);
  not g39454 (n_18430, n21408);
  and g39455 (n21409, \a[26] , n_18430);
  and g39456 (n21410, n_18429, n_18430);
  not g39457 (n_18431, n21409);
  not g39458 (n_18432, n21410);
  and g39459 (n21411, n_18431, n_18432);
  and g39460 (n21412, n_18214, n_18396);
  and g39461 (n21413, n21411, n21412);
  not g39462 (n_18433, n21411);
  not g39463 (n_18434, n21412);
  and g39464 (n21414, n_18433, n_18434);
  not g39465 (n_18435, n21413);
  not g39466 (n_18436, n21414);
  and g39467 (n21415, n_18435, n_18436);
  and g39468 (n21416, \b[59] , n3050);
  and g39469 (n21417, \b[57] , n3243);
  and g39470 (n21418, \b[58] , n3045);
  and g39476 (n21421, n3053, n12179);
  not g39479 (n_18441, n21422);
  and g39480 (n21423, \a[29] , n_18441);
  not g39481 (n_18442, n21423);
  and g39482 (n21424, \a[29] , n_18442);
  and g39483 (n21425, n_18441, n_18442);
  not g39484 (n_18443, n21424);
  not g39485 (n_18444, n21425);
  and g39486 (n21426, n_18443, n_18444);
  and g39487 (n21427, n_18224, n_18225);
  not g39488 (n_18445, n21427);
  and g39489 (n21428, n_18395, n_18445);
  not g39490 (n_18446, n21426);
  not g39491 (n_18447, n21428);
  and g39492 (n21429, n_18446, n_18447);
  not g39493 (n_18448, n21429);
  and g39494 (n21430, n_18446, n_18448);
  and g39495 (n21431, n_18447, n_18448);
  not g39496 (n_18449, n21430);
  not g39497 (n_18450, n21431);
  and g39498 (n21432, n_18449, n_18450);
  and g39499 (n21433, \b[56] , n3638);
  and g39500 (n21434, \b[54] , n3843);
  and g39501 (n21435, \b[55] , n3633);
  and g39507 (n21438, n3641, n10708);
  not g39510 (n_18455, n21439);
  and g39511 (n21440, \a[32] , n_18455);
  not g39512 (n_18456, n21440);
  and g39513 (n21441, \a[32] , n_18456);
  and g39514 (n21442, n_18455, n_18456);
  not g39515 (n_18457, n21441);
  not g39516 (n_18458, n21442);
  and g39517 (n21443, n_18457, n_18458);
  and g39518 (n21444, n_18379, n_18389);
  and g39519 (n21445, n21443, n21444);
  not g39520 (n_18459, n21443);
  not g39521 (n_18460, n21444);
  and g39522 (n21446, n_18459, n_18460);
  not g39523 (n_18461, n21445);
  not g39524 (n_18462, n21446);
  and g39525 (n21447, n_18461, n_18462);
  and g39526 (n21448, \b[53] , n4287);
  and g39527 (n21449, \b[51] , n4532);
  and g39528 (n21450, \b[52] , n4282);
  and g39534 (n21453, n4290, n9972);
  not g39537 (n_18467, n21454);
  and g39538 (n21455, \a[35] , n_18467);
  not g39539 (n_18468, n21455);
  and g39540 (n21456, \a[35] , n_18468);
  and g39541 (n21457, n_18467, n_18468);
  not g39542 (n_18469, n21456);
  not g39543 (n_18470, n21457);
  and g39544 (n21458, n_18469, n_18470);
  and g39545 (n21459, n_18363, n_18373);
  and g39546 (n21460, n_18338, n_18341);
  and g39547 (n21461, \b[44] , n6595);
  and g39548 (n21462, \b[42] , n6902);
  and g39549 (n21463, \b[43] , n6590);
  and g39555 (n21466, n6598, n7072);
  not g39558 (n_18475, n21467);
  and g39559 (n21468, \a[44] , n_18475);
  not g39560 (n_18476, n21468);
  and g39561 (n21469, \a[44] , n_18476);
  and g39562 (n21470, n_18475, n_18476);
  not g39563 (n_18477, n21469);
  not g39564 (n_18478, n21470);
  and g39565 (n21471, n_18477, n_18478);
  and g39566 (n21472, n_18329, n_18334);
  and g39567 (n21473, n_18298, n_18308);
  and g39568 (n21474, \b[35] , n9339);
  and g39569 (n21475, \b[33] , n9732);
  and g39570 (n21476, \b[34] , n9334);
  and g39576 (n21479, n4696, n9342);
  not g39579 (n_18483, n21480);
  and g39580 (n21481, \a[53] , n_18483);
  not g39581 (n_18484, n21481);
  and g39582 (n21482, \a[53] , n_18484);
  and g39583 (n21483, n_18483, n_18484);
  not g39584 (n_18485, n21482);
  not g39585 (n_18486, n21483);
  and g39586 (n21484, n_18485, n_18486);
  and g39587 (n21485, n_18281, n_18292);
  and g39588 (n21486, n_18257, n_18269);
  and g39589 (n21487, \b[22] , n13903);
  and g39590 (n21488, \b[23] , n_11555);
  not g39591 (n_18487, n21487);
  not g39592 (n_18488, n21488);
  and g39593 (n21489, n_18487, n_18488);
  and g39594 (n21490, n_18254, n21489);
  not g39595 (n_18489, n21489);
  and g39596 (n21491, n21210, n_18489);
  not g39597 (n_18490, n21490);
  not g39598 (n_18491, n21491);
  and g39599 (n21492, n_18490, n_18491);
  and g39600 (n21493, \b[26] , n12668);
  and g39601 (n21494, \b[24] , n13047);
  and g39602 (n21495, \b[25] , n12663);
  not g39603 (n_18492, n21494);
  not g39604 (n_18493, n21495);
  and g39605 (n21496, n_18492, n_18493);
  not g39606 (n_18494, n21493);
  and g39607 (n21497, n_18494, n21496);
  and g39608 (n21498, n_12644, n21497);
  not g39609 (n_18495, n2813);
  and g39610 (n21499, n_18495, n21497);
  not g39611 (n_18496, n21498);
  not g39612 (n_18497, n21499);
  and g39613 (n21500, n_18496, n_18497);
  not g39614 (n_18498, n21500);
  and g39615 (n21501, \a[62] , n_18498);
  and g39616 (n21502, n_10843, n21500);
  not g39617 (n_18499, n21501);
  not g39618 (n_18500, n21502);
  and g39619 (n21503, n_18499, n_18500);
  not g39620 (n_18501, n21503);
  and g39621 (n21504, n21492, n_18501);
  not g39622 (n_18502, n21492);
  and g39623 (n21505, n_18502, n21503);
  not g39624 (n_18503, n21504);
  not g39625 (n_18504, n21505);
  and g39626 (n21506, n_18503, n_18504);
  not g39627 (n_18505, n21486);
  and g39628 (n21507, n_18505, n21506);
  not g39629 (n_18506, n21506);
  and g39630 (n21508, n21486, n_18506);
  not g39631 (n_18507, n21507);
  not g39632 (n_18508, n21508);
  and g39633 (n21509, n_18507, n_18508);
  and g39634 (n21510, \b[29] , n11531);
  and g39635 (n21511, \b[27] , n11896);
  and g39636 (n21512, \b[28] , n11526);
  and g39642 (n21515, n3383, n11534);
  not g39645 (n_18513, n21516);
  and g39646 (n21517, \a[59] , n_18513);
  not g39647 (n_18514, n21517);
  and g39648 (n21518, \a[59] , n_18514);
  and g39649 (n21519, n_18513, n_18514);
  not g39650 (n_18515, n21518);
  not g39651 (n_18516, n21519);
  and g39652 (n21520, n_18515, n_18516);
  not g39653 (n_18517, n21520);
  and g39654 (n21521, n21509, n_18517);
  not g39655 (n_18518, n21521);
  and g39656 (n21522, n21509, n_18518);
  and g39657 (n21523, n_18517, n_18518);
  not g39658 (n_18519, n21522);
  not g39659 (n_18520, n21523);
  and g39660 (n21524, n_18519, n_18520);
  and g39661 (n21525, n_18273, n_18277);
  and g39662 (n21526, n21524, n21525);
  not g39663 (n_18521, n21524);
  not g39664 (n_18522, n21525);
  and g39665 (n21527, n_18521, n_18522);
  not g39666 (n_18523, n21526);
  not g39667 (n_18524, n21527);
  and g39668 (n21528, n_18523, n_18524);
  and g39669 (n21529, \b[32] , n10426);
  and g39670 (n21530, \b[30] , n10796);
  and g39671 (n21531, \b[31] , n10421);
  and g39677 (n21534, n4013, n10429);
  not g39680 (n_18529, n21535);
  and g39681 (n21536, \a[56] , n_18529);
  not g39682 (n_18530, n21536);
  and g39683 (n21537, \a[56] , n_18530);
  and g39684 (n21538, n_18529, n_18530);
  not g39685 (n_18531, n21537);
  not g39686 (n_18532, n21538);
  and g39687 (n21539, n_18531, n_18532);
  not g39688 (n_18533, n21528);
  and g39689 (n21540, n_18533, n21539);
  not g39690 (n_18534, n21539);
  and g39691 (n21541, n21528, n_18534);
  not g39692 (n_18535, n21540);
  not g39693 (n_18536, n21541);
  and g39694 (n21542, n_18535, n_18536);
  not g39695 (n_18537, n21485);
  and g39696 (n21543, n_18537, n21542);
  not g39697 (n_18538, n21542);
  and g39698 (n21544, n21485, n_18538);
  not g39699 (n_18539, n21543);
  not g39700 (n_18540, n21544);
  and g39701 (n21545, n_18539, n_18540);
  not g39702 (n_18541, n21484);
  and g39703 (n21546, n_18541, n21545);
  not g39704 (n_18542, n21545);
  and g39705 (n21547, n21484, n_18542);
  not g39706 (n_18543, n21546);
  not g39707 (n_18544, n21547);
  and g39708 (n21548, n_18543, n_18544);
  not g39709 (n_18545, n21473);
  and g39710 (n21549, n_18545, n21548);
  not g39711 (n_18546, n21548);
  and g39712 (n21550, n21473, n_18546);
  not g39713 (n_18547, n21549);
  not g39714 (n_18548, n21550);
  and g39715 (n21551, n_18547, n_18548);
  and g39716 (n21552, \b[38] , n8362);
  and g39717 (n21553, \b[36] , n8715);
  and g39718 (n21554, \b[37] , n8357);
  and g39724 (n21557, n5205, n8365);
  not g39727 (n_18553, n21558);
  and g39728 (n21559, \a[50] , n_18553);
  not g39729 (n_18554, n21559);
  and g39730 (n21560, \a[50] , n_18554);
  and g39731 (n21561, n_18553, n_18554);
  not g39732 (n_18555, n21560);
  not g39733 (n_18556, n21561);
  and g39734 (n21562, n_18555, n_18556);
  not g39735 (n_18557, n21562);
  and g39736 (n21563, n21551, n_18557);
  not g39737 (n_18558, n21563);
  and g39738 (n21564, n21551, n_18558);
  and g39739 (n21565, n_18557, n_18558);
  not g39740 (n_18559, n21564);
  not g39741 (n_18560, n21565);
  and g39742 (n21566, n_18559, n_18560);
  and g39743 (n21567, n_18315, n_18327);
  not g39744 (n_18561, n21566);
  not g39745 (n_18562, n21567);
  and g39746 (n21568, n_18561, n_18562);
  not g39747 (n_18563, n21568);
  and g39748 (n21569, n_18561, n_18563);
  and g39749 (n21570, n_18562, n_18563);
  not g39750 (n_18564, n21569);
  not g39751 (n_18565, n21570);
  and g39752 (n21571, n_18564, n_18565);
  and g39753 (n21572, \b[41] , n7446);
  and g39754 (n21573, \b[39] , n7787);
  and g39755 (n21574, \b[40] , n7441);
  and g39761 (n21577, n6219, n7449);
  not g39764 (n_18570, n21578);
  and g39765 (n21579, \a[47] , n_18570);
  not g39766 (n_18571, n21579);
  and g39767 (n21580, \a[47] , n_18571);
  and g39768 (n21581, n_18570, n_18571);
  not g39769 (n_18572, n21580);
  not g39770 (n_18573, n21581);
  and g39771 (n21582, n_18572, n_18573);
  not g39772 (n_18574, n21571);
  and g39773 (n21583, n_18574, n21582);
  not g39774 (n_18575, n21582);
  and g39775 (n21584, n21571, n_18575);
  not g39776 (n_18576, n21583);
  not g39777 (n_18577, n21584);
  and g39778 (n21585, n_18576, n_18577);
  not g39779 (n_18578, n21472);
  not g39780 (n_18579, n21585);
  and g39781 (n21586, n_18578, n_18579);
  and g39782 (n21587, n21472, n21585);
  not g39783 (n_18580, n21586);
  not g39784 (n_18581, n21587);
  and g39785 (n21588, n_18580, n_18581);
  not g39786 (n_18582, n21471);
  and g39787 (n21589, n_18582, n21588);
  not g39788 (n_18583, n21588);
  and g39789 (n21590, n21471, n_18583);
  not g39790 (n_18584, n21589);
  not g39791 (n_18585, n21590);
  and g39792 (n21591, n_18584, n_18585);
  not g39793 (n_18586, n21460);
  and g39794 (n21592, n_18586, n21591);
  not g39795 (n_18587, n21591);
  and g39796 (n21593, n21460, n_18587);
  not g39797 (n_18588, n21592);
  not g39798 (n_18589, n21593);
  and g39799 (n21594, n_18588, n_18589);
  and g39800 (n21595, \b[47] , n5777);
  and g39801 (n21596, \b[45] , n6059);
  and g39802 (n21597, \b[46] , n5772);
  and g39808 (n21600, n5780, n7703);
  not g39811 (n_18594, n21601);
  and g39812 (n21602, \a[41] , n_18594);
  not g39813 (n_18595, n21602);
  and g39814 (n21603, \a[41] , n_18595);
  and g39815 (n21604, n_18594, n_18595);
  not g39816 (n_18596, n21603);
  not g39817 (n_18597, n21604);
  and g39818 (n21605, n_18596, n_18597);
  not g39819 (n_18598, n21605);
  and g39820 (n21606, n21594, n_18598);
  not g39821 (n_18599, n21606);
  and g39822 (n21607, n21594, n_18599);
  and g39823 (n21608, n_18598, n_18599);
  not g39824 (n_18600, n21607);
  not g39825 (n_18601, n21608);
  and g39826 (n21609, n_18600, n_18601);
  and g39827 (n21610, n_18347, n_18357);
  and g39828 (n21611, n21609, n21610);
  not g39829 (n_18602, n21609);
  not g39830 (n_18603, n21610);
  and g39831 (n21612, n_18602, n_18603);
  not g39832 (n_18604, n21611);
  not g39833 (n_18605, n21612);
  and g39834 (n21613, n_18604, n_18605);
  and g39835 (n21614, \b[50] , n5035);
  and g39836 (n21615, \b[48] , n5277);
  and g39837 (n21616, \b[49] , n5030);
  and g39843 (n21619, n5038, n8949);
  not g39846 (n_18610, n21620);
  and g39847 (n21621, \a[38] , n_18610);
  not g39848 (n_18611, n21621);
  and g39849 (n21622, \a[38] , n_18611);
  and g39850 (n21623, n_18610, n_18611);
  not g39851 (n_18612, n21622);
  not g39852 (n_18613, n21623);
  and g39853 (n21624, n_18612, n_18613);
  not g39854 (n_18614, n21613);
  and g39855 (n21625, n_18614, n21624);
  not g39856 (n_18615, n21624);
  and g39857 (n21626, n21613, n_18615);
  not g39858 (n_18616, n21625);
  not g39859 (n_18617, n21626);
  and g39860 (n21627, n_18616, n_18617);
  not g39861 (n_18618, n21459);
  and g39862 (n21628, n_18618, n21627);
  not g39863 (n_18619, n21628);
  and g39864 (n21629, n_18618, n_18619);
  and g39865 (n21630, n21627, n_18619);
  not g39866 (n_18620, n21629);
  not g39867 (n_18621, n21630);
  and g39868 (n21631, n_18620, n_18621);
  not g39869 (n_18622, n21458);
  not g39870 (n_18623, n21631);
  and g39871 (n21632, n_18622, n_18623);
  not g39872 (n_18624, n21632);
  and g39873 (n21633, n_18622, n_18624);
  and g39874 (n21634, n_18623, n_18624);
  not g39875 (n_18625, n21633);
  not g39876 (n_18626, n21634);
  and g39877 (n21635, n_18625, n_18626);
  not g39878 (n_18627, n21635);
  and g39879 (n21636, n21447, n_18627);
  not g39880 (n_18628, n21636);
  and g39881 (n21637, n21447, n_18628);
  and g39882 (n21638, n_18627, n_18628);
  not g39883 (n_18629, n21637);
  not g39884 (n_18630, n21638);
  and g39885 (n21639, n_18629, n_18630);
  not g39886 (n_18631, n21432);
  and g39887 (n21640, n_18631, n21639);
  not g39888 (n_18632, n21639);
  and g39889 (n21641, n21432, n_18632);
  not g39890 (n_18633, n21640);
  not g39891 (n_18634, n21641);
  and g39892 (n21642, n_18633, n_18634);
  not g39893 (n_18635, n21642);
  and g39894 (n21643, n21415, n_18635);
  not g39895 (n_18636, n21643);
  and g39896 (n21644, n21415, n_18636);
  and g39897 (n21645, n_18635, n_18636);
  not g39898 (n_18637, n21644);
  not g39899 (n_18638, n21645);
  and g39900 (n21646, n_18637, n_18638);
  not g39901 (n_18639, n21400);
  and g39902 (n21647, n_18639, n21646);
  not g39903 (n_18640, n21646);
  and g39904 (n21648, n21400, n_18640);
  not g39905 (n_18641, n21647);
  not g39906 (n_18642, n21648);
  and g39907 (n21649, n_18641, n_18642);
  not g39908 (n_18643, n21388);
  not g39909 (n_18644, n21649);
  and g39910 (n21650, n_18643, n_18644);
  not g39911 (n_18645, n21650);
  and g39912 (n21651, n_18643, n_18645);
  and g39913 (n21652, n_18644, n_18645);
  not g39914 (n_18646, n21651);
  not g39915 (n_18647, n21652);
  and g39916 (n21653, n_18646, n_18647);
  not g39917 (n_18648, n21387);
  not g39918 (n_18649, n21653);
  and g39919 (n21654, n_18648, n_18649);
  and g39920 (n21655, n21387, n_18647);
  and g39921 (n21656, n_18646, n21655);
  not g39922 (n_18650, n21654);
  not g39923 (n_18651, n21656);
  and g39924 (\f[86] , n_18650, n_18651);
  and g39925 (n21658, n_18645, n_18650);
  and g39926 (n21659, n_18639, n_18640);
  not g39927 (n_18652, n21659);
  and g39928 (n21660, n_18422, n_18652);
  and g39929 (n21661, n_18436, n_18636);
  and g39930 (n21662, \b[63] , n2539);
  and g39931 (n21663, \b[61] , n2685);
  and g39932 (n21664, \b[62] , n2534);
  and g39938 (n21667, n2542, n13771);
  not g39941 (n_18657, n21668);
  and g39942 (n21669, \a[26] , n_18657);
  not g39943 (n_18658, n21669);
  and g39944 (n21670, \a[26] , n_18658);
  and g39945 (n21671, n_18657, n_18658);
  not g39946 (n_18659, n21670);
  not g39947 (n_18660, n21671);
  and g39948 (n21672, n_18659, n_18660);
  not g39949 (n_18661, n21661);
  not g39950 (n_18662, n21672);
  and g39951 (n21673, n_18661, n_18662);
  not g39952 (n_18663, n21673);
  and g39953 (n21674, n_18661, n_18663);
  and g39954 (n21675, n_18662, n_18663);
  not g39955 (n_18664, n21674);
  not g39956 (n_18665, n21675);
  and g39957 (n21676, n_18664, n_18665);
  and g39958 (n21677, n_18631, n_18632);
  not g39959 (n_18666, n21677);
  and g39960 (n21678, n_18448, n_18666);
  and g39961 (n21679, \b[60] , n3050);
  and g39962 (n21680, \b[58] , n3243);
  and g39963 (n21681, \b[59] , n3045);
  and g39969 (n21684, n3053, n12211);
  not g39972 (n_18671, n21685);
  and g39973 (n21686, \a[29] , n_18671);
  not g39974 (n_18672, n21686);
  and g39975 (n21687, \a[29] , n_18672);
  and g39976 (n21688, n_18671, n_18672);
  not g39977 (n_18673, n21687);
  not g39978 (n_18674, n21688);
  and g39979 (n21689, n_18673, n_18674);
  not g39980 (n_18675, n21678);
  and g39981 (n21690, n_18675, n21689);
  not g39982 (n_18676, n21689);
  and g39983 (n21691, n21678, n_18676);
  not g39984 (n_18677, n21690);
  not g39985 (n_18678, n21691);
  and g39986 (n21692, n_18677, n_18678);
  and g39987 (n21693, \b[57] , n3638);
  and g39988 (n21694, \b[55] , n3843);
  and g39989 (n21695, \b[56] , n3633);
  and g39995 (n21698, n3641, n11410);
  not g39998 (n_18683, n21699);
  and g39999 (n21700, \a[32] , n_18683);
  not g40000 (n_18684, n21700);
  and g40001 (n21701, \a[32] , n_18684);
  and g40002 (n21702, n_18683, n_18684);
  not g40003 (n_18685, n21701);
  not g40004 (n_18686, n21702);
  and g40005 (n21703, n_18685, n_18686);
  and g40006 (n21704, n_18462, n_18628);
  and g40007 (n21705, n21703, n21704);
  not g40008 (n_18687, n21703);
  not g40009 (n_18688, n21704);
  and g40010 (n21706, n_18687, n_18688);
  not g40011 (n_18689, n21705);
  not g40012 (n_18690, n21706);
  and g40013 (n21707, n_18689, n_18690);
  and g40014 (n21708, n_18619, n_18624);
  and g40015 (n21709, n_18605, n_18617);
  and g40016 (n21710, n_18580, n_18584);
  and g40017 (n21711, n_18574, n_18575);
  not g40018 (n_18691, n21711);
  and g40019 (n21712, n_18563, n_18691);
  and g40020 (n21713, \b[36] , n9339);
  and g40021 (n21714, \b[34] , n9732);
  and g40022 (n21715, \b[35] , n9334);
  and g40028 (n21718, n4922, n9342);
  not g40031 (n_18696, n21719);
  and g40032 (n21720, \a[53] , n_18696);
  not g40033 (n_18697, n21720);
  and g40034 (n21721, \a[53] , n_18697);
  and g40035 (n21722, n_18696, n_18697);
  not g40036 (n_18698, n21721);
  not g40037 (n_18699, n21722);
  and g40038 (n21723, n_18698, n_18699);
  and g40039 (n21724, n_18507, n_18518);
  and g40040 (n21725, n_18490, n_18503);
  and g40041 (n21726, \b[23] , n13903);
  and g40042 (n21727, \b[24] , n_11555);
  not g40043 (n_18700, n21726);
  not g40044 (n_18701, n21727);
  and g40045 (n21728, n_18700, n_18701);
  not g40046 (n_18702, n21728);
  and g40047 (n21729, n_1590, n_18702);
  and g40048 (n21730, \a[23] , n21728);
  not g40049 (n_18703, n21729);
  not g40050 (n_18704, n21730);
  and g40051 (n21731, n_18703, n_18704);
  and g40052 (n21732, n_18489, n21731);
  not g40053 (n_18705, n21731);
  and g40054 (n21733, n21489, n_18705);
  not g40055 (n_18706, n21732);
  not g40056 (n_18707, n21733);
  and g40057 (n21734, n_18706, n_18707);
  and g40058 (n21735, \b[27] , n12668);
  and g40059 (n21736, \b[25] , n13047);
  and g40060 (n21737, \b[26] , n12663);
  and g40066 (n21740, n2990, n12671);
  not g40069 (n_18712, n21741);
  and g40070 (n21742, \a[62] , n_18712);
  not g40071 (n_18713, n21742);
  and g40072 (n21743, \a[62] , n_18713);
  and g40073 (n21744, n_18712, n_18713);
  not g40074 (n_18714, n21743);
  not g40075 (n_18715, n21744);
  and g40076 (n21745, n_18714, n_18715);
  not g40077 (n_18716, n21745);
  and g40078 (n21746, n21734, n_18716);
  not g40079 (n_18717, n21746);
  and g40080 (n21747, n21734, n_18717);
  and g40081 (n21748, n_18716, n_18717);
  not g40082 (n_18718, n21747);
  not g40083 (n_18719, n21748);
  and g40084 (n21749, n_18718, n_18719);
  not g40085 (n_18720, n21725);
  and g40086 (n21750, n_18720, n21749);
  not g40087 (n_18721, n21749);
  and g40088 (n21751, n21725, n_18721);
  not g40089 (n_18722, n21750);
  not g40090 (n_18723, n21751);
  and g40091 (n21752, n_18722, n_18723);
  and g40092 (n21753, \b[30] , n11531);
  and g40093 (n21754, \b[28] , n11896);
  and g40094 (n21755, \b[29] , n11526);
  and g40100 (n21758, n3577, n11534);
  not g40103 (n_18728, n21759);
  and g40104 (n21760, \a[59] , n_18728);
  not g40105 (n_18729, n21760);
  and g40106 (n21761, \a[59] , n_18729);
  and g40107 (n21762, n_18728, n_18729);
  not g40108 (n_18730, n21761);
  not g40109 (n_18731, n21762);
  and g40110 (n21763, n_18730, n_18731);
  not g40111 (n_18732, n21752);
  not g40112 (n_18733, n21763);
  and g40113 (n21764, n_18732, n_18733);
  and g40114 (n21765, n21752, n21763);
  not g40115 (n_18734, n21764);
  not g40116 (n_18735, n21765);
  and g40117 (n21766, n_18734, n_18735);
  not g40118 (n_18736, n21766);
  and g40119 (n21767, n21724, n_18736);
  not g40120 (n_18737, n21724);
  and g40121 (n21768, n_18737, n21766);
  not g40122 (n_18738, n21767);
  not g40123 (n_18739, n21768);
  and g40124 (n21769, n_18738, n_18739);
  and g40125 (n21770, \b[33] , n10426);
  and g40126 (n21771, \b[31] , n10796);
  and g40127 (n21772, \b[32] , n10421);
  and g40133 (n21775, n4223, n10429);
  not g40136 (n_18744, n21776);
  and g40137 (n21777, \a[56] , n_18744);
  not g40138 (n_18745, n21777);
  and g40139 (n21778, \a[56] , n_18745);
  and g40140 (n21779, n_18744, n_18745);
  not g40141 (n_18746, n21778);
  not g40142 (n_18747, n21779);
  and g40143 (n21780, n_18746, n_18747);
  and g40144 (n21781, n_18524, n_18536);
  not g40145 (n_18748, n21780);
  not g40146 (n_18749, n21781);
  and g40147 (n21782, n_18748, n_18749);
  and g40148 (n21783, n21780, n21781);
  not g40149 (n_18750, n21782);
  not g40150 (n_18751, n21783);
  and g40151 (n21784, n_18750, n_18751);
  and g40152 (n21785, n21769, n21784);
  not g40153 (n_18752, n21769);
  not g40154 (n_18753, n21784);
  and g40155 (n21786, n_18752, n_18753);
  not g40156 (n_18754, n21785);
  not g40157 (n_18755, n21786);
  and g40158 (n21787, n_18754, n_18755);
  not g40159 (n_18756, n21723);
  and g40160 (n21788, n_18756, n21787);
  not g40161 (n_18757, n21788);
  and g40162 (n21789, n21787, n_18757);
  and g40163 (n21790, n_18756, n_18757);
  not g40164 (n_18758, n21789);
  not g40165 (n_18759, n21790);
  and g40166 (n21791, n_18758, n_18759);
  and g40167 (n21792, n_18539, n_18543);
  and g40168 (n21793, n21791, n21792);
  not g40169 (n_18760, n21791);
  not g40170 (n_18761, n21792);
  and g40171 (n21794, n_18760, n_18761);
  not g40172 (n_18762, n21793);
  not g40173 (n_18763, n21794);
  and g40174 (n21795, n_18762, n_18763);
  and g40175 (n21796, \b[39] , n8362);
  and g40176 (n21797, \b[37] , n8715);
  and g40177 (n21798, \b[38] , n8357);
  and g40183 (n21801, n5451, n8365);
  not g40186 (n_18768, n21802);
  and g40187 (n21803, \a[50] , n_18768);
  not g40188 (n_18769, n21803);
  and g40189 (n21804, \a[50] , n_18769);
  and g40190 (n21805, n_18768, n_18769);
  not g40191 (n_18770, n21804);
  not g40192 (n_18771, n21805);
  and g40193 (n21806, n_18770, n_18771);
  not g40194 (n_18772, n21806);
  and g40195 (n21807, n21795, n_18772);
  not g40196 (n_18773, n21807);
  and g40197 (n21808, n21795, n_18773);
  and g40198 (n21809, n_18772, n_18773);
  not g40199 (n_18774, n21808);
  not g40200 (n_18775, n21809);
  and g40201 (n21810, n_18774, n_18775);
  and g40202 (n21811, n_18547, n_18558);
  and g40203 (n21812, n21810, n21811);
  not g40204 (n_18776, n21810);
  not g40205 (n_18777, n21811);
  and g40206 (n21813, n_18776, n_18777);
  not g40207 (n_18778, n21812);
  not g40208 (n_18779, n21813);
  and g40209 (n21814, n_18778, n_18779);
  and g40210 (n21815, \b[42] , n7446);
  and g40211 (n21816, \b[40] , n7787);
  and g40212 (n21817, \b[41] , n7441);
  and g40218 (n21820, n6489, n7449);
  not g40221 (n_18784, n21821);
  and g40222 (n21822, \a[47] , n_18784);
  not g40223 (n_18785, n21822);
  and g40224 (n21823, \a[47] , n_18785);
  and g40225 (n21824, n_18784, n_18785);
  not g40226 (n_18786, n21823);
  not g40227 (n_18787, n21824);
  and g40228 (n21825, n_18786, n_18787);
  not g40229 (n_18788, n21825);
  and g40230 (n21826, n21814, n_18788);
  not g40231 (n_18789, n21826);
  and g40232 (n21827, n21814, n_18789);
  and g40233 (n21828, n_18788, n_18789);
  not g40234 (n_18790, n21827);
  not g40235 (n_18791, n21828);
  and g40236 (n21829, n_18790, n_18791);
  not g40237 (n_18792, n21712);
  and g40238 (n21830, n_18792, n21829);
  not g40239 (n_18793, n21829);
  and g40240 (n21831, n21712, n_18793);
  not g40241 (n_18794, n21830);
  not g40242 (n_18795, n21831);
  and g40243 (n21832, n_18794, n_18795);
  and g40244 (n21833, \b[45] , n6595);
  and g40245 (n21834, \b[43] , n6902);
  and g40246 (n21835, \b[44] , n6590);
  and g40252 (n21838, n6598, n7361);
  not g40255 (n_18800, n21839);
  and g40256 (n21840, \a[44] , n_18800);
  not g40257 (n_18801, n21840);
  and g40258 (n21841, \a[44] , n_18801);
  and g40259 (n21842, n_18800, n_18801);
  not g40260 (n_18802, n21841);
  not g40261 (n_18803, n21842);
  and g40262 (n21843, n_18802, n_18803);
  not g40263 (n_18804, n21832);
  not g40264 (n_18805, n21843);
  and g40265 (n21844, n_18804, n_18805);
  and g40266 (n21845, n21832, n21843);
  not g40267 (n_18806, n21844);
  not g40268 (n_18807, n21845);
  and g40269 (n21846, n_18806, n_18807);
  not g40270 (n_18808, n21846);
  and g40271 (n21847, n21710, n_18808);
  not g40272 (n_18809, n21710);
  and g40273 (n21848, n_18809, n21846);
  not g40274 (n_18810, n21847);
  not g40275 (n_18811, n21848);
  and g40276 (n21849, n_18810, n_18811);
  and g40277 (n21850, \b[48] , n5777);
  and g40278 (n21851, \b[46] , n6059);
  and g40279 (n21852, \b[47] , n5772);
  and g40285 (n21855, n5780, n8009);
  not g40288 (n_18816, n21856);
  and g40289 (n21857, \a[41] , n_18816);
  not g40290 (n_18817, n21857);
  and g40291 (n21858, \a[41] , n_18817);
  and g40292 (n21859, n_18816, n_18817);
  not g40293 (n_18818, n21858);
  not g40294 (n_18819, n21859);
  and g40295 (n21860, n_18818, n_18819);
  not g40296 (n_18820, n21860);
  and g40297 (n21861, n21849, n_18820);
  not g40298 (n_18821, n21861);
  and g40299 (n21862, n21849, n_18821);
  and g40300 (n21863, n_18820, n_18821);
  not g40301 (n_18822, n21862);
  not g40302 (n_18823, n21863);
  and g40303 (n21864, n_18822, n_18823);
  and g40304 (n21865, n_18588, n_18599);
  and g40305 (n21866, n21864, n21865);
  not g40306 (n_18824, n21864);
  not g40307 (n_18825, n21865);
  and g40308 (n21867, n_18824, n_18825);
  not g40309 (n_18826, n21866);
  not g40310 (n_18827, n21867);
  and g40311 (n21868, n_18826, n_18827);
  and g40312 (n21869, \b[51] , n5035);
  and g40313 (n21870, \b[49] , n5277);
  and g40314 (n21871, \b[50] , n5030);
  and g40320 (n21874, n5038, n8976);
  not g40323 (n_18832, n21875);
  and g40324 (n21876, \a[38] , n_18832);
  not g40325 (n_18833, n21876);
  and g40326 (n21877, \a[38] , n_18833);
  and g40327 (n21878, n_18832, n_18833);
  not g40328 (n_18834, n21877);
  not g40329 (n_18835, n21878);
  and g40330 (n21879, n_18834, n_18835);
  not g40331 (n_18836, n21879);
  and g40332 (n21880, n21868, n_18836);
  not g40333 (n_18837, n21868);
  and g40334 (n21881, n_18837, n21879);
  not g40335 (n_18838, n21709);
  not g40336 (n_18839, n21881);
  and g40337 (n21882, n_18838, n_18839);
  not g40338 (n_18840, n21880);
  and g40339 (n21883, n_18840, n21882);
  not g40340 (n_18841, n21883);
  and g40341 (n21884, n_18838, n_18841);
  and g40342 (n21885, n_18840, n_18841);
  and g40343 (n21886, n_18839, n21885);
  not g40344 (n_18842, n21884);
  not g40345 (n_18843, n21886);
  and g40346 (n21887, n_18842, n_18843);
  and g40347 (n21888, \b[54] , n4287);
  and g40348 (n21889, \b[52] , n4532);
  and g40349 (n21890, \b[53] , n4282);
  and g40355 (n21893, n4290, n9998);
  not g40358 (n_18848, n21894);
  and g40359 (n21895, \a[35] , n_18848);
  not g40360 (n_18849, n21895);
  and g40361 (n21896, \a[35] , n_18849);
  and g40362 (n21897, n_18848, n_18849);
  not g40363 (n_18850, n21896);
  not g40364 (n_18851, n21897);
  and g40365 (n21898, n_18850, n_18851);
  and g40366 (n21899, n21887, n21898);
  not g40367 (n_18852, n21887);
  not g40368 (n_18853, n21898);
  and g40369 (n21900, n_18852, n_18853);
  not g40370 (n_18854, n21899);
  not g40371 (n_18855, n21900);
  and g40372 (n21901, n_18854, n_18855);
  not g40373 (n_18856, n21708);
  and g40374 (n21902, n_18856, n21901);
  not g40375 (n_18857, n21901);
  and g40376 (n21903, n21708, n_18857);
  not g40377 (n_18858, n21902);
  not g40378 (n_18859, n21903);
  and g40379 (n21904, n_18858, n_18859);
  and g40380 (n21905, n21707, n21904);
  not g40381 (n_18860, n21707);
  not g40382 (n_18861, n21904);
  and g40383 (n21906, n_18860, n_18861);
  not g40384 (n_18862, n21692);
  not g40385 (n_18863, n21906);
  and g40386 (n21907, n_18862, n_18863);
  not g40387 (n_18864, n21905);
  and g40388 (n21908, n_18864, n21907);
  not g40389 (n_18865, n21908);
  and g40390 (n21909, n_18862, n_18865);
  and g40391 (n21910, n_18863, n_18865);
  and g40392 (n21911, n_18864, n21910);
  not g40393 (n_18866, n21909);
  not g40394 (n_18867, n21911);
  and g40395 (n21912, n_18866, n_18867);
  not g40396 (n_18868, n21676);
  and g40397 (n21913, n_18868, n21912);
  not g40398 (n_18869, n21912);
  and g40399 (n21914, n21676, n_18869);
  not g40400 (n_18870, n21913);
  not g40401 (n_18871, n21914);
  and g40402 (n21915, n_18870, n_18871);
  not g40403 (n_18872, n21660);
  not g40404 (n_18873, n21915);
  and g40405 (n21916, n_18872, n_18873);
  not g40406 (n_18874, n21916);
  and g40407 (n21917, n_18872, n_18874);
  and g40408 (n21918, n_18873, n_18874);
  not g40409 (n_18875, n21917);
  not g40410 (n_18876, n21918);
  and g40411 (n21919, n_18875, n_18876);
  not g40412 (n_18877, n21658);
  not g40413 (n_18878, n21919);
  and g40414 (n21920, n_18877, n_18878);
  and g40415 (n21921, n21658, n_18876);
  and g40416 (n21922, n_18875, n21921);
  not g40417 (n_18879, n21920);
  not g40418 (n_18880, n21922);
  and g40419 (\f[87] , n_18879, n_18880);
  and g40420 (n21924, n_18874, n_18879);
  and g40421 (n21925, n_18868, n_18869);
  not g40422 (n_18881, n21925);
  and g40423 (n21926, n_18663, n_18881);
  and g40424 (n21927, \b[61] , n3050);
  and g40425 (n21928, \b[59] , n3243);
  and g40426 (n21929, \b[60] , n3045);
  and g40432 (n21932, n3053, n12969);
  not g40435 (n_18886, n21933);
  and g40436 (n21934, \a[29] , n_18886);
  not g40437 (n_18887, n21934);
  and g40438 (n21935, \a[29] , n_18887);
  and g40439 (n21936, n_18886, n_18887);
  not g40440 (n_18888, n21935);
  not g40441 (n_18889, n21936);
  and g40442 (n21937, n_18888, n_18889);
  and g40443 (n21938, n_18690, n_18864);
  not g40444 (n_18890, n21937);
  not g40445 (n_18891, n21938);
  and g40446 (n21939, n_18890, n_18891);
  not g40447 (n_18892, n21939);
  and g40448 (n21940, n_18890, n_18892);
  and g40449 (n21941, n_18891, n_18892);
  not g40450 (n_18893, n21940);
  not g40451 (n_18894, n21941);
  and g40452 (n21942, n_18893, n_18894);
  and g40453 (n21943, n_18855, n_18858);
  and g40454 (n21944, \b[58] , n3638);
  and g40455 (n21945, \b[56] , n3843);
  and g40456 (n21946, \b[57] , n3633);
  not g40457 (n_18895, n21945);
  not g40458 (n_18896, n21946);
  and g40459 (n21947, n_18895, n_18896);
  not g40460 (n_18897, n21944);
  and g40461 (n21948, n_18897, n21947);
  and g40462 (n21949, n_12780, n21948);
  and g40463 (n21950, n_13160, n21948);
  not g40464 (n_18898, n21949);
  not g40465 (n_18899, n21950);
  and g40466 (n21951, n_18898, n_18899);
  not g40467 (n_18900, n21951);
  and g40468 (n21952, \a[32] , n_18900);
  and g40469 (n21953, n_2992, n21951);
  not g40470 (n_18901, n21952);
  not g40471 (n_18902, n21953);
  and g40472 (n21954, n_18901, n_18902);
  not g40473 (n_18903, n21943);
  not g40474 (n_18904, n21954);
  and g40475 (n21955, n_18903, n_18904);
  and g40476 (n21956, n21943, n21954);
  not g40477 (n_18905, n21955);
  not g40478 (n_18906, n21956);
  and g40479 (n21957, n_18905, n_18906);
  and g40480 (n21958, \b[43] , n7446);
  and g40481 (n21959, \b[41] , n7787);
  and g40482 (n21960, \b[42] , n7441);
  and g40488 (n21963, n6515, n7449);
  not g40491 (n_18911, n21964);
  and g40492 (n21965, \a[47] , n_18911);
  not g40493 (n_18912, n21965);
  and g40494 (n21966, \a[47] , n_18912);
  and g40495 (n21967, n_18911, n_18912);
  not g40496 (n_18913, n21966);
  not g40497 (n_18914, n21967);
  and g40498 (n21968, n_18913, n_18914);
  and g40499 (n21969, n_18773, n_18779);
  and g40500 (n21970, \b[40] , n8362);
  and g40501 (n21971, \b[38] , n8715);
  and g40502 (n21972, \b[39] , n8357);
  and g40508 (n21975, n5955, n8365);
  not g40511 (n_18919, n21976);
  and g40512 (n21977, \a[50] , n_18919);
  not g40513 (n_18920, n21977);
  and g40514 (n21978, \a[50] , n_18920);
  and g40515 (n21979, n_18919, n_18920);
  not g40516 (n_18921, n21978);
  not g40517 (n_18922, n21979);
  and g40518 (n21980, n_18921, n_18922);
  and g40519 (n21981, n_18757, n_18763);
  and g40520 (n21982, n_18720, n_18721);
  not g40521 (n_18923, n21982);
  and g40522 (n21983, n_18717, n_18923);
  and g40523 (n21984, \b[24] , n13903);
  and g40524 (n21985, \b[25] , n_11555);
  not g40525 (n_18924, n21984);
  not g40526 (n_18925, n21985);
  and g40527 (n21986, n_18924, n_18925);
  and g40528 (n21987, n_18703, n_18706);
  not g40529 (n_18926, n21986);
  and g40530 (n21988, n_18926, n21987);
  not g40531 (n_18927, n21987);
  and g40532 (n21989, n21986, n_18927);
  not g40533 (n_18928, n21988);
  not g40534 (n_18929, n21989);
  and g40535 (n21990, n_18928, n_18929);
  and g40536 (n21991, \b[28] , n12668);
  and g40537 (n21992, \b[26] , n13047);
  and g40538 (n21993, \b[27] , n12663);
  not g40539 (n_18930, n21992);
  not g40540 (n_18931, n21993);
  and g40541 (n21994, n_18930, n_18931);
  not g40542 (n_18932, n21991);
  and g40543 (n21995, n_18932, n21994);
  and g40544 (n21996, n_12644, n21995);
  not g40545 (n_18933, n3189);
  and g40546 (n21997, n_18933, n21995);
  not g40547 (n_18934, n21996);
  not g40548 (n_18935, n21997);
  and g40549 (n21998, n_18934, n_18935);
  not g40550 (n_18936, n21998);
  and g40551 (n21999, \a[62] , n_18936);
  and g40552 (n22000, n_10843, n21998);
  not g40553 (n_18937, n21999);
  not g40554 (n_18938, n22000);
  and g40555 (n22001, n_18937, n_18938);
  not g40556 (n_18939, n22001);
  and g40557 (n22002, n21990, n_18939);
  not g40558 (n_18940, n21990);
  and g40559 (n22003, n_18940, n22001);
  not g40560 (n_18941, n22002);
  not g40561 (n_18942, n22003);
  and g40562 (n22004, n_18941, n_18942);
  not g40563 (n_18943, n21983);
  and g40564 (n22005, n_18943, n22004);
  not g40565 (n_18944, n22004);
  and g40566 (n22006, n21983, n_18944);
  not g40567 (n_18945, n22005);
  not g40568 (n_18946, n22006);
  and g40569 (n22007, n_18945, n_18946);
  and g40570 (n22008, \b[31] , n11531);
  and g40571 (n22009, \b[29] , n11896);
  and g40572 (n22010, \b[30] , n11526);
  and g40578 (n22013, n3796, n11534);
  not g40581 (n_18951, n22014);
  and g40582 (n22015, \a[59] , n_18951);
  not g40583 (n_18952, n22015);
  and g40584 (n22016, \a[59] , n_18952);
  and g40585 (n22017, n_18951, n_18952);
  not g40586 (n_18953, n22016);
  not g40587 (n_18954, n22017);
  and g40588 (n22018, n_18953, n_18954);
  not g40589 (n_18955, n22018);
  and g40590 (n22019, n22007, n_18955);
  not g40591 (n_18956, n22019);
  and g40592 (n22020, n22007, n_18956);
  and g40593 (n22021, n_18955, n_18956);
  not g40594 (n_18957, n22020);
  not g40595 (n_18958, n22021);
  and g40596 (n22022, n_18957, n_18958);
  and g40597 (n22023, n_18734, n_18739);
  and g40598 (n22024, n22022, n22023);
  not g40599 (n_18959, n22022);
  not g40600 (n_18960, n22023);
  and g40601 (n22025, n_18959, n_18960);
  not g40602 (n_18961, n22024);
  not g40603 (n_18962, n22025);
  and g40604 (n22026, n_18961, n_18962);
  and g40605 (n22027, \b[34] , n10426);
  and g40606 (n22028, \b[32] , n10796);
  and g40607 (n22029, \b[33] , n10421);
  and g40613 (n22032, n4466, n10429);
  not g40616 (n_18967, n22033);
  and g40617 (n22034, \a[56] , n_18967);
  not g40618 (n_18968, n22034);
  and g40619 (n22035, \a[56] , n_18968);
  and g40620 (n22036, n_18967, n_18968);
  not g40621 (n_18969, n22035);
  not g40622 (n_18970, n22036);
  and g40623 (n22037, n_18969, n_18970);
  not g40624 (n_18971, n22037);
  and g40625 (n22038, n22026, n_18971);
  not g40626 (n_18972, n22038);
  and g40627 (n22039, n22026, n_18972);
  and g40628 (n22040, n_18971, n_18972);
  not g40629 (n_18973, n22039);
  not g40630 (n_18974, n22040);
  and g40631 (n22041, n_18973, n_18974);
  and g40632 (n22042, n_18750, n_18754);
  and g40633 (n22043, n22041, n22042);
  not g40634 (n_18975, n22041);
  not g40635 (n_18976, n22042);
  and g40636 (n22044, n_18975, n_18976);
  not g40637 (n_18977, n22043);
  not g40638 (n_18978, n22044);
  and g40639 (n22045, n_18977, n_18978);
  and g40640 (n22046, \b[37] , n9339);
  and g40641 (n22047, \b[35] , n9732);
  and g40642 (n22048, \b[36] , n9334);
  and g40648 (n22051, n5181, n9342);
  not g40651 (n_18983, n22052);
  and g40652 (n22053, \a[53] , n_18983);
  not g40653 (n_18984, n22053);
  and g40654 (n22054, \a[53] , n_18984);
  and g40655 (n22055, n_18983, n_18984);
  not g40656 (n_18985, n22054);
  not g40657 (n_18986, n22055);
  and g40658 (n22056, n_18985, n_18986);
  not g40659 (n_18987, n22045);
  and g40660 (n22057, n_18987, n22056);
  not g40661 (n_18988, n22056);
  and g40662 (n22058, n22045, n_18988);
  not g40663 (n_18989, n22057);
  not g40664 (n_18990, n22058);
  and g40665 (n22059, n_18989, n_18990);
  not g40666 (n_18991, n21981);
  and g40667 (n22060, n_18991, n22059);
  not g40668 (n_18992, n22060);
  and g40669 (n22061, n_18991, n_18992);
  and g40670 (n22062, n22059, n_18992);
  not g40671 (n_18993, n22061);
  not g40672 (n_18994, n22062);
  and g40673 (n22063, n_18993, n_18994);
  not g40674 (n_18995, n21980);
  not g40675 (n_18996, n22063);
  and g40676 (n22064, n_18995, n_18996);
  and g40677 (n22065, n21980, n_18994);
  and g40678 (n22066, n_18993, n22065);
  not g40679 (n_18997, n22064);
  not g40680 (n_18998, n22066);
  and g40681 (n22067, n_18997, n_18998);
  not g40682 (n_18999, n21969);
  and g40683 (n22068, n_18999, n22067);
  not g40684 (n_19000, n22067);
  and g40685 (n22069, n21969, n_19000);
  not g40686 (n_19001, n22068);
  not g40687 (n_19002, n22069);
  and g40688 (n22070, n_19001, n_19002);
  not g40689 (n_19003, n21968);
  and g40690 (n22071, n_19003, n22070);
  not g40691 (n_19004, n22071);
  and g40692 (n22072, n22070, n_19004);
  and g40693 (n22073, n_19003, n_19004);
  not g40694 (n_19005, n22072);
  not g40695 (n_19006, n22073);
  and g40696 (n22074, n_19005, n_19006);
  and g40697 (n22075, n_18792, n_18793);
  not g40698 (n_19007, n22075);
  and g40699 (n22076, n_18789, n_19007);
  and g40700 (n22077, n22074, n22076);
  not g40701 (n_19008, n22074);
  not g40702 (n_19009, n22076);
  and g40703 (n22078, n_19008, n_19009);
  not g40704 (n_19010, n22077);
  not g40705 (n_19011, n22078);
  and g40706 (n22079, n_19010, n_19011);
  and g40707 (n22080, \b[46] , n6595);
  and g40708 (n22081, \b[44] , n6902);
  and g40709 (n22082, \b[45] , n6590);
  and g40715 (n22085, n6598, n7677);
  not g40718 (n_19016, n22086);
  and g40719 (n22087, \a[44] , n_19016);
  not g40720 (n_19017, n22087);
  and g40721 (n22088, \a[44] , n_19017);
  and g40722 (n22089, n_19016, n_19017);
  not g40723 (n_19018, n22088);
  not g40724 (n_19019, n22089);
  and g40725 (n22090, n_19018, n_19019);
  not g40726 (n_19020, n22090);
  and g40727 (n22091, n22079, n_19020);
  not g40728 (n_19021, n22091);
  and g40729 (n22092, n22079, n_19021);
  and g40730 (n22093, n_19020, n_19021);
  not g40731 (n_19022, n22092);
  not g40732 (n_19023, n22093);
  and g40733 (n22094, n_19022, n_19023);
  and g40734 (n22095, n_18806, n_18811);
  and g40735 (n22096, n22094, n22095);
  not g40736 (n_19024, n22094);
  not g40737 (n_19025, n22095);
  and g40738 (n22097, n_19024, n_19025);
  not g40739 (n_19026, n22096);
  not g40740 (n_19027, n22097);
  and g40741 (n22098, n_19026, n_19027);
  and g40742 (n22099, \b[49] , n5777);
  and g40743 (n22100, \b[47] , n6059);
  and g40744 (n22101, \b[48] , n5772);
  and g40750 (n22104, n5780, n8625);
  not g40753 (n_19032, n22105);
  and g40754 (n22106, \a[41] , n_19032);
  not g40755 (n_19033, n22106);
  and g40756 (n22107, \a[41] , n_19033);
  and g40757 (n22108, n_19032, n_19033);
  not g40758 (n_19034, n22107);
  not g40759 (n_19035, n22108);
  and g40760 (n22109, n_19034, n_19035);
  not g40761 (n_19036, n22109);
  and g40762 (n22110, n22098, n_19036);
  not g40763 (n_19037, n22110);
  and g40764 (n22111, n22098, n_19037);
  and g40765 (n22112, n_19036, n_19037);
  not g40766 (n_19038, n22111);
  not g40767 (n_19039, n22112);
  and g40768 (n22113, n_19038, n_19039);
  and g40769 (n22114, n_18821, n_18827);
  and g40770 (n22115, n22113, n22114);
  not g40771 (n_19040, n22113);
  not g40772 (n_19041, n22114);
  and g40773 (n22116, n_19040, n_19041);
  not g40774 (n_19042, n22115);
  not g40775 (n_19043, n22116);
  and g40776 (n22117, n_19042, n_19043);
  and g40777 (n22118, \b[52] , n5035);
  and g40778 (n22119, \b[50] , n5277);
  and g40779 (n22120, \b[51] , n5030);
  and g40785 (n22123, n5038, n9628);
  not g40788 (n_19048, n22124);
  and g40789 (n22125, \a[38] , n_19048);
  not g40790 (n_19049, n22125);
  and g40791 (n22126, \a[38] , n_19049);
  and g40792 (n22127, n_19048, n_19049);
  not g40793 (n_19050, n22126);
  not g40794 (n_19051, n22127);
  and g40795 (n22128, n_19050, n_19051);
  not g40796 (n_19052, n22128);
  and g40797 (n22129, n22117, n_19052);
  not g40798 (n_19053, n22129);
  and g40799 (n22130, n22117, n_19053);
  and g40800 (n22131, n_19052, n_19053);
  not g40801 (n_19054, n22130);
  not g40802 (n_19055, n22131);
  and g40803 (n22132, n_19054, n_19055);
  not g40804 (n_19056, n21885);
  and g40805 (n22133, n_19056, n22132);
  not g40806 (n_19057, n22132);
  and g40807 (n22134, n21885, n_19057);
  not g40808 (n_19058, n22133);
  not g40809 (n_19059, n22134);
  and g40810 (n22135, n_19058, n_19059);
  and g40811 (n22136, \b[55] , n4287);
  and g40812 (n22137, \b[53] , n4532);
  and g40813 (n22138, \b[54] , n4282);
  and g40819 (n22141, n4290, n10684);
  not g40822 (n_19064, n22142);
  and g40823 (n22143, \a[35] , n_19064);
  not g40824 (n_19065, n22143);
  and g40825 (n22144, \a[35] , n_19065);
  and g40826 (n22145, n_19064, n_19065);
  not g40827 (n_19066, n22144);
  not g40828 (n_19067, n22145);
  and g40829 (n22146, n_19066, n_19067);
  not g40830 (n_19068, n22135);
  not g40831 (n_19069, n22146);
  and g40832 (n22147, n_19068, n_19069);
  and g40833 (n22148, n22135, n22146);
  not g40834 (n_19070, n22147);
  not g40835 (n_19071, n22148);
  and g40836 (n22149, n_19070, n_19071);
  and g40837 (n22150, n21957, n22149);
  not g40838 (n_19072, n21957);
  not g40839 (n_19073, n22149);
  and g40840 (n22151, n_19072, n_19073);
  not g40841 (n_19074, n22150);
  not g40842 (n_19075, n22151);
  and g40843 (n22152, n_19074, n_19075);
  not g40844 (n_19076, n21942);
  and g40845 (n22153, n_19076, n22152);
  not g40846 (n_19077, n22153);
  and g40847 (n22154, n_19076, n_19077);
  and g40848 (n22155, n22152, n_19077);
  not g40849 (n_19078, n22154);
  not g40850 (n_19079, n22155);
  and g40851 (n22156, n_19078, n_19079);
  and g40852 (n22157, n_18675, n_18676);
  not g40853 (n_19080, n22157);
  and g40854 (n22158, n_18865, n_19080);
  and g40855 (n22159, \b[62] , n2685);
  and g40856 (n22160, \b[63] , n2534);
  not g40857 (n_19081, n22159);
  not g40858 (n_19082, n22160);
  and g40859 (n22161, n_19081, n_19082);
  and g40860 (n22162, n_13498, n22161);
  and g40861 (n22163, n13800, n22161);
  not g40862 (n_19083, n22162);
  not g40863 (n_19084, n22163);
  and g40864 (n22164, n_19083, n_19084);
  not g40865 (n_19085, n22164);
  and g40866 (n22165, \a[26] , n_19085);
  and g40867 (n22166, n_2025, n22164);
  not g40868 (n_19086, n22165);
  not g40869 (n_19087, n22166);
  and g40870 (n22167, n_19086, n_19087);
  not g40871 (n_19088, n22158);
  not g40872 (n_19089, n22167);
  and g40873 (n22168, n_19088, n_19089);
  not g40874 (n_19090, n22168);
  and g40875 (n22169, n_19088, n_19090);
  and g40876 (n22170, n_19089, n_19090);
  not g40877 (n_19091, n22169);
  not g40878 (n_19092, n22170);
  and g40879 (n22171, n_19091, n_19092);
  not g40880 (n_19093, n22156);
  not g40881 (n_19094, n22171);
  and g40882 (n22172, n_19093, n_19094);
  and g40883 (n22173, n22156, n_19092);
  and g40884 (n22174, n_19091, n22173);
  not g40885 (n_19095, n22172);
  not g40886 (n_19096, n22174);
  and g40887 (n22175, n_19095, n_19096);
  not g40888 (n_19097, n21926);
  and g40889 (n22176, n_19097, n22175);
  not g40890 (n_19098, n22176);
  and g40891 (n22177, n_19097, n_19098);
  and g40892 (n22178, n22175, n_19098);
  not g40893 (n_19099, n22177);
  not g40894 (n_19100, n22178);
  and g40895 (n22179, n_19099, n_19100);
  not g40896 (n_19101, n21924);
  not g40897 (n_19102, n22179);
  and g40898 (n22180, n_19101, n_19102);
  and g40899 (n22181, n21924, n_19100);
  and g40900 (n22182, n_19099, n22181);
  not g40901 (n_19103, n22180);
  not g40902 (n_19104, n22182);
  and g40903 (\f[88] , n_19103, n_19104);
  and g40904 (n22184, n_19098, n_19103);
  and g40905 (n22185, n_19090, n_19095);
  and g40906 (n22186, n_18892, n_19077);
  and g40907 (n22187, \b[63] , n2685);
  and g40908 (n22188, n2542, n13797);
  not g40909 (n_19105, n22187);
  not g40910 (n_19106, n22188);
  and g40911 (n22189, n_19105, n_19106);
  not g40912 (n_19107, n22189);
  and g40913 (n22190, \a[26] , n_19107);
  not g40914 (n_19108, n22190);
  and g40915 (n22191, \a[26] , n_19108);
  and g40916 (n22192, n_19107, n_19108);
  not g40917 (n_19109, n22191);
  not g40918 (n_19110, n22192);
  and g40919 (n22193, n_19109, n_19110);
  not g40920 (n_19111, n22186);
  not g40921 (n_19112, n22193);
  and g40922 (n22194, n_19111, n_19112);
  not g40923 (n_19113, n22194);
  and g40924 (n22195, n_19111, n_19113);
  and g40925 (n22196, n_19112, n_19113);
  not g40926 (n_19114, n22195);
  not g40927 (n_19115, n22196);
  and g40928 (n22197, n_19114, n_19115);
  and g40929 (n22198, \b[62] , n3050);
  and g40930 (n22199, \b[60] , n3243);
  and g40931 (n22200, \b[61] , n3045);
  and g40937 (n22203, n3053, n13370);
  not g40940 (n_19120, n22204);
  and g40941 (n22205, \a[29] , n_19120);
  not g40942 (n_19121, n22205);
  and g40943 (n22206, \a[29] , n_19121);
  and g40944 (n22207, n_19120, n_19121);
  not g40945 (n_19122, n22206);
  not g40946 (n_19123, n22207);
  and g40947 (n22208, n_19122, n_19123);
  and g40948 (n22209, n_18905, n_19074);
  and g40949 (n22210, n22208, n22209);
  not g40950 (n_19124, n22208);
  not g40951 (n_19125, n22209);
  and g40952 (n22211, n_19124, n_19125);
  not g40953 (n_19126, n22210);
  not g40954 (n_19127, n22211);
  and g40955 (n22212, n_19126, n_19127);
  and g40956 (n22213, \b[59] , n3638);
  and g40957 (n22214, \b[57] , n3843);
  and g40958 (n22215, \b[58] , n3633);
  and g40964 (n22218, n3641, n12179);
  not g40967 (n_19132, n22219);
  and g40968 (n22220, \a[32] , n_19132);
  not g40969 (n_19133, n22220);
  and g40970 (n22221, \a[32] , n_19133);
  and g40971 (n22222, n_19132, n_19133);
  not g40972 (n_19134, n22221);
  not g40973 (n_19135, n22222);
  and g40974 (n22223, n_19134, n_19135);
  and g40975 (n22224, n_19056, n_19057);
  not g40976 (n_19136, n22224);
  and g40977 (n22225, n_19070, n_19136);
  and g40978 (n22226, n22223, n22225);
  not g40979 (n_19137, n22223);
  not g40980 (n_19138, n22225);
  and g40981 (n22227, n_19137, n_19138);
  not g40982 (n_19139, n22226);
  not g40983 (n_19140, n22227);
  and g40984 (n22228, n_19139, n_19140);
  and g40985 (n22229, \b[56] , n4287);
  and g40986 (n22230, \b[54] , n4532);
  and g40987 (n22231, \b[55] , n4282);
  and g40993 (n22234, n4290, n10708);
  not g40996 (n_19145, n22235);
  and g40997 (n22236, \a[35] , n_19145);
  not g40998 (n_19146, n22236);
  and g40999 (n22237, \a[35] , n_19146);
  and g41000 (n22238, n_19145, n_19146);
  not g41001 (n_19147, n22237);
  not g41002 (n_19148, n22238);
  and g41003 (n22239, n_19147, n_19148);
  and g41004 (n22240, n_19043, n_19053);
  and g41005 (n22241, \b[53] , n5035);
  and g41006 (n22242, \b[51] , n5277);
  and g41007 (n22243, \b[52] , n5030);
  and g41013 (n22246, n5038, n9972);
  not g41016 (n_19153, n22247);
  and g41017 (n22248, \a[38] , n_19153);
  not g41018 (n_19154, n22248);
  and g41019 (n22249, \a[38] , n_19154);
  and g41020 (n22250, n_19153, n_19154);
  not g41021 (n_19155, n22249);
  not g41022 (n_19156, n22250);
  and g41023 (n22251, n_19155, n_19156);
  and g41024 (n22252, n_19027, n_19037);
  and g41025 (n22253, n_19001, n_19004);
  and g41026 (n22254, \b[44] , n7446);
  and g41027 (n22255, \b[42] , n7787);
  and g41028 (n22256, \b[43] , n7441);
  and g41034 (n22259, n7072, n7449);
  not g41037 (n_19161, n22260);
  and g41038 (n22261, \a[47] , n_19161);
  not g41039 (n_19162, n22261);
  and g41040 (n22262, \a[47] , n_19162);
  and g41041 (n22263, n_19161, n_19162);
  not g41042 (n_19163, n22262);
  not g41043 (n_19164, n22263);
  and g41044 (n22264, n_19163, n_19164);
  and g41045 (n22265, n_18992, n_18997);
  and g41046 (n22266, n_18962, n_18972);
  and g41047 (n22267, \b[35] , n10426);
  and g41048 (n22268, \b[33] , n10796);
  and g41049 (n22269, \b[34] , n10421);
  and g41055 (n22272, n4696, n10429);
  not g41058 (n_19169, n22273);
  and g41059 (n22274, \a[56] , n_19169);
  not g41060 (n_19170, n22274);
  and g41061 (n22275, \a[56] , n_19170);
  and g41062 (n22276, n_19169, n_19170);
  not g41063 (n_19171, n22275);
  not g41064 (n_19172, n22276);
  and g41065 (n22277, n_19171, n_19172);
  and g41066 (n22278, n_18945, n_18956);
  and g41067 (n22279, \b[32] , n11531);
  and g41068 (n22280, \b[30] , n11896);
  and g41069 (n22281, \b[31] , n11526);
  and g41075 (n22284, n4013, n11534);
  not g41078 (n_19177, n22285);
  and g41079 (n22286, \a[59] , n_19177);
  not g41080 (n_19178, n22286);
  and g41081 (n22287, \a[59] , n_19178);
  and g41082 (n22288, n_19177, n_19178);
  not g41083 (n_19179, n22287);
  not g41084 (n_19180, n22288);
  and g41085 (n22289, n_19179, n_19180);
  and g41086 (n22290, n_18929, n_18941);
  and g41087 (n22291, \b[25] , n13903);
  and g41088 (n22292, \b[26] , n_11555);
  not g41089 (n_19181, n22291);
  not g41090 (n_19182, n22292);
  and g41091 (n22293, n_19181, n_19182);
  and g41092 (n22294, n_18926, n22293);
  not g41093 (n_19183, n22293);
  and g41094 (n22295, n21986, n_19183);
  not g41095 (n_19184, n22294);
  not g41096 (n_19185, n22295);
  and g41097 (n22296, n_19184, n_19185);
  and g41098 (n22297, \b[29] , n12668);
  and g41099 (n22298, \b[27] , n13047);
  and g41100 (n22299, \b[28] , n12663);
  not g41101 (n_19186, n22298);
  not g41102 (n_19187, n22299);
  and g41103 (n22300, n_19186, n_19187);
  not g41104 (n_19188, n22297);
  and g41105 (n22301, n_19188, n22300);
  and g41106 (n22302, n_12644, n22301);
  not g41107 (n_19189, n3383);
  and g41108 (n22303, n_19189, n22301);
  not g41109 (n_19190, n22302);
  not g41110 (n_19191, n22303);
  and g41111 (n22304, n_19190, n_19191);
  not g41112 (n_19192, n22304);
  and g41113 (n22305, \a[62] , n_19192);
  and g41114 (n22306, n_10843, n22304);
  not g41115 (n_19193, n22305);
  not g41116 (n_19194, n22306);
  and g41117 (n22307, n_19193, n_19194);
  not g41118 (n_19195, n22307);
  and g41119 (n22308, n22296, n_19195);
  not g41120 (n_19196, n22296);
  and g41121 (n22309, n_19196, n22307);
  not g41122 (n_19197, n22308);
  not g41123 (n_19198, n22309);
  and g41124 (n22310, n_19197, n_19198);
  not g41125 (n_19199, n22290);
  and g41126 (n22311, n_19199, n22310);
  not g41127 (n_19200, n22310);
  and g41128 (n22312, n22290, n_19200);
  not g41129 (n_19201, n22311);
  not g41130 (n_19202, n22312);
  and g41131 (n22313, n_19201, n_19202);
  not g41132 (n_19203, n22289);
  and g41133 (n22314, n_19203, n22313);
  not g41134 (n_19204, n22313);
  and g41135 (n22315, n22289, n_19204);
  not g41136 (n_19205, n22314);
  not g41137 (n_19206, n22315);
  and g41138 (n22316, n_19205, n_19206);
  not g41139 (n_19207, n22278);
  and g41140 (n22317, n_19207, n22316);
  not g41141 (n_19208, n22316);
  and g41142 (n22318, n22278, n_19208);
  not g41143 (n_19209, n22317);
  not g41144 (n_19210, n22318);
  and g41145 (n22319, n_19209, n_19210);
  not g41146 (n_19211, n22277);
  and g41147 (n22320, n_19211, n22319);
  not g41148 (n_19212, n22319);
  and g41149 (n22321, n22277, n_19212);
  not g41150 (n_19213, n22320);
  not g41151 (n_19214, n22321);
  and g41152 (n22322, n_19213, n_19214);
  not g41153 (n_19215, n22266);
  and g41154 (n22323, n_19215, n22322);
  not g41155 (n_19216, n22322);
  and g41156 (n22324, n22266, n_19216);
  not g41157 (n_19217, n22323);
  not g41158 (n_19218, n22324);
  and g41159 (n22325, n_19217, n_19218);
  and g41160 (n22326, \b[38] , n9339);
  and g41161 (n22327, \b[36] , n9732);
  and g41162 (n22328, \b[37] , n9334);
  and g41168 (n22331, n5205, n9342);
  not g41171 (n_19223, n22332);
  and g41172 (n22333, \a[53] , n_19223);
  not g41173 (n_19224, n22333);
  and g41174 (n22334, \a[53] , n_19224);
  and g41175 (n22335, n_19223, n_19224);
  not g41176 (n_19225, n22334);
  not g41177 (n_19226, n22335);
  and g41178 (n22336, n_19225, n_19226);
  not g41179 (n_19227, n22336);
  and g41180 (n22337, n22325, n_19227);
  not g41181 (n_19228, n22337);
  and g41182 (n22338, n22325, n_19228);
  and g41183 (n22339, n_19227, n_19228);
  not g41184 (n_19229, n22338);
  not g41185 (n_19230, n22339);
  and g41186 (n22340, n_19229, n_19230);
  and g41187 (n22341, n_18978, n_18990);
  not g41188 (n_19231, n22340);
  not g41189 (n_19232, n22341);
  and g41190 (n22342, n_19231, n_19232);
  not g41191 (n_19233, n22342);
  and g41192 (n22343, n_19231, n_19233);
  and g41193 (n22344, n_19232, n_19233);
  not g41194 (n_19234, n22343);
  not g41195 (n_19235, n22344);
  and g41196 (n22345, n_19234, n_19235);
  and g41197 (n22346, \b[41] , n8362);
  and g41198 (n22347, \b[39] , n8715);
  and g41199 (n22348, \b[40] , n8357);
  and g41205 (n22351, n6219, n8365);
  not g41208 (n_19240, n22352);
  and g41209 (n22353, \a[50] , n_19240);
  not g41210 (n_19241, n22353);
  and g41211 (n22354, \a[50] , n_19241);
  and g41212 (n22355, n_19240, n_19241);
  not g41213 (n_19242, n22354);
  not g41214 (n_19243, n22355);
  and g41215 (n22356, n_19242, n_19243);
  not g41216 (n_19244, n22345);
  and g41217 (n22357, n_19244, n22356);
  not g41218 (n_19245, n22356);
  and g41219 (n22358, n22345, n_19245);
  not g41220 (n_19246, n22357);
  not g41221 (n_19247, n22358);
  and g41222 (n22359, n_19246, n_19247);
  not g41223 (n_19248, n22265);
  not g41224 (n_19249, n22359);
  and g41225 (n22360, n_19248, n_19249);
  and g41226 (n22361, n22265, n22359);
  not g41227 (n_19250, n22360);
  not g41228 (n_19251, n22361);
  and g41229 (n22362, n_19250, n_19251);
  not g41230 (n_19252, n22264);
  and g41231 (n22363, n_19252, n22362);
  not g41232 (n_19253, n22362);
  and g41233 (n22364, n22264, n_19253);
  not g41234 (n_19254, n22363);
  not g41235 (n_19255, n22364);
  and g41236 (n22365, n_19254, n_19255);
  not g41237 (n_19256, n22253);
  and g41238 (n22366, n_19256, n22365);
  not g41239 (n_19257, n22365);
  and g41240 (n22367, n22253, n_19257);
  not g41241 (n_19258, n22366);
  not g41242 (n_19259, n22367);
  and g41243 (n22368, n_19258, n_19259);
  and g41244 (n22369, \b[47] , n6595);
  and g41245 (n22370, \b[45] , n6902);
  and g41246 (n22371, \b[46] , n6590);
  and g41252 (n22374, n6598, n7703);
  not g41255 (n_19264, n22375);
  and g41256 (n22376, \a[44] , n_19264);
  not g41257 (n_19265, n22376);
  and g41258 (n22377, \a[44] , n_19265);
  and g41259 (n22378, n_19264, n_19265);
  not g41260 (n_19266, n22377);
  not g41261 (n_19267, n22378);
  and g41262 (n22379, n_19266, n_19267);
  not g41263 (n_19268, n22379);
  and g41264 (n22380, n22368, n_19268);
  not g41265 (n_19269, n22380);
  and g41266 (n22381, n22368, n_19269);
  and g41267 (n22382, n_19268, n_19269);
  not g41268 (n_19270, n22381);
  not g41269 (n_19271, n22382);
  and g41270 (n22383, n_19270, n_19271);
  and g41271 (n22384, n_19011, n_19021);
  and g41272 (n22385, n22383, n22384);
  not g41273 (n_19272, n22383);
  not g41274 (n_19273, n22384);
  and g41275 (n22386, n_19272, n_19273);
  not g41276 (n_19274, n22385);
  not g41277 (n_19275, n22386);
  and g41278 (n22387, n_19274, n_19275);
  and g41279 (n22388, \b[50] , n5777);
  and g41280 (n22389, \b[48] , n6059);
  and g41281 (n22390, \b[49] , n5772);
  and g41287 (n22393, n5780, n8949);
  not g41290 (n_19280, n22394);
  and g41291 (n22395, \a[41] , n_19280);
  not g41292 (n_19281, n22395);
  and g41293 (n22396, \a[41] , n_19281);
  and g41294 (n22397, n_19280, n_19281);
  not g41295 (n_19282, n22396);
  not g41296 (n_19283, n22397);
  and g41297 (n22398, n_19282, n_19283);
  not g41298 (n_19284, n22387);
  and g41299 (n22399, n_19284, n22398);
  not g41300 (n_19285, n22398);
  and g41301 (n22400, n22387, n_19285);
  not g41302 (n_19286, n22399);
  not g41303 (n_19287, n22400);
  and g41304 (n22401, n_19286, n_19287);
  not g41305 (n_19288, n22252);
  and g41306 (n22402, n_19288, n22401);
  not g41307 (n_19289, n22402);
  and g41308 (n22403, n_19288, n_19289);
  and g41309 (n22404, n22401, n_19289);
  not g41310 (n_19290, n22403);
  not g41311 (n_19291, n22404);
  and g41312 (n22405, n_19290, n_19291);
  not g41313 (n_19292, n22251);
  not g41314 (n_19293, n22405);
  and g41315 (n22406, n_19292, n_19293);
  and g41316 (n22407, n22251, n_19291);
  and g41317 (n22408, n_19290, n22407);
  not g41318 (n_19294, n22406);
  not g41319 (n_19295, n22408);
  and g41320 (n22409, n_19294, n_19295);
  not g41321 (n_19296, n22240);
  and g41322 (n22410, n_19296, n22409);
  not g41323 (n_19297, n22409);
  and g41324 (n22411, n22240, n_19297);
  not g41325 (n_19298, n22410);
  not g41326 (n_19299, n22411);
  and g41327 (n22412, n_19298, n_19299);
  not g41328 (n_19300, n22239);
  and g41329 (n22413, n_19300, n22412);
  not g41330 (n_19301, n22413);
  and g41331 (n22414, n_19300, n_19301);
  and g41332 (n22415, n22412, n_19301);
  not g41333 (n_19302, n22414);
  not g41334 (n_19303, n22415);
  and g41335 (n22416, n_19302, n_19303);
  not g41336 (n_19304, n22416);
  and g41337 (n22417, n22228, n_19304);
  not g41338 (n_19305, n22417);
  and g41339 (n22418, n22228, n_19305);
  and g41340 (n22419, n_19304, n_19305);
  not g41341 (n_19306, n22418);
  not g41342 (n_19307, n22419);
  and g41343 (n22420, n_19306, n_19307);
  not g41344 (n_19308, n22212);
  and g41345 (n22421, n_19308, n22420);
  not g41346 (n_19309, n22420);
  and g41347 (n22422, n22212, n_19309);
  not g41348 (n_19310, n22421);
  not g41349 (n_19311, n22422);
  and g41350 (n22423, n_19310, n_19311);
  not g41351 (n_19312, n22197);
  and g41352 (n22424, n_19312, n22423);
  not g41353 (n_19313, n22423);
  and g41354 (n22425, n22197, n_19313);
  not g41355 (n_19314, n22424);
  not g41356 (n_19315, n22425);
  and g41357 (n22426, n_19314, n_19315);
  not g41358 (n_19316, n22185);
  and g41359 (n22427, n_19316, n22426);
  not g41360 (n_19317, n22426);
  and g41361 (n22428, n22185, n_19317);
  not g41362 (n_19318, n22427);
  not g41363 (n_19319, n22428);
  and g41364 (n22429, n_19318, n_19319);
  not g41365 (n_19320, n22184);
  and g41366 (n22430, n_19320, n22429);
  not g41367 (n_19321, n22429);
  and g41368 (n22431, n22184, n_19321);
  not g41369 (n_19322, n22430);
  not g41370 (n_19323, n22431);
  and g41371 (\f[89] , n_19322, n_19323);
  and g41372 (n22433, n_19113, n_19314);
  and g41373 (n22434, n_19127, n_19311);
  and g41374 (n22435, \b[63] , n3050);
  and g41375 (n22436, \b[61] , n3243);
  and g41376 (n22437, \b[62] , n3045);
  and g41382 (n22440, n3053, n13771);
  not g41385 (n_19328, n22441);
  and g41386 (n22442, \a[29] , n_19328);
  not g41387 (n_19329, n22442);
  and g41388 (n22443, \a[29] , n_19329);
  and g41389 (n22444, n_19328, n_19329);
  not g41390 (n_19330, n22443);
  not g41391 (n_19331, n22444);
  and g41392 (n22445, n_19330, n_19331);
  not g41393 (n_19332, n22434);
  not g41394 (n_19333, n22445);
  and g41395 (n22446, n_19332, n_19333);
  not g41396 (n_19334, n22446);
  and g41397 (n22447, n_19332, n_19334);
  and g41398 (n22448, n_19333, n_19334);
  not g41399 (n_19335, n22447);
  not g41400 (n_19336, n22448);
  and g41401 (n22449, n_19335, n_19336);
  and g41402 (n22450, \b[57] , n4287);
  and g41403 (n22451, \b[55] , n4532);
  and g41404 (n22452, \b[56] , n4282);
  and g41410 (n22455, n4290, n11410);
  not g41413 (n_19341, n22456);
  and g41414 (n22457, \a[35] , n_19341);
  not g41415 (n_19342, n22457);
  and g41416 (n22458, \a[35] , n_19342);
  and g41417 (n22459, n_19341, n_19342);
  not g41418 (n_19343, n22458);
  not g41419 (n_19344, n22459);
  and g41420 (n22460, n_19343, n_19344);
  and g41421 (n22461, n_19289, n_19294);
  and g41422 (n22462, n_19275, n_19287);
  and g41423 (n22463, n_19250, n_19254);
  and g41424 (n22464, n_19244, n_19245);
  not g41425 (n_19345, n22464);
  and g41426 (n22465, n_19233, n_19345);
  and g41427 (n22466, \b[33] , n11531);
  and g41428 (n22467, \b[31] , n11896);
  and g41429 (n22468, \b[32] , n11526);
  and g41435 (n22471, n4223, n11534);
  not g41438 (n_19350, n22472);
  and g41439 (n22473, \a[59] , n_19350);
  not g41440 (n_19351, n22473);
  and g41441 (n22474, \a[59] , n_19351);
  and g41442 (n22475, n_19350, n_19351);
  not g41443 (n_19352, n22474);
  not g41444 (n_19353, n22475);
  and g41445 (n22476, n_19352, n_19353);
  and g41446 (n22477, n_19201, n_19205);
  and g41447 (n22478, n22476, n22477);
  not g41448 (n_19354, n22476);
  not g41449 (n_19355, n22477);
  and g41450 (n22479, n_19354, n_19355);
  not g41451 (n_19356, n22478);
  not g41452 (n_19357, n22479);
  and g41453 (n22480, n_19356, n_19357);
  and g41454 (n22481, n_19184, n_19197);
  and g41455 (n22482, \b[26] , n13903);
  and g41456 (n22483, \b[27] , n_11555);
  not g41457 (n_19358, n22482);
  not g41458 (n_19359, n22483);
  and g41459 (n22484, n_19358, n_19359);
  not g41460 (n_19360, n22484);
  and g41461 (n22485, n_2025, n_19360);
  and g41462 (n22486, \a[26] , n22484);
  not g41463 (n_19361, n22485);
  not g41464 (n_19362, n22486);
  and g41465 (n22487, n_19361, n_19362);
  and g41466 (n22488, n_19183, n22487);
  not g41467 (n_19363, n22487);
  and g41468 (n22489, n22293, n_19363);
  not g41469 (n_19364, n22488);
  not g41470 (n_19365, n22489);
  and g41471 (n22490, n_19364, n_19365);
  not g41472 (n_19366, n22481);
  and g41473 (n22491, n_19366, n22490);
  not g41474 (n_19367, n22490);
  and g41475 (n22492, n22481, n_19367);
  not g41476 (n_19368, n22491);
  not g41477 (n_19369, n22492);
  and g41478 (n22493, n_19368, n_19369);
  and g41479 (n22494, \b[30] , n12668);
  and g41480 (n22495, \b[28] , n13047);
  and g41481 (n22496, \b[29] , n12663);
  and g41487 (n22499, n3577, n12671);
  not g41490 (n_19374, n22500);
  and g41491 (n22501, \a[62] , n_19374);
  not g41492 (n_19375, n22501);
  and g41493 (n22502, \a[62] , n_19375);
  and g41494 (n22503, n_19374, n_19375);
  not g41495 (n_19376, n22502);
  not g41496 (n_19377, n22503);
  and g41497 (n22504, n_19376, n_19377);
  not g41498 (n_19378, n22504);
  and g41499 (n22505, n22493, n_19378);
  not g41500 (n_19379, n22505);
  and g41501 (n22506, n22493, n_19379);
  and g41502 (n22507, n_19378, n_19379);
  not g41503 (n_19380, n22506);
  not g41504 (n_19381, n22507);
  and g41505 (n22508, n_19380, n_19381);
  not g41506 (n_19382, n22480);
  and g41507 (n22509, n_19382, n22508);
  not g41508 (n_19383, n22508);
  and g41509 (n22510, n22480, n_19383);
  not g41510 (n_19384, n22509);
  not g41511 (n_19385, n22510);
  and g41512 (n22511, n_19384, n_19385);
  and g41513 (n22512, \b[36] , n10426);
  and g41514 (n22513, \b[34] , n10796);
  and g41515 (n22514, \b[35] , n10421);
  and g41521 (n22517, n4922, n10429);
  not g41524 (n_19390, n22518);
  and g41525 (n22519, \a[56] , n_19390);
  not g41526 (n_19391, n22519);
  and g41527 (n22520, \a[56] , n_19391);
  and g41528 (n22521, n_19390, n_19391);
  not g41529 (n_19392, n22520);
  not g41530 (n_19393, n22521);
  and g41531 (n22522, n_19392, n_19393);
  not g41532 (n_19394, n22522);
  and g41533 (n22523, n22511, n_19394);
  not g41534 (n_19395, n22523);
  and g41535 (n22524, n22511, n_19395);
  and g41536 (n22525, n_19394, n_19395);
  not g41537 (n_19396, n22524);
  not g41538 (n_19397, n22525);
  and g41539 (n22526, n_19396, n_19397);
  and g41540 (n22527, n_19209, n_19213);
  and g41541 (n22528, n22526, n22527);
  not g41542 (n_19398, n22526);
  not g41543 (n_19399, n22527);
  and g41544 (n22529, n_19398, n_19399);
  not g41545 (n_19400, n22528);
  not g41546 (n_19401, n22529);
  and g41547 (n22530, n_19400, n_19401);
  and g41548 (n22531, \b[39] , n9339);
  and g41549 (n22532, \b[37] , n9732);
  and g41550 (n22533, \b[38] , n9334);
  and g41556 (n22536, n5451, n9342);
  not g41559 (n_19406, n22537);
  and g41560 (n22538, \a[53] , n_19406);
  not g41561 (n_19407, n22538);
  and g41562 (n22539, \a[53] , n_19407);
  and g41563 (n22540, n_19406, n_19407);
  not g41564 (n_19408, n22539);
  not g41565 (n_19409, n22540);
  and g41566 (n22541, n_19408, n_19409);
  not g41567 (n_19410, n22541);
  and g41568 (n22542, n22530, n_19410);
  not g41569 (n_19411, n22542);
  and g41570 (n22543, n22530, n_19411);
  and g41571 (n22544, n_19410, n_19411);
  not g41572 (n_19412, n22543);
  not g41573 (n_19413, n22544);
  and g41574 (n22545, n_19412, n_19413);
  and g41575 (n22546, n_19217, n_19228);
  and g41576 (n22547, n22545, n22546);
  not g41577 (n_19414, n22545);
  not g41578 (n_19415, n22546);
  and g41579 (n22548, n_19414, n_19415);
  not g41580 (n_19416, n22547);
  not g41581 (n_19417, n22548);
  and g41582 (n22549, n_19416, n_19417);
  and g41583 (n22550, \b[42] , n8362);
  and g41584 (n22551, \b[40] , n8715);
  and g41585 (n22552, \b[41] , n8357);
  and g41591 (n22555, n6489, n8365);
  not g41594 (n_19422, n22556);
  and g41595 (n22557, \a[50] , n_19422);
  not g41596 (n_19423, n22557);
  and g41597 (n22558, \a[50] , n_19423);
  and g41598 (n22559, n_19422, n_19423);
  not g41599 (n_19424, n22558);
  not g41600 (n_19425, n22559);
  and g41601 (n22560, n_19424, n_19425);
  not g41602 (n_19426, n22560);
  and g41603 (n22561, n22549, n_19426);
  not g41604 (n_19427, n22561);
  and g41605 (n22562, n22549, n_19427);
  and g41606 (n22563, n_19426, n_19427);
  not g41607 (n_19428, n22562);
  not g41608 (n_19429, n22563);
  and g41609 (n22564, n_19428, n_19429);
  not g41610 (n_19430, n22465);
  and g41611 (n22565, n_19430, n22564);
  not g41612 (n_19431, n22564);
  and g41613 (n22566, n22465, n_19431);
  not g41614 (n_19432, n22565);
  not g41615 (n_19433, n22566);
  and g41616 (n22567, n_19432, n_19433);
  and g41617 (n22568, \b[45] , n7446);
  and g41618 (n22569, \b[43] , n7787);
  and g41619 (n22570, \b[44] , n7441);
  and g41625 (n22573, n7361, n7449);
  not g41628 (n_19438, n22574);
  and g41629 (n22575, \a[47] , n_19438);
  not g41630 (n_19439, n22575);
  and g41631 (n22576, \a[47] , n_19439);
  and g41632 (n22577, n_19438, n_19439);
  not g41633 (n_19440, n22576);
  not g41634 (n_19441, n22577);
  and g41635 (n22578, n_19440, n_19441);
  not g41636 (n_19442, n22567);
  not g41637 (n_19443, n22578);
  and g41638 (n22579, n_19442, n_19443);
  and g41639 (n22580, n22567, n22578);
  not g41640 (n_19444, n22579);
  not g41641 (n_19445, n22580);
  and g41642 (n22581, n_19444, n_19445);
  not g41643 (n_19446, n22581);
  and g41644 (n22582, n22463, n_19446);
  not g41645 (n_19447, n22463);
  and g41646 (n22583, n_19447, n22581);
  not g41647 (n_19448, n22582);
  not g41648 (n_19449, n22583);
  and g41649 (n22584, n_19448, n_19449);
  and g41650 (n22585, \b[48] , n6595);
  and g41651 (n22586, \b[46] , n6902);
  and g41652 (n22587, \b[47] , n6590);
  and g41658 (n22590, n6598, n8009);
  not g41661 (n_19454, n22591);
  and g41662 (n22592, \a[44] , n_19454);
  not g41663 (n_19455, n22592);
  and g41664 (n22593, \a[44] , n_19455);
  and g41665 (n22594, n_19454, n_19455);
  not g41666 (n_19456, n22593);
  not g41667 (n_19457, n22594);
  and g41668 (n22595, n_19456, n_19457);
  not g41669 (n_19458, n22595);
  and g41670 (n22596, n22584, n_19458);
  not g41671 (n_19459, n22596);
  and g41672 (n22597, n22584, n_19459);
  and g41673 (n22598, n_19458, n_19459);
  not g41674 (n_19460, n22597);
  not g41675 (n_19461, n22598);
  and g41676 (n22599, n_19460, n_19461);
  and g41677 (n22600, n_19258, n_19269);
  and g41678 (n22601, n22599, n22600);
  not g41679 (n_19462, n22599);
  not g41680 (n_19463, n22600);
  and g41681 (n22602, n_19462, n_19463);
  not g41682 (n_19464, n22601);
  not g41683 (n_19465, n22602);
  and g41684 (n22603, n_19464, n_19465);
  and g41685 (n22604, \b[51] , n5777);
  and g41686 (n22605, \b[49] , n6059);
  and g41687 (n22606, \b[50] , n5772);
  and g41693 (n22609, n5780, n8976);
  not g41696 (n_19470, n22610);
  and g41697 (n22611, \a[41] , n_19470);
  not g41698 (n_19471, n22611);
  and g41699 (n22612, \a[41] , n_19471);
  and g41700 (n22613, n_19470, n_19471);
  not g41701 (n_19472, n22612);
  not g41702 (n_19473, n22613);
  and g41703 (n22614, n_19472, n_19473);
  not g41704 (n_19474, n22614);
  and g41705 (n22615, n22603, n_19474);
  not g41706 (n_19475, n22603);
  and g41707 (n22616, n_19475, n22614);
  not g41708 (n_19476, n22462);
  not g41709 (n_19477, n22616);
  and g41710 (n22617, n_19476, n_19477);
  not g41711 (n_19478, n22615);
  and g41712 (n22618, n_19478, n22617);
  not g41713 (n_19479, n22618);
  and g41714 (n22619, n_19476, n_19479);
  and g41715 (n22620, n_19478, n_19479);
  and g41716 (n22621, n_19477, n22620);
  not g41717 (n_19480, n22619);
  not g41718 (n_19481, n22621);
  and g41719 (n22622, n_19480, n_19481);
  and g41720 (n22623, \b[54] , n5035);
  and g41721 (n22624, \b[52] , n5277);
  and g41722 (n22625, \b[53] , n5030);
  and g41728 (n22628, n5038, n9998);
  not g41731 (n_19486, n22629);
  and g41732 (n22630, \a[38] , n_19486);
  not g41733 (n_19487, n22630);
  and g41734 (n22631, \a[38] , n_19487);
  and g41735 (n22632, n_19486, n_19487);
  not g41736 (n_19488, n22631);
  not g41737 (n_19489, n22632);
  and g41738 (n22633, n_19488, n_19489);
  and g41739 (n22634, n22622, n22633);
  not g41740 (n_19490, n22622);
  not g41741 (n_19491, n22633);
  and g41742 (n22635, n_19490, n_19491);
  not g41743 (n_19492, n22634);
  not g41744 (n_19493, n22635);
  and g41745 (n22636, n_19492, n_19493);
  not g41746 (n_19494, n22461);
  and g41747 (n22637, n_19494, n22636);
  not g41748 (n_19495, n22636);
  and g41749 (n22638, n22461, n_19495);
  not g41750 (n_19496, n22637);
  not g41751 (n_19497, n22638);
  and g41752 (n22639, n_19496, n_19497);
  not g41753 (n_19498, n22460);
  and g41754 (n22640, n_19498, n22639);
  not g41755 (n_19499, n22640);
  and g41756 (n22641, n22639, n_19499);
  and g41757 (n22642, n_19498, n_19499);
  not g41758 (n_19500, n22641);
  not g41759 (n_19501, n22642);
  and g41760 (n22643, n_19500, n_19501);
  and g41761 (n22644, n_19298, n_19301);
  and g41762 (n22645, n22643, n22644);
  not g41763 (n_19502, n22643);
  not g41764 (n_19503, n22644);
  and g41765 (n22646, n_19502, n_19503);
  not g41766 (n_19504, n22645);
  not g41767 (n_19505, n22646);
  and g41768 (n22647, n_19504, n_19505);
  and g41769 (n22648, \b[60] , n3638);
  and g41770 (n22649, \b[58] , n3843);
  and g41771 (n22650, \b[59] , n3633);
  and g41777 (n22653, n3641, n12211);
  not g41780 (n_19510, n22654);
  and g41781 (n22655, \a[32] , n_19510);
  not g41782 (n_19511, n22655);
  and g41783 (n22656, \a[32] , n_19511);
  and g41784 (n22657, n_19510, n_19511);
  not g41785 (n_19512, n22656);
  not g41786 (n_19513, n22657);
  and g41787 (n22658, n_19512, n_19513);
  and g41788 (n22659, n_19140, n_19305);
  and g41789 (n22660, n22658, n22659);
  not g41790 (n_19514, n22658);
  not g41791 (n_19515, n22659);
  and g41792 (n22661, n_19514, n_19515);
  not g41793 (n_19516, n22660);
  not g41794 (n_19517, n22661);
  and g41795 (n22662, n_19516, n_19517);
  not g41796 (n_19518, n22662);
  and g41797 (n22663, n22647, n_19518);
  not g41798 (n_19519, n22647);
  and g41799 (n22664, n_19519, n22662);
  not g41800 (n_19520, n22663);
  not g41801 (n_19521, n22664);
  and g41802 (n22665, n_19520, n_19521);
  not g41803 (n_19522, n22449);
  not g41804 (n_19523, n22665);
  and g41805 (n22666, n_19522, n_19523);
  and g41806 (n22667, n22449, n22665);
  not g41807 (n_19524, n22666);
  not g41808 (n_19525, n22667);
  and g41809 (n22668, n_19524, n_19525);
  not g41810 (n_19526, n22668);
  and g41811 (n22669, n22433, n_19526);
  not g41812 (n_19527, n22433);
  and g41813 (n22670, n_19527, n22668);
  not g41814 (n_19528, n22669);
  not g41815 (n_19529, n22670);
  and g41816 (n22671, n_19528, n_19529);
  and g41817 (n22672, n_19318, n_19322);
  not g41818 (n_19530, n22672);
  and g41819 (n22673, n22671, n_19530);
  not g41820 (n_19531, n22671);
  and g41821 (n22674, n_19531, n22672);
  not g41822 (n_19532, n22673);
  not g41823 (n_19533, n22674);
  and g41824 (\f[90] , n_19532, n_19533);
  and g41825 (n22676, n22647, n22662);
  not g41826 (n_19534, n22676);
  and g41827 (n22677, n_19517, n_19534);
  and g41828 (n22678, \b[62] , n3243);
  and g41829 (n22679, \b[63] , n3045);
  not g41830 (n_19535, n22678);
  not g41831 (n_19536, n22679);
  and g41832 (n22680, n_19535, n_19536);
  and g41833 (n22681, n_12601, n22680);
  and g41834 (n22682, n13800, n22680);
  not g41835 (n_19537, n22681);
  not g41836 (n_19538, n22682);
  and g41837 (n22683, n_19537, n_19538);
  not g41838 (n_19539, n22683);
  and g41839 (n22684, \a[29] , n_19539);
  and g41840 (n22685, n_2476, n22683);
  not g41841 (n_19540, n22684);
  not g41842 (n_19541, n22685);
  and g41843 (n22686, n_19540, n_19541);
  not g41844 (n_19542, n22677);
  not g41845 (n_19543, n22686);
  and g41846 (n22687, n_19542, n_19543);
  and g41847 (n22688, n22677, n22686);
  not g41848 (n_19544, n22687);
  not g41849 (n_19545, n22688);
  and g41850 (n22689, n_19544, n_19545);
  and g41851 (n22690, \b[61] , n3638);
  and g41852 (n22691, \b[59] , n3843);
  and g41853 (n22692, \b[60] , n3633);
  and g41859 (n22695, n3641, n12969);
  not g41862 (n_19550, n22696);
  and g41863 (n22697, \a[32] , n_19550);
  not g41864 (n_19551, n22697);
  and g41865 (n22698, \a[32] , n_19551);
  and g41866 (n22699, n_19550, n_19551);
  not g41867 (n_19552, n22698);
  not g41868 (n_19553, n22699);
  and g41869 (n22700, n_19552, n_19553);
  and g41870 (n22701, n_19499, n_19505);
  and g41871 (n22702, n22700, n22701);
  not g41872 (n_19554, n22700);
  not g41873 (n_19555, n22701);
  and g41874 (n22703, n_19554, n_19555);
  not g41875 (n_19556, n22702);
  not g41876 (n_19557, n22703);
  and g41877 (n22704, n_19556, n_19557);
  and g41878 (n22705, \b[58] , n4287);
  and g41879 (n22706, \b[56] , n4532);
  and g41880 (n22707, \b[57] , n4282);
  and g41886 (n22710, n4290, n11436);
  not g41889 (n_19562, n22711);
  and g41890 (n22712, \a[35] , n_19562);
  not g41891 (n_19563, n22712);
  and g41892 (n22713, \a[35] , n_19563);
  and g41893 (n22714, n_19562, n_19563);
  not g41894 (n_19564, n22713);
  not g41895 (n_19565, n22714);
  and g41896 (n22715, n_19564, n_19565);
  and g41897 (n22716, n_19493, n_19496);
  and g41898 (n22717, \b[43] , n8362);
  and g41899 (n22718, \b[41] , n8715);
  and g41900 (n22719, \b[42] , n8357);
  and g41906 (n22722, n6515, n8365);
  not g41909 (n_19570, n22723);
  and g41910 (n22724, \a[50] , n_19570);
  not g41911 (n_19571, n22724);
  and g41912 (n22725, \a[50] , n_19571);
  and g41913 (n22726, n_19570, n_19571);
  not g41914 (n_19572, n22725);
  not g41915 (n_19573, n22726);
  and g41916 (n22727, n_19572, n_19573);
  and g41917 (n22728, n_19411, n_19417);
  and g41918 (n22729, \b[40] , n9339);
  and g41919 (n22730, \b[38] , n9732);
  and g41920 (n22731, \b[39] , n9334);
  and g41926 (n22734, n5955, n9342);
  not g41929 (n_19578, n22735);
  and g41930 (n22736, \a[53] , n_19578);
  not g41931 (n_19579, n22736);
  and g41932 (n22737, \a[53] , n_19579);
  and g41933 (n22738, n_19578, n_19579);
  not g41934 (n_19580, n22737);
  not g41935 (n_19581, n22738);
  and g41936 (n22739, n_19580, n_19581);
  and g41937 (n22740, n_19395, n_19401);
  and g41938 (n22741, \b[34] , n11531);
  and g41939 (n22742, \b[32] , n11896);
  and g41940 (n22743, \b[33] , n11526);
  and g41946 (n22746, n4466, n11534);
  not g41949 (n_19586, n22747);
  and g41950 (n22748, \a[59] , n_19586);
  not g41951 (n_19587, n22748);
  and g41952 (n22749, \a[59] , n_19587);
  and g41953 (n22750, n_19586, n_19587);
  not g41954 (n_19588, n22749);
  not g41955 (n_19589, n22750);
  and g41956 (n22751, n_19588, n_19589);
  and g41957 (n22752, \b[27] , n13903);
  and g41958 (n22753, \b[28] , n_11555);
  not g41959 (n_19590, n22752);
  not g41960 (n_19591, n22753);
  and g41961 (n22754, n_19590, n_19591);
  and g41962 (n22755, n_19361, n_19364);
  not g41963 (n_19592, n22754);
  and g41964 (n22756, n_19592, n22755);
  not g41965 (n_19593, n22755);
  and g41966 (n22757, n22754, n_19593);
  not g41967 (n_19594, n22756);
  not g41968 (n_19595, n22757);
  and g41969 (n22758, n_19594, n_19595);
  and g41970 (n22759, \b[31] , n12668);
  and g41971 (n22760, \b[29] , n13047);
  and g41972 (n22761, \b[30] , n12663);
  and g41978 (n22764, n3796, n12671);
  not g41981 (n_19600, n22765);
  and g41982 (n22766, \a[62] , n_19600);
  not g41983 (n_19601, n22766);
  and g41984 (n22767, \a[62] , n_19601);
  and g41985 (n22768, n_19600, n_19601);
  not g41986 (n_19602, n22767);
  not g41987 (n_19603, n22768);
  and g41988 (n22769, n_19602, n_19603);
  not g41989 (n_19604, n22758);
  and g41990 (n22770, n_19604, n22769);
  not g41991 (n_19605, n22769);
  and g41992 (n22771, n22758, n_19605);
  not g41993 (n_19606, n22770);
  not g41994 (n_19607, n22771);
  and g41995 (n22772, n_19606, n_19607);
  and g41996 (n22773, n_19368, n_19379);
  not g41997 (n_19608, n22773);
  and g41998 (n22774, n22772, n_19608);
  not g41999 (n_19609, n22772);
  and g42000 (n22775, n_19609, n22773);
  not g42001 (n_19610, n22774);
  not g42002 (n_19611, n22775);
  and g42003 (n22776, n_19610, n_19611);
  not g42004 (n_19612, n22751);
  and g42005 (n22777, n_19612, n22776);
  not g42006 (n_19613, n22777);
  and g42007 (n22778, n22776, n_19613);
  and g42008 (n22779, n_19612, n_19613);
  not g42009 (n_19614, n22778);
  not g42010 (n_19615, n22779);
  and g42011 (n22780, n_19614, n_19615);
  and g42012 (n22781, n_19357, n_19385);
  not g42013 (n_19616, n22780);
  not g42014 (n_19617, n22781);
  and g42015 (n22782, n_19616, n_19617);
  not g42016 (n_19618, n22782);
  and g42017 (n22783, n_19616, n_19618);
  and g42018 (n22784, n_19617, n_19618);
  not g42019 (n_19619, n22783);
  not g42020 (n_19620, n22784);
  and g42021 (n22785, n_19619, n_19620);
  and g42022 (n22786, \b[37] , n10426);
  and g42023 (n22787, \b[35] , n10796);
  and g42024 (n22788, \b[36] , n10421);
  and g42030 (n22791, n5181, n10429);
  not g42033 (n_19625, n22792);
  and g42034 (n22793, \a[56] , n_19625);
  not g42035 (n_19626, n22793);
  and g42036 (n22794, \a[56] , n_19626);
  and g42037 (n22795, n_19625, n_19626);
  not g42038 (n_19627, n22794);
  not g42039 (n_19628, n22795);
  and g42040 (n22796, n_19627, n_19628);
  not g42041 (n_19629, n22785);
  and g42042 (n22797, n_19629, n22796);
  not g42043 (n_19630, n22796);
  and g42044 (n22798, n22785, n_19630);
  not g42045 (n_19631, n22797);
  not g42046 (n_19632, n22798);
  and g42047 (n22799, n_19631, n_19632);
  not g42048 (n_19633, n22740);
  not g42049 (n_19634, n22799);
  and g42050 (n22800, n_19633, n_19634);
  not g42051 (n_19635, n22800);
  and g42052 (n22801, n_19633, n_19635);
  and g42053 (n22802, n_19634, n_19635);
  not g42054 (n_19636, n22801);
  not g42055 (n_19637, n22802);
  and g42056 (n22803, n_19636, n_19637);
  not g42057 (n_19638, n22739);
  not g42058 (n_19639, n22803);
  and g42059 (n22804, n_19638, n_19639);
  and g42060 (n22805, n22739, n_19637);
  and g42061 (n22806, n_19636, n22805);
  not g42062 (n_19640, n22804);
  not g42063 (n_19641, n22806);
  and g42064 (n22807, n_19640, n_19641);
  not g42065 (n_19642, n22728);
  and g42066 (n22808, n_19642, n22807);
  not g42067 (n_19643, n22807);
  and g42068 (n22809, n22728, n_19643);
  not g42069 (n_19644, n22808);
  not g42070 (n_19645, n22809);
  and g42071 (n22810, n_19644, n_19645);
  not g42072 (n_19646, n22727);
  and g42073 (n22811, n_19646, n22810);
  not g42074 (n_19647, n22811);
  and g42075 (n22812, n22810, n_19647);
  and g42076 (n22813, n_19646, n_19647);
  not g42077 (n_19648, n22812);
  not g42078 (n_19649, n22813);
  and g42079 (n22814, n_19648, n_19649);
  and g42080 (n22815, n_19430, n_19431);
  not g42081 (n_19650, n22815);
  and g42082 (n22816, n_19427, n_19650);
  and g42083 (n22817, n22814, n22816);
  not g42084 (n_19651, n22814);
  not g42085 (n_19652, n22816);
  and g42086 (n22818, n_19651, n_19652);
  not g42087 (n_19653, n22817);
  not g42088 (n_19654, n22818);
  and g42089 (n22819, n_19653, n_19654);
  and g42090 (n22820, \b[46] , n7446);
  and g42091 (n22821, \b[44] , n7787);
  and g42092 (n22822, \b[45] , n7441);
  and g42098 (n22825, n7449, n7677);
  not g42101 (n_19659, n22826);
  and g42102 (n22827, \a[47] , n_19659);
  not g42103 (n_19660, n22827);
  and g42104 (n22828, \a[47] , n_19660);
  and g42105 (n22829, n_19659, n_19660);
  not g42106 (n_19661, n22828);
  not g42107 (n_19662, n22829);
  and g42108 (n22830, n_19661, n_19662);
  not g42109 (n_19663, n22830);
  and g42110 (n22831, n22819, n_19663);
  not g42111 (n_19664, n22831);
  and g42112 (n22832, n22819, n_19664);
  and g42113 (n22833, n_19663, n_19664);
  not g42114 (n_19665, n22832);
  not g42115 (n_19666, n22833);
  and g42116 (n22834, n_19665, n_19666);
  and g42117 (n22835, n_19444, n_19449);
  and g42118 (n22836, n22834, n22835);
  not g42119 (n_19667, n22834);
  not g42120 (n_19668, n22835);
  and g42121 (n22837, n_19667, n_19668);
  not g42122 (n_19669, n22836);
  not g42123 (n_19670, n22837);
  and g42124 (n22838, n_19669, n_19670);
  and g42125 (n22839, \b[49] , n6595);
  and g42126 (n22840, \b[47] , n6902);
  and g42127 (n22841, \b[48] , n6590);
  and g42133 (n22844, n6598, n8625);
  not g42136 (n_19675, n22845);
  and g42137 (n22846, \a[44] , n_19675);
  not g42138 (n_19676, n22846);
  and g42139 (n22847, \a[44] , n_19676);
  and g42140 (n22848, n_19675, n_19676);
  not g42141 (n_19677, n22847);
  not g42142 (n_19678, n22848);
  and g42143 (n22849, n_19677, n_19678);
  not g42144 (n_19679, n22849);
  and g42145 (n22850, n22838, n_19679);
  not g42146 (n_19680, n22850);
  and g42147 (n22851, n22838, n_19680);
  and g42148 (n22852, n_19679, n_19680);
  not g42149 (n_19681, n22851);
  not g42150 (n_19682, n22852);
  and g42151 (n22853, n_19681, n_19682);
  and g42152 (n22854, n_19459, n_19465);
  and g42153 (n22855, n22853, n22854);
  not g42154 (n_19683, n22853);
  not g42155 (n_19684, n22854);
  and g42156 (n22856, n_19683, n_19684);
  not g42157 (n_19685, n22855);
  not g42158 (n_19686, n22856);
  and g42159 (n22857, n_19685, n_19686);
  and g42160 (n22858, \b[52] , n5777);
  and g42161 (n22859, \b[50] , n6059);
  and g42162 (n22860, \b[51] , n5772);
  and g42168 (n22863, n5780, n9628);
  not g42171 (n_19691, n22864);
  and g42172 (n22865, \a[41] , n_19691);
  not g42173 (n_19692, n22865);
  and g42174 (n22866, \a[41] , n_19692);
  and g42175 (n22867, n_19691, n_19692);
  not g42176 (n_19693, n22866);
  not g42177 (n_19694, n22867);
  and g42178 (n22868, n_19693, n_19694);
  not g42179 (n_19695, n22868);
  and g42180 (n22869, n22857, n_19695);
  not g42181 (n_19696, n22869);
  and g42182 (n22870, n22857, n_19696);
  and g42183 (n22871, n_19695, n_19696);
  not g42184 (n_19697, n22870);
  not g42185 (n_19698, n22871);
  and g42186 (n22872, n_19697, n_19698);
  not g42187 (n_19699, n22620);
  and g42188 (n22873, n_19699, n22872);
  not g42189 (n_19700, n22872);
  and g42190 (n22874, n22620, n_19700);
  not g42191 (n_19701, n22873);
  not g42192 (n_19702, n22874);
  and g42193 (n22875, n_19701, n_19702);
  and g42194 (n22876, \b[55] , n5035);
  and g42195 (n22877, \b[53] , n5277);
  and g42196 (n22878, \b[54] , n5030);
  and g42202 (n22881, n5038, n10684);
  not g42205 (n_19707, n22882);
  and g42206 (n22883, \a[38] , n_19707);
  not g42207 (n_19708, n22883);
  and g42208 (n22884, \a[38] , n_19708);
  and g42209 (n22885, n_19707, n_19708);
  not g42210 (n_19709, n22884);
  not g42211 (n_19710, n22885);
  and g42212 (n22886, n_19709, n_19710);
  not g42213 (n_19711, n22875);
  not g42214 (n_19712, n22886);
  and g42215 (n22887, n_19711, n_19712);
  and g42216 (n22888, n22875, n22886);
  not g42217 (n_19713, n22887);
  not g42218 (n_19714, n22888);
  and g42219 (n22889, n_19713, n_19714);
  not g42220 (n_19715, n22716);
  and g42221 (n22890, n_19715, n22889);
  not g42222 (n_19716, n22889);
  and g42223 (n22891, n22716, n_19716);
  not g42224 (n_19717, n22890);
  not g42225 (n_19718, n22891);
  and g42226 (n22892, n_19717, n_19718);
  not g42227 (n_19719, n22715);
  and g42228 (n22893, n_19719, n22892);
  not g42229 (n_19720, n22893);
  and g42230 (n22894, n22892, n_19720);
  and g42231 (n22895, n_19719, n_19720);
  not g42232 (n_19721, n22894);
  not g42233 (n_19722, n22895);
  and g42234 (n22896, n_19721, n_19722);
  not g42235 (n_19723, n22896);
  and g42236 (n22897, n22704, n_19723);
  not g42237 (n_19724, n22704);
  and g42238 (n22898, n_19724, n22896);
  not g42239 (n_19725, n22898);
  and g42240 (n22899, n22689, n_19725);
  not g42241 (n_19726, n22897);
  and g42242 (n22900, n_19726, n22899);
  not g42243 (n_19727, n22900);
  and g42244 (n22901, n22689, n_19727);
  and g42245 (n22902, n_19725, n_19727);
  and g42246 (n22903, n_19726, n22902);
  not g42247 (n_19728, n22901);
  not g42248 (n_19729, n22903);
  and g42249 (n22904, n_19728, n_19729);
  and g42250 (n22905, n_19334, n_19524);
  and g42251 (n22906, n22904, n22905);
  not g42252 (n_19730, n22904);
  not g42253 (n_19731, n22905);
  and g42254 (n22907, n_19730, n_19731);
  not g42255 (n_19732, n22906);
  not g42256 (n_19733, n22907);
  and g42257 (n22908, n_19732, n_19733);
  and g42258 (n22909, n_19529, n_19532);
  not g42259 (n_19734, n22909);
  and g42260 (n22910, n22908, n_19734);
  not g42261 (n_19735, n22908);
  and g42262 (n22911, n_19735, n22909);
  not g42263 (n_19736, n22910);
  not g42264 (n_19737, n22911);
  and g42265 (\f[91] , n_19736, n_19737);
  and g42266 (n22913, n_19733, n_19736);
  and g42267 (n22914, n_19544, n_19727);
  and g42268 (n22915, n_19557, n_19726);
  and g42269 (n22916, \b[63] , n3243);
  and g42270 (n22917, n3053, n13797);
  not g42271 (n_19738, n22916);
  not g42272 (n_19739, n22917);
  and g42273 (n22918, n_19738, n_19739);
  not g42274 (n_19740, n22918);
  and g42275 (n22919, \a[29] , n_19740);
  not g42276 (n_19741, n22919);
  and g42277 (n22920, \a[29] , n_19741);
  and g42278 (n22921, n_19740, n_19741);
  not g42279 (n_19742, n22920);
  not g42280 (n_19743, n22921);
  and g42281 (n22922, n_19742, n_19743);
  not g42282 (n_19744, n22915);
  not g42283 (n_19745, n22922);
  and g42284 (n22923, n_19744, n_19745);
  not g42285 (n_19746, n22923);
  and g42286 (n22924, n_19744, n_19746);
  and g42287 (n22925, n_19745, n_19746);
  not g42288 (n_19747, n22924);
  not g42289 (n_19748, n22925);
  and g42290 (n22926, n_19747, n_19748);
  and g42291 (n22927, \b[62] , n3638);
  and g42292 (n22928, \b[60] , n3843);
  and g42293 (n22929, \b[61] , n3633);
  and g42299 (n22932, n3641, n13370);
  not g42302 (n_19753, n22933);
  and g42303 (n22934, \a[32] , n_19753);
  not g42304 (n_19754, n22934);
  and g42305 (n22935, \a[32] , n_19754);
  and g42306 (n22936, n_19753, n_19754);
  not g42307 (n_19755, n22935);
  not g42308 (n_19756, n22936);
  and g42309 (n22937, n_19755, n_19756);
  and g42310 (n22938, n_19717, n_19720);
  and g42311 (n22939, n22937, n22938);
  not g42312 (n_19757, n22937);
  not g42313 (n_19758, n22938);
  and g42314 (n22940, n_19757, n_19758);
  not g42315 (n_19759, n22939);
  not g42316 (n_19760, n22940);
  and g42317 (n22941, n_19759, n_19760);
  and g42318 (n22942, n_19699, n_19700);
  not g42319 (n_19761, n22942);
  and g42320 (n22943, n_19713, n_19761);
  and g42321 (n22944, \b[56] , n5035);
  and g42322 (n22945, \b[54] , n5277);
  and g42323 (n22946, \b[55] , n5030);
  and g42329 (n22949, n5038, n10708);
  not g42332 (n_19766, n22950);
  and g42333 (n22951, \a[38] , n_19766);
  not g42334 (n_19767, n22951);
  and g42335 (n22952, \a[38] , n_19767);
  and g42336 (n22953, n_19766, n_19767);
  not g42337 (n_19768, n22952);
  not g42338 (n_19769, n22953);
  and g42339 (n22954, n_19768, n_19769);
  and g42340 (n22955, n_19686, n_19696);
  and g42341 (n22956, \b[53] , n5777);
  and g42342 (n22957, \b[51] , n6059);
  and g42343 (n22958, \b[52] , n5772);
  and g42349 (n22961, n5780, n9972);
  not g42352 (n_19774, n22962);
  and g42353 (n22963, \a[41] , n_19774);
  not g42354 (n_19775, n22963);
  and g42355 (n22964, \a[41] , n_19775);
  and g42356 (n22965, n_19774, n_19775);
  not g42357 (n_19776, n22964);
  not g42358 (n_19777, n22965);
  and g42359 (n22966, n_19776, n_19777);
  and g42360 (n22967, n_19670, n_19680);
  and g42361 (n22968, n_19644, n_19647);
  and g42362 (n22969, \b[44] , n8362);
  and g42363 (n22970, \b[42] , n8715);
  and g42364 (n22971, \b[43] , n8357);
  and g42370 (n22974, n7072, n8365);
  not g42373 (n_19782, n22975);
  and g42374 (n22976, \a[50] , n_19782);
  not g42375 (n_19783, n22976);
  and g42376 (n22977, \a[50] , n_19783);
  and g42377 (n22978, n_19782, n_19783);
  not g42378 (n_19784, n22977);
  not g42379 (n_19785, n22978);
  and g42380 (n22979, n_19784, n_19785);
  and g42381 (n22980, n_19635, n_19640);
  and g42382 (n22981, n_19610, n_19613);
  and g42383 (n22982, \b[35] , n11531);
  and g42384 (n22983, \b[33] , n11896);
  and g42385 (n22984, \b[34] , n11526);
  and g42391 (n22987, n4696, n11534);
  not g42394 (n_19790, n22988);
  and g42395 (n22989, \a[59] , n_19790);
  not g42396 (n_19791, n22989);
  and g42397 (n22990, \a[59] , n_19791);
  and g42398 (n22991, n_19790, n_19791);
  not g42399 (n_19792, n22990);
  not g42400 (n_19793, n22991);
  and g42401 (n22992, n_19792, n_19793);
  and g42402 (n22993, n_19595, n_19607);
  and g42403 (n22994, \b[28] , n13903);
  and g42404 (n22995, \b[29] , n_11555);
  not g42405 (n_19794, n22994);
  not g42406 (n_19795, n22995);
  and g42407 (n22996, n_19794, n_19795);
  not g42408 (n_19796, n22996);
  and g42409 (n22997, n22754, n_19796);
  and g42410 (n22998, n_19592, n22996);
  not g42411 (n_19797, n22993);
  not g42412 (n_19798, n22998);
  and g42413 (n22999, n_19797, n_19798);
  not g42414 (n_19799, n22997);
  and g42415 (n23000, n_19799, n22999);
  not g42416 (n_19800, n23000);
  and g42417 (n23001, n_19797, n_19800);
  and g42418 (n23002, n_19798, n_19800);
  and g42419 (n23003, n_19799, n23002);
  not g42420 (n_19801, n23001);
  not g42421 (n_19802, n23003);
  and g42422 (n23004, n_19801, n_19802);
  and g42423 (n23005, \b[32] , n12668);
  and g42424 (n23006, \b[30] , n13047);
  and g42425 (n23007, \b[31] , n12663);
  and g42431 (n23010, n4013, n12671);
  not g42434 (n_19807, n23011);
  and g42435 (n23012, \a[62] , n_19807);
  not g42436 (n_19808, n23012);
  and g42437 (n23013, \a[62] , n_19808);
  and g42438 (n23014, n_19807, n_19808);
  not g42439 (n_19809, n23013);
  not g42440 (n_19810, n23014);
  and g42441 (n23015, n_19809, n_19810);
  not g42442 (n_19811, n23004);
  and g42443 (n23016, n_19811, n23015);
  not g42444 (n_19812, n23015);
  and g42445 (n23017, n23004, n_19812);
  not g42446 (n_19813, n23016);
  not g42447 (n_19814, n23017);
  and g42448 (n23018, n_19813, n_19814);
  not g42449 (n_19815, n22992);
  not g42450 (n_19816, n23018);
  and g42451 (n23019, n_19815, n_19816);
  and g42452 (n23020, n22992, n23018);
  not g42453 (n_19817, n23019);
  not g42454 (n_19818, n23020);
  and g42455 (n23021, n_19817, n_19818);
  not g42456 (n_19819, n22981);
  and g42457 (n23022, n_19819, n23021);
  not g42458 (n_19820, n23021);
  and g42459 (n23023, n22981, n_19820);
  not g42460 (n_19821, n23022);
  not g42461 (n_19822, n23023);
  and g42462 (n23024, n_19821, n_19822);
  and g42463 (n23025, \b[38] , n10426);
  and g42464 (n23026, \b[36] , n10796);
  and g42465 (n23027, \b[37] , n10421);
  and g42471 (n23030, n5205, n10429);
  not g42474 (n_19827, n23031);
  and g42475 (n23032, \a[56] , n_19827);
  not g42476 (n_19828, n23032);
  and g42477 (n23033, \a[56] , n_19828);
  and g42478 (n23034, n_19827, n_19828);
  not g42479 (n_19829, n23033);
  not g42480 (n_19830, n23034);
  and g42481 (n23035, n_19829, n_19830);
  not g42482 (n_19831, n23035);
  and g42483 (n23036, n23024, n_19831);
  not g42484 (n_19832, n23036);
  and g42485 (n23037, n23024, n_19832);
  and g42486 (n23038, n_19831, n_19832);
  not g42487 (n_19833, n23037);
  not g42488 (n_19834, n23038);
  and g42489 (n23039, n_19833, n_19834);
  and g42490 (n23040, n_19629, n_19630);
  not g42491 (n_19835, n23040);
  and g42492 (n23041, n_19618, n_19835);
  not g42493 (n_19836, n23039);
  not g42494 (n_19837, n23041);
  and g42495 (n23042, n_19836, n_19837);
  not g42496 (n_19838, n23042);
  and g42497 (n23043, n_19836, n_19838);
  and g42498 (n23044, n_19837, n_19838);
  not g42499 (n_19839, n23043);
  not g42500 (n_19840, n23044);
  and g42501 (n23045, n_19839, n_19840);
  and g42502 (n23046, \b[41] , n9339);
  and g42503 (n23047, \b[39] , n9732);
  and g42504 (n23048, \b[40] , n9334);
  and g42510 (n23051, n6219, n9342);
  not g42513 (n_19845, n23052);
  and g42514 (n23053, \a[53] , n_19845);
  not g42515 (n_19846, n23053);
  and g42516 (n23054, \a[53] , n_19846);
  and g42517 (n23055, n_19845, n_19846);
  not g42518 (n_19847, n23054);
  not g42519 (n_19848, n23055);
  and g42520 (n23056, n_19847, n_19848);
  not g42521 (n_19849, n23045);
  and g42522 (n23057, n_19849, n23056);
  not g42523 (n_19850, n23056);
  and g42524 (n23058, n23045, n_19850);
  not g42525 (n_19851, n23057);
  not g42526 (n_19852, n23058);
  and g42527 (n23059, n_19851, n_19852);
  not g42528 (n_19853, n22980);
  not g42529 (n_19854, n23059);
  and g42530 (n23060, n_19853, n_19854);
  and g42531 (n23061, n22980, n23059);
  not g42532 (n_19855, n23060);
  not g42533 (n_19856, n23061);
  and g42534 (n23062, n_19855, n_19856);
  not g42535 (n_19857, n22979);
  and g42536 (n23063, n_19857, n23062);
  not g42537 (n_19858, n23062);
  and g42538 (n23064, n22979, n_19858);
  not g42539 (n_19859, n23063);
  not g42540 (n_19860, n23064);
  and g42541 (n23065, n_19859, n_19860);
  not g42542 (n_19861, n22968);
  and g42543 (n23066, n_19861, n23065);
  not g42544 (n_19862, n23065);
  and g42545 (n23067, n22968, n_19862);
  not g42546 (n_19863, n23066);
  not g42547 (n_19864, n23067);
  and g42548 (n23068, n_19863, n_19864);
  and g42549 (n23069, \b[47] , n7446);
  and g42550 (n23070, \b[45] , n7787);
  and g42551 (n23071, \b[46] , n7441);
  and g42557 (n23074, n7449, n7703);
  not g42560 (n_19869, n23075);
  and g42561 (n23076, \a[47] , n_19869);
  not g42562 (n_19870, n23076);
  and g42563 (n23077, \a[47] , n_19870);
  and g42564 (n23078, n_19869, n_19870);
  not g42565 (n_19871, n23077);
  not g42566 (n_19872, n23078);
  and g42567 (n23079, n_19871, n_19872);
  not g42568 (n_19873, n23079);
  and g42569 (n23080, n23068, n_19873);
  not g42570 (n_19874, n23080);
  and g42571 (n23081, n23068, n_19874);
  and g42572 (n23082, n_19873, n_19874);
  not g42573 (n_19875, n23081);
  not g42574 (n_19876, n23082);
  and g42575 (n23083, n_19875, n_19876);
  and g42576 (n23084, n_19654, n_19664);
  and g42577 (n23085, n23083, n23084);
  not g42578 (n_19877, n23083);
  not g42579 (n_19878, n23084);
  and g42580 (n23086, n_19877, n_19878);
  not g42581 (n_19879, n23085);
  not g42582 (n_19880, n23086);
  and g42583 (n23087, n_19879, n_19880);
  and g42584 (n23088, \b[50] , n6595);
  and g42585 (n23089, \b[48] , n6902);
  and g42586 (n23090, \b[49] , n6590);
  and g42592 (n23093, n6598, n8949);
  not g42595 (n_19885, n23094);
  and g42596 (n23095, \a[44] , n_19885);
  not g42597 (n_19886, n23095);
  and g42598 (n23096, \a[44] , n_19886);
  and g42599 (n23097, n_19885, n_19886);
  not g42600 (n_19887, n23096);
  not g42601 (n_19888, n23097);
  and g42602 (n23098, n_19887, n_19888);
  not g42603 (n_19889, n23087);
  and g42604 (n23099, n_19889, n23098);
  not g42605 (n_19890, n23098);
  and g42606 (n23100, n23087, n_19890);
  not g42607 (n_19891, n23099);
  not g42608 (n_19892, n23100);
  and g42609 (n23101, n_19891, n_19892);
  not g42610 (n_19893, n22967);
  and g42611 (n23102, n_19893, n23101);
  not g42612 (n_19894, n23102);
  and g42613 (n23103, n_19893, n_19894);
  and g42614 (n23104, n23101, n_19894);
  not g42615 (n_19895, n23103);
  not g42616 (n_19896, n23104);
  and g42617 (n23105, n_19895, n_19896);
  not g42618 (n_19897, n22966);
  not g42619 (n_19898, n23105);
  and g42620 (n23106, n_19897, n_19898);
  and g42621 (n23107, n22966, n_19896);
  and g42622 (n23108, n_19895, n23107);
  not g42623 (n_19899, n23106);
  not g42624 (n_19900, n23108);
  and g42625 (n23109, n_19899, n_19900);
  not g42626 (n_19901, n22955);
  and g42627 (n23110, n_19901, n23109);
  not g42628 (n_19902, n23109);
  and g42629 (n23111, n22955, n_19902);
  not g42630 (n_19903, n23110);
  not g42631 (n_19904, n23111);
  and g42632 (n23112, n_19903, n_19904);
  not g42633 (n_19905, n22954);
  and g42634 (n23113, n_19905, n23112);
  not g42635 (n_19906, n23112);
  and g42636 (n23114, n22954, n_19906);
  not g42637 (n_19907, n23113);
  not g42638 (n_19908, n23114);
  and g42639 (n23115, n_19907, n_19908);
  not g42640 (n_19909, n22943);
  and g42641 (n23116, n_19909, n23115);
  not g42642 (n_19910, n23115);
  and g42643 (n23117, n22943, n_19910);
  not g42644 (n_19911, n23116);
  not g42645 (n_19912, n23117);
  and g42646 (n23118, n_19911, n_19912);
  and g42647 (n23119, \b[59] , n4287);
  and g42648 (n23120, \b[57] , n4532);
  and g42649 (n23121, \b[58] , n4282);
  and g42655 (n23124, n4290, n12179);
  not g42658 (n_19917, n23125);
  and g42659 (n23126, \a[35] , n_19917);
  not g42660 (n_19918, n23126);
  and g42661 (n23127, \a[35] , n_19918);
  and g42662 (n23128, n_19917, n_19918);
  not g42663 (n_19919, n23127);
  not g42664 (n_19920, n23128);
  and g42665 (n23129, n_19919, n_19920);
  not g42666 (n_19921, n23129);
  and g42667 (n23130, n23118, n_19921);
  not g42668 (n_19922, n23130);
  and g42669 (n23131, n23118, n_19922);
  and g42670 (n23132, n_19921, n_19922);
  not g42671 (n_19923, n23131);
  not g42672 (n_19924, n23132);
  and g42673 (n23133, n_19923, n_19924);
  not g42674 (n_19925, n22941);
  and g42675 (n23134, n_19925, n23133);
  not g42676 (n_19926, n23133);
  and g42677 (n23135, n22941, n_19926);
  not g42678 (n_19927, n23134);
  not g42679 (n_19928, n23135);
  and g42680 (n23136, n_19927, n_19928);
  not g42681 (n_19929, n22926);
  and g42682 (n23137, n_19929, n23136);
  not g42683 (n_19930, n23136);
  and g42684 (n23138, n22926, n_19930);
  not g42685 (n_19931, n23137);
  not g42686 (n_19932, n23138);
  and g42687 (n23139, n_19931, n_19932);
  not g42688 (n_19933, n22914);
  and g42689 (n23140, n_19933, n23139);
  not g42690 (n_19934, n23140);
  and g42691 (n23141, n_19933, n_19934);
  and g42692 (n23142, n23139, n_19934);
  not g42693 (n_19935, n23141);
  not g42694 (n_19936, n23142);
  and g42695 (n23143, n_19935, n_19936);
  not g42696 (n_19937, n22913);
  not g42697 (n_19938, n23143);
  and g42698 (n23144, n_19937, n_19938);
  and g42699 (n23145, n22913, n_19936);
  and g42700 (n23146, n_19935, n23145);
  not g42701 (n_19939, n23144);
  not g42702 (n_19940, n23146);
  and g42703 (\f[92] , n_19939, n_19940);
  and g42704 (n23148, n_19934, n_19939);
  and g42705 (n23149, n_19746, n_19931);
  and g42706 (n23150, \b[57] , n5035);
  and g42707 (n23151, \b[55] , n5277);
  and g42708 (n23152, \b[56] , n5030);
  and g42714 (n23155, n5038, n11410);
  not g42717 (n_19945, n23156);
  and g42718 (n23157, \a[38] , n_19945);
  not g42719 (n_19946, n23157);
  and g42720 (n23158, \a[38] , n_19946);
  and g42721 (n23159, n_19945, n_19946);
  not g42722 (n_19947, n23158);
  not g42723 (n_19948, n23159);
  and g42724 (n23160, n_19947, n_19948);
  and g42725 (n23161, n_19894, n_19899);
  and g42726 (n23162, n_19880, n_19892);
  and g42727 (n23163, n_19855, n_19859);
  and g42728 (n23164, n_19849, n_19850);
  not g42729 (n_19949, n23164);
  and g42730 (n23165, n_19838, n_19949);
  and g42731 (n23166, \b[39] , n10426);
  and g42732 (n23167, \b[37] , n10796);
  and g42733 (n23168, \b[38] , n10421);
  and g42739 (n23171, n5451, n10429);
  not g42742 (n_19954, n23172);
  and g42743 (n23173, \a[56] , n_19954);
  not g42744 (n_19955, n23173);
  and g42745 (n23174, \a[56] , n_19955);
  and g42746 (n23175, n_19954, n_19955);
  not g42747 (n_19956, n23174);
  not g42748 (n_19957, n23175);
  and g42749 (n23176, n_19956, n_19957);
  and g42750 (n23177, n_19811, n_19812);
  not g42751 (n_19958, n23177);
  and g42752 (n23178, n_19817, n_19958);
  and g42753 (n23179, \b[29] , n13903);
  and g42754 (n23180, \b[30] , n_11555);
  not g42755 (n_19959, n23179);
  not g42756 (n_19960, n23180);
  and g42757 (n23181, n_19959, n_19960);
  not g42758 (n_19961, n23181);
  and g42759 (n23182, n_2476, n_19961);
  and g42760 (n23183, \a[29] , n23181);
  not g42761 (n_19962, n23182);
  not g42762 (n_19963, n23183);
  and g42763 (n23184, n_19962, n_19963);
  and g42764 (n23185, n_19796, n23184);
  not g42765 (n_19964, n23185);
  and g42766 (n23186, n_19796, n_19964);
  and g42767 (n23187, n23184, n_19964);
  not g42768 (n_19965, n23186);
  not g42769 (n_19966, n23187);
  and g42770 (n23188, n_19965, n_19966);
  not g42771 (n_19967, n23002);
  not g42772 (n_19968, n23188);
  and g42773 (n23189, n_19967, n_19968);
  not g42774 (n_19969, n23189);
  and g42775 (n23190, n_19967, n_19969);
  and g42776 (n23191, n_19968, n_19969);
  not g42777 (n_19970, n23190);
  not g42778 (n_19971, n23191);
  and g42779 (n23192, n_19970, n_19971);
  and g42780 (n23193, \b[33] , n12668);
  and g42781 (n23194, \b[31] , n13047);
  and g42782 (n23195, \b[32] , n12663);
  and g42788 (n23198, n4223, n12671);
  not g42791 (n_19976, n23199);
  and g42792 (n23200, \a[62] , n_19976);
  not g42793 (n_19977, n23200);
  and g42794 (n23201, \a[62] , n_19977);
  and g42795 (n23202, n_19976, n_19977);
  not g42796 (n_19978, n23201);
  not g42797 (n_19979, n23202);
  and g42798 (n23203, n_19978, n_19979);
  not g42799 (n_19980, n23192);
  and g42800 (n23204, n_19980, n23203);
  not g42801 (n_19981, n23203);
  and g42802 (n23205, n23192, n_19981);
  not g42803 (n_19982, n23204);
  not g42804 (n_19983, n23205);
  and g42805 (n23206, n_19982, n_19983);
  and g42806 (n23207, \b[36] , n11531);
  and g42807 (n23208, \b[34] , n11896);
  and g42808 (n23209, \b[35] , n11526);
  and g42814 (n23212, n4922, n11534);
  not g42817 (n_19988, n23213);
  and g42818 (n23214, \a[59] , n_19988);
  not g42819 (n_19989, n23214);
  and g42820 (n23215, \a[59] , n_19989);
  and g42821 (n23216, n_19988, n_19989);
  not g42822 (n_19990, n23215);
  not g42823 (n_19991, n23216);
  and g42824 (n23217, n_19990, n_19991);
  not g42825 (n_19992, n23206);
  not g42826 (n_19993, n23217);
  and g42827 (n23218, n_19992, n_19993);
  and g42828 (n23219, n23206, n23217);
  not g42829 (n_19994, n23218);
  not g42830 (n_19995, n23219);
  and g42831 (n23220, n_19994, n_19995);
  not g42832 (n_19996, n23178);
  and g42833 (n23221, n_19996, n23220);
  not g42834 (n_19997, n23220);
  and g42835 (n23222, n23178, n_19997);
  not g42836 (n_19998, n23221);
  not g42837 (n_19999, n23222);
  and g42838 (n23223, n_19998, n_19999);
  not g42839 (n_20000, n23176);
  and g42840 (n23224, n_20000, n23223);
  not g42841 (n_20001, n23224);
  and g42842 (n23225, n23223, n_20001);
  and g42843 (n23226, n_20000, n_20001);
  not g42844 (n_20002, n23225);
  not g42845 (n_20003, n23226);
  and g42846 (n23227, n_20002, n_20003);
  and g42847 (n23228, n_19821, n_19832);
  and g42848 (n23229, n23227, n23228);
  not g42849 (n_20004, n23227);
  not g42850 (n_20005, n23228);
  and g42851 (n23230, n_20004, n_20005);
  not g42852 (n_20006, n23229);
  not g42853 (n_20007, n23230);
  and g42854 (n23231, n_20006, n_20007);
  and g42855 (n23232, \b[42] , n9339);
  and g42856 (n23233, \b[40] , n9732);
  and g42857 (n23234, \b[41] , n9334);
  and g42863 (n23237, n6489, n9342);
  not g42866 (n_20012, n23238);
  and g42867 (n23239, \a[53] , n_20012);
  not g42868 (n_20013, n23239);
  and g42869 (n23240, \a[53] , n_20013);
  and g42870 (n23241, n_20012, n_20013);
  not g42871 (n_20014, n23240);
  not g42872 (n_20015, n23241);
  and g42873 (n23242, n_20014, n_20015);
  not g42874 (n_20016, n23242);
  and g42875 (n23243, n23231, n_20016);
  not g42876 (n_20017, n23243);
  and g42877 (n23244, n23231, n_20017);
  and g42878 (n23245, n_20016, n_20017);
  not g42879 (n_20018, n23244);
  not g42880 (n_20019, n23245);
  and g42881 (n23246, n_20018, n_20019);
  not g42882 (n_20020, n23165);
  and g42883 (n23247, n_20020, n23246);
  not g42884 (n_20021, n23246);
  and g42885 (n23248, n23165, n_20021);
  not g42886 (n_20022, n23247);
  not g42887 (n_20023, n23248);
  and g42888 (n23249, n_20022, n_20023);
  and g42889 (n23250, \b[45] , n8362);
  and g42890 (n23251, \b[43] , n8715);
  and g42891 (n23252, \b[44] , n8357);
  and g42897 (n23255, n7361, n8365);
  not g42900 (n_20028, n23256);
  and g42901 (n23257, \a[50] , n_20028);
  not g42902 (n_20029, n23257);
  and g42903 (n23258, \a[50] , n_20029);
  and g42904 (n23259, n_20028, n_20029);
  not g42905 (n_20030, n23258);
  not g42906 (n_20031, n23259);
  and g42907 (n23260, n_20030, n_20031);
  not g42908 (n_20032, n23249);
  not g42909 (n_20033, n23260);
  and g42910 (n23261, n_20032, n_20033);
  and g42911 (n23262, n23249, n23260);
  not g42912 (n_20034, n23261);
  not g42913 (n_20035, n23262);
  and g42914 (n23263, n_20034, n_20035);
  not g42915 (n_20036, n23263);
  and g42916 (n23264, n23163, n_20036);
  not g42917 (n_20037, n23163);
  and g42918 (n23265, n_20037, n23263);
  not g42919 (n_20038, n23264);
  not g42920 (n_20039, n23265);
  and g42921 (n23266, n_20038, n_20039);
  and g42922 (n23267, \b[48] , n7446);
  and g42923 (n23268, \b[46] , n7787);
  and g42924 (n23269, \b[47] , n7441);
  and g42930 (n23272, n7449, n8009);
  not g42933 (n_20044, n23273);
  and g42934 (n23274, \a[47] , n_20044);
  not g42935 (n_20045, n23274);
  and g42936 (n23275, \a[47] , n_20045);
  and g42937 (n23276, n_20044, n_20045);
  not g42938 (n_20046, n23275);
  not g42939 (n_20047, n23276);
  and g42940 (n23277, n_20046, n_20047);
  not g42941 (n_20048, n23277);
  and g42942 (n23278, n23266, n_20048);
  not g42943 (n_20049, n23278);
  and g42944 (n23279, n23266, n_20049);
  and g42945 (n23280, n_20048, n_20049);
  not g42946 (n_20050, n23279);
  not g42947 (n_20051, n23280);
  and g42948 (n23281, n_20050, n_20051);
  and g42949 (n23282, n_19863, n_19874);
  and g42950 (n23283, n23281, n23282);
  not g42951 (n_20052, n23281);
  not g42952 (n_20053, n23282);
  and g42953 (n23284, n_20052, n_20053);
  not g42954 (n_20054, n23283);
  not g42955 (n_20055, n23284);
  and g42956 (n23285, n_20054, n_20055);
  and g42957 (n23286, \b[51] , n6595);
  and g42958 (n23287, \b[49] , n6902);
  and g42959 (n23288, \b[50] , n6590);
  and g42965 (n23291, n6598, n8976);
  not g42968 (n_20060, n23292);
  and g42969 (n23293, \a[44] , n_20060);
  not g42970 (n_20061, n23293);
  and g42971 (n23294, \a[44] , n_20061);
  and g42972 (n23295, n_20060, n_20061);
  not g42973 (n_20062, n23294);
  not g42974 (n_20063, n23295);
  and g42975 (n23296, n_20062, n_20063);
  not g42976 (n_20064, n23296);
  and g42977 (n23297, n23285, n_20064);
  not g42978 (n_20065, n23285);
  and g42979 (n23298, n_20065, n23296);
  not g42980 (n_20066, n23162);
  not g42981 (n_20067, n23298);
  and g42982 (n23299, n_20066, n_20067);
  not g42983 (n_20068, n23297);
  and g42984 (n23300, n_20068, n23299);
  not g42985 (n_20069, n23300);
  and g42986 (n23301, n_20066, n_20069);
  and g42987 (n23302, n_20068, n_20069);
  and g42988 (n23303, n_20067, n23302);
  not g42989 (n_20070, n23301);
  not g42990 (n_20071, n23303);
  and g42991 (n23304, n_20070, n_20071);
  and g42992 (n23305, \b[54] , n5777);
  and g42993 (n23306, \b[52] , n6059);
  and g42994 (n23307, \b[53] , n5772);
  and g43000 (n23310, n5780, n9998);
  not g43003 (n_20076, n23311);
  and g43004 (n23312, \a[41] , n_20076);
  not g43005 (n_20077, n23312);
  and g43006 (n23313, \a[41] , n_20077);
  and g43007 (n23314, n_20076, n_20077);
  not g43008 (n_20078, n23313);
  not g43009 (n_20079, n23314);
  and g43010 (n23315, n_20078, n_20079);
  and g43011 (n23316, n23304, n23315);
  not g43012 (n_20080, n23304);
  not g43013 (n_20081, n23315);
  and g43014 (n23317, n_20080, n_20081);
  not g43015 (n_20082, n23316);
  not g43016 (n_20083, n23317);
  and g43017 (n23318, n_20082, n_20083);
  not g43018 (n_20084, n23161);
  and g43019 (n23319, n_20084, n23318);
  not g43020 (n_20085, n23318);
  and g43021 (n23320, n23161, n_20085);
  not g43022 (n_20086, n23319);
  not g43023 (n_20087, n23320);
  and g43024 (n23321, n_20086, n_20087);
  not g43025 (n_20088, n23160);
  and g43026 (n23322, n_20088, n23321);
  not g43027 (n_20089, n23322);
  and g43028 (n23323, n23321, n_20089);
  and g43029 (n23324, n_20088, n_20089);
  not g43030 (n_20090, n23323);
  not g43031 (n_20091, n23324);
  and g43032 (n23325, n_20090, n_20091);
  and g43033 (n23326, n_19903, n_19907);
  and g43034 (n23327, n23325, n23326);
  not g43035 (n_20092, n23325);
  not g43036 (n_20093, n23326);
  and g43037 (n23328, n_20092, n_20093);
  not g43038 (n_20094, n23327);
  not g43039 (n_20095, n23328);
  and g43040 (n23329, n_20094, n_20095);
  and g43041 (n23330, \b[60] , n4287);
  and g43042 (n23331, \b[58] , n4532);
  and g43043 (n23332, \b[59] , n4282);
  and g43049 (n23335, n4290, n12211);
  not g43052 (n_20100, n23336);
  and g43053 (n23337, \a[35] , n_20100);
  not g43054 (n_20101, n23337);
  and g43055 (n23338, \a[35] , n_20101);
  and g43056 (n23339, n_20100, n_20101);
  not g43057 (n_20102, n23338);
  not g43058 (n_20103, n23339);
  and g43059 (n23340, n_20102, n_20103);
  not g43060 (n_20104, n23340);
  and g43061 (n23341, n23329, n_20104);
  not g43062 (n_20105, n23341);
  and g43063 (n23342, n23329, n_20105);
  and g43064 (n23343, n_20104, n_20105);
  not g43065 (n_20106, n23342);
  not g43066 (n_20107, n23343);
  and g43067 (n23344, n_20106, n_20107);
  and g43068 (n23345, n_19911, n_19922);
  and g43069 (n23346, n23344, n23345);
  not g43070 (n_20108, n23344);
  not g43071 (n_20109, n23345);
  and g43072 (n23347, n_20108, n_20109);
  not g43073 (n_20110, n23346);
  not g43074 (n_20111, n23347);
  and g43075 (n23348, n_20110, n_20111);
  and g43076 (n23349, n_19760, n_19928);
  and g43077 (n23350, \b[63] , n3638);
  and g43078 (n23351, \b[61] , n3843);
  and g43079 (n23352, \b[62] , n3633);
  and g43085 (n23355, n3641, n13771);
  not g43088 (n_20116, n23356);
  and g43089 (n23357, \a[32] , n_20116);
  not g43090 (n_20117, n23357);
  and g43091 (n23358, \a[32] , n_20117);
  and g43092 (n23359, n_20116, n_20117);
  not g43093 (n_20118, n23358);
  not g43094 (n_20119, n23359);
  and g43095 (n23360, n_20118, n_20119);
  not g43096 (n_20120, n23349);
  not g43097 (n_20121, n23360);
  and g43098 (n23361, n_20120, n_20121);
  not g43099 (n_20122, n23361);
  and g43100 (n23362, n_20120, n_20122);
  and g43101 (n23363, n_20121, n_20122);
  not g43102 (n_20123, n23362);
  not g43103 (n_20124, n23363);
  and g43104 (n23364, n_20123, n_20124);
  not g43105 (n_20125, n23348);
  and g43106 (n23365, n_20125, n23364);
  not g43107 (n_20126, n23364);
  and g43108 (n23366, n23348, n_20126);
  not g43109 (n_20127, n23365);
  not g43110 (n_20128, n23366);
  and g43111 (n23367, n_20127, n_20128);
  not g43112 (n_20129, n23149);
  and g43113 (n23368, n_20129, n23367);
  not g43114 (n_20130, n23367);
  and g43115 (n23369, n23149, n_20130);
  not g43116 (n_20131, n23368);
  not g43117 (n_20132, n23369);
  and g43118 (n23370, n_20131, n_20132);
  not g43119 (n_20133, n23148);
  and g43120 (n23371, n_20133, n23370);
  not g43121 (n_20134, n23370);
  and g43122 (n23372, n23148, n_20134);
  not g43123 (n_20135, n23371);
  not g43124 (n_20136, n23372);
  and g43125 (\f[93] , n_20135, n_20136);
  and g43126 (n23374, n_20105, n_20111);
  and g43127 (n23375, \b[62] , n3843);
  and g43128 (n23376, \b[63] , n3633);
  not g43129 (n_20137, n23375);
  not g43130 (n_20138, n23376);
  and g43131 (n23377, n_20137, n_20138);
  and g43132 (n23378, n_12780, n23377);
  and g43133 (n23379, n13800, n23377);
  not g43134 (n_20139, n23378);
  not g43135 (n_20140, n23379);
  and g43136 (n23380, n_20139, n_20140);
  not g43137 (n_20141, n23380);
  and g43138 (n23381, \a[32] , n_20141);
  and g43139 (n23382, n_2992, n23380);
  not g43140 (n_20142, n23381);
  not g43141 (n_20143, n23382);
  and g43142 (n23383, n_20142, n_20143);
  not g43143 (n_20144, n23374);
  not g43144 (n_20145, n23383);
  and g43145 (n23384, n_20144, n_20145);
  and g43146 (n23385, n23374, n23383);
  not g43147 (n_20146, n23384);
  not g43148 (n_20147, n23385);
  and g43149 (n23386, n_20146, n_20147);
  and g43150 (n23387, \b[58] , n5035);
  and g43151 (n23388, \b[56] , n5277);
  and g43152 (n23389, \b[57] , n5030);
  and g43158 (n23392, n5038, n11436);
  not g43161 (n_20152, n23393);
  and g43162 (n23394, \a[38] , n_20152);
  not g43163 (n_20153, n23394);
  and g43164 (n23395, \a[38] , n_20153);
  and g43165 (n23396, n_20152, n_20153);
  not g43166 (n_20154, n23395);
  not g43167 (n_20155, n23396);
  and g43168 (n23397, n_20154, n_20155);
  and g43169 (n23398, n_20083, n_20086);
  and g43170 (n23399, \b[43] , n9339);
  and g43171 (n23400, \b[41] , n9732);
  and g43172 (n23401, \b[42] , n9334);
  and g43178 (n23404, n6515, n9342);
  not g43181 (n_20160, n23405);
  and g43182 (n23406, \a[53] , n_20160);
  not g43183 (n_20161, n23406);
  and g43184 (n23407, \a[53] , n_20161);
  and g43185 (n23408, n_20160, n_20161);
  not g43186 (n_20162, n23407);
  not g43187 (n_20163, n23408);
  and g43188 (n23409, n_20162, n_20163);
  and g43189 (n23410, n_20001, n_20007);
  and g43190 (n23411, \b[40] , n10426);
  and g43191 (n23412, \b[38] , n10796);
  and g43192 (n23413, \b[39] , n10421);
  and g43198 (n23416, n5955, n10429);
  not g43201 (n_20168, n23417);
  and g43202 (n23418, \a[56] , n_20168);
  not g43203 (n_20169, n23418);
  and g43204 (n23419, \a[56] , n_20169);
  and g43205 (n23420, n_20168, n_20169);
  not g43206 (n_20170, n23419);
  not g43207 (n_20171, n23420);
  and g43208 (n23421, n_20170, n_20171);
  and g43209 (n23422, n_19994, n_19998);
  and g43210 (n23423, \b[37] , n11531);
  and g43211 (n23424, \b[35] , n11896);
  and g43212 (n23425, \b[36] , n11526);
  and g43218 (n23428, n5181, n11534);
  not g43221 (n_20176, n23429);
  and g43222 (n23430, \a[59] , n_20176);
  not g43223 (n_20177, n23430);
  and g43224 (n23431, \a[59] , n_20177);
  and g43225 (n23432, n_20176, n_20177);
  not g43226 (n_20178, n23431);
  not g43227 (n_20179, n23432);
  and g43228 (n23433, n_20178, n_20179);
  and g43229 (n23434, n_19980, n_19981);
  not g43230 (n_20180, n23434);
  and g43231 (n23435, n_19969, n_20180);
  and g43232 (n23436, \b[30] , n13903);
  and g43233 (n23437, \b[31] , n_11555);
  not g43234 (n_20181, n23436);
  not g43235 (n_20182, n23437);
  and g43236 (n23438, n_20181, n_20182);
  and g43237 (n23439, n_19962, n_19964);
  not g43238 (n_20183, n23438);
  and g43239 (n23440, n_20183, n23439);
  not g43240 (n_20184, n23439);
  and g43241 (n23441, n23438, n_20184);
  not g43242 (n_20185, n23440);
  not g43243 (n_20186, n23441);
  and g43244 (n23442, n_20185, n_20186);
  and g43245 (n23443, \b[34] , n12668);
  and g43246 (n23444, \b[32] , n13047);
  and g43247 (n23445, \b[33] , n12663);
  and g43253 (n23448, n4466, n12671);
  not g43256 (n_20191, n23449);
  and g43257 (n23450, \a[62] , n_20191);
  not g43258 (n_20192, n23450);
  and g43259 (n23451, \a[62] , n_20192);
  and g43260 (n23452, n_20191, n_20192);
  not g43261 (n_20193, n23451);
  not g43262 (n_20194, n23452);
  and g43263 (n23453, n_20193, n_20194);
  not g43264 (n_20195, n23442);
  and g43265 (n23454, n_20195, n23453);
  not g43266 (n_20196, n23453);
  and g43267 (n23455, n23442, n_20196);
  not g43268 (n_20197, n23454);
  not g43269 (n_20198, n23455);
  and g43270 (n23456, n_20197, n_20198);
  not g43271 (n_20199, n23435);
  and g43272 (n23457, n_20199, n23456);
  not g43273 (n_20200, n23457);
  and g43274 (n23458, n_20199, n_20200);
  and g43275 (n23459, n23456, n_20200);
  not g43276 (n_20201, n23458);
  not g43277 (n_20202, n23459);
  and g43278 (n23460, n_20201, n_20202);
  not g43279 (n_20203, n23433);
  not g43280 (n_20204, n23460);
  and g43281 (n23461, n_20203, n_20204);
  and g43282 (n23462, n23433, n_20202);
  and g43283 (n23463, n_20201, n23462);
  not g43284 (n_20205, n23461);
  not g43285 (n_20206, n23463);
  and g43286 (n23464, n_20205, n_20206);
  not g43287 (n_20207, n23422);
  and g43288 (n23465, n_20207, n23464);
  not g43289 (n_20208, n23465);
  and g43290 (n23466, n_20207, n_20208);
  and g43291 (n23467, n23464, n_20208);
  not g43292 (n_20209, n23466);
  not g43293 (n_20210, n23467);
  and g43294 (n23468, n_20209, n_20210);
  not g43295 (n_20211, n23421);
  not g43296 (n_20212, n23468);
  and g43297 (n23469, n_20211, n_20212);
  and g43298 (n23470, n23421, n_20210);
  and g43299 (n23471, n_20209, n23470);
  not g43300 (n_20213, n23469);
  not g43301 (n_20214, n23471);
  and g43302 (n23472, n_20213, n_20214);
  not g43303 (n_20215, n23410);
  and g43304 (n23473, n_20215, n23472);
  not g43305 (n_20216, n23472);
  and g43306 (n23474, n23410, n_20216);
  not g43307 (n_20217, n23473);
  not g43308 (n_20218, n23474);
  and g43309 (n23475, n_20217, n_20218);
  not g43310 (n_20219, n23409);
  and g43311 (n23476, n_20219, n23475);
  not g43312 (n_20220, n23476);
  and g43313 (n23477, n23475, n_20220);
  and g43314 (n23478, n_20219, n_20220);
  not g43315 (n_20221, n23477);
  not g43316 (n_20222, n23478);
  and g43317 (n23479, n_20221, n_20222);
  and g43318 (n23480, n_20020, n_20021);
  not g43319 (n_20223, n23480);
  and g43320 (n23481, n_20017, n_20223);
  and g43321 (n23482, n23479, n23481);
  not g43322 (n_20224, n23479);
  not g43323 (n_20225, n23481);
  and g43324 (n23483, n_20224, n_20225);
  not g43325 (n_20226, n23482);
  not g43326 (n_20227, n23483);
  and g43327 (n23484, n_20226, n_20227);
  and g43328 (n23485, \b[46] , n8362);
  and g43329 (n23486, \b[44] , n8715);
  and g43330 (n23487, \b[45] , n8357);
  and g43336 (n23490, n7677, n8365);
  not g43339 (n_20232, n23491);
  and g43340 (n23492, \a[50] , n_20232);
  not g43341 (n_20233, n23492);
  and g43342 (n23493, \a[50] , n_20233);
  and g43343 (n23494, n_20232, n_20233);
  not g43344 (n_20234, n23493);
  not g43345 (n_20235, n23494);
  and g43346 (n23495, n_20234, n_20235);
  not g43347 (n_20236, n23495);
  and g43348 (n23496, n23484, n_20236);
  not g43349 (n_20237, n23496);
  and g43350 (n23497, n23484, n_20237);
  and g43351 (n23498, n_20236, n_20237);
  not g43352 (n_20238, n23497);
  not g43353 (n_20239, n23498);
  and g43354 (n23499, n_20238, n_20239);
  and g43355 (n23500, n_20034, n_20039);
  and g43356 (n23501, n23499, n23500);
  not g43357 (n_20240, n23499);
  not g43358 (n_20241, n23500);
  and g43359 (n23502, n_20240, n_20241);
  not g43360 (n_20242, n23501);
  not g43361 (n_20243, n23502);
  and g43362 (n23503, n_20242, n_20243);
  and g43363 (n23504, \b[49] , n7446);
  and g43364 (n23505, \b[47] , n7787);
  and g43365 (n23506, \b[48] , n7441);
  and g43371 (n23509, n7449, n8625);
  not g43374 (n_20248, n23510);
  and g43375 (n23511, \a[47] , n_20248);
  not g43376 (n_20249, n23511);
  and g43377 (n23512, \a[47] , n_20249);
  and g43378 (n23513, n_20248, n_20249);
  not g43379 (n_20250, n23512);
  not g43380 (n_20251, n23513);
  and g43381 (n23514, n_20250, n_20251);
  not g43382 (n_20252, n23514);
  and g43383 (n23515, n23503, n_20252);
  not g43384 (n_20253, n23515);
  and g43385 (n23516, n23503, n_20253);
  and g43386 (n23517, n_20252, n_20253);
  not g43387 (n_20254, n23516);
  not g43388 (n_20255, n23517);
  and g43389 (n23518, n_20254, n_20255);
  and g43390 (n23519, n_20049, n_20055);
  and g43391 (n23520, n23518, n23519);
  not g43392 (n_20256, n23518);
  not g43393 (n_20257, n23519);
  and g43394 (n23521, n_20256, n_20257);
  not g43395 (n_20258, n23520);
  not g43396 (n_20259, n23521);
  and g43397 (n23522, n_20258, n_20259);
  and g43398 (n23523, \b[52] , n6595);
  and g43399 (n23524, \b[50] , n6902);
  and g43400 (n23525, \b[51] , n6590);
  and g43406 (n23528, n6598, n9628);
  not g43409 (n_20264, n23529);
  and g43410 (n23530, \a[44] , n_20264);
  not g43411 (n_20265, n23530);
  and g43412 (n23531, \a[44] , n_20265);
  and g43413 (n23532, n_20264, n_20265);
  not g43414 (n_20266, n23531);
  not g43415 (n_20267, n23532);
  and g43416 (n23533, n_20266, n_20267);
  not g43417 (n_20268, n23533);
  and g43418 (n23534, n23522, n_20268);
  not g43419 (n_20269, n23534);
  and g43420 (n23535, n23522, n_20269);
  and g43421 (n23536, n_20268, n_20269);
  not g43422 (n_20270, n23535);
  not g43423 (n_20271, n23536);
  and g43424 (n23537, n_20270, n_20271);
  not g43425 (n_20272, n23302);
  and g43426 (n23538, n_20272, n23537);
  not g43427 (n_20273, n23537);
  and g43428 (n23539, n23302, n_20273);
  not g43429 (n_20274, n23538);
  not g43430 (n_20275, n23539);
  and g43431 (n23540, n_20274, n_20275);
  and g43432 (n23541, \b[55] , n5777);
  and g43433 (n23542, \b[53] , n6059);
  and g43434 (n23543, \b[54] , n5772);
  and g43440 (n23546, n5780, n10684);
  not g43443 (n_20280, n23547);
  and g43444 (n23548, \a[41] , n_20280);
  not g43445 (n_20281, n23548);
  and g43446 (n23549, \a[41] , n_20281);
  and g43447 (n23550, n_20280, n_20281);
  not g43448 (n_20282, n23549);
  not g43449 (n_20283, n23550);
  and g43450 (n23551, n_20282, n_20283);
  not g43451 (n_20284, n23540);
  not g43452 (n_20285, n23551);
  and g43453 (n23552, n_20284, n_20285);
  and g43454 (n23553, n23540, n23551);
  not g43455 (n_20286, n23552);
  not g43456 (n_20287, n23553);
  and g43457 (n23554, n_20286, n_20287);
  not g43458 (n_20288, n23398);
  and g43459 (n23555, n_20288, n23554);
  not g43460 (n_20289, n23554);
  and g43461 (n23556, n23398, n_20289);
  not g43462 (n_20290, n23555);
  not g43463 (n_20291, n23556);
  and g43464 (n23557, n_20290, n_20291);
  not g43465 (n_20292, n23397);
  and g43466 (n23558, n_20292, n23557);
  not g43467 (n_20293, n23558);
  and g43468 (n23559, n23557, n_20293);
  and g43469 (n23560, n_20292, n_20293);
  not g43470 (n_20294, n23559);
  not g43471 (n_20295, n23560);
  and g43472 (n23561, n_20294, n_20295);
  and g43473 (n23562, n_20089, n_20095);
  and g43474 (n23563, n23561, n23562);
  not g43475 (n_20296, n23561);
  not g43476 (n_20297, n23562);
  and g43477 (n23564, n_20296, n_20297);
  not g43478 (n_20298, n23563);
  not g43479 (n_20299, n23564);
  and g43480 (n23565, n_20298, n_20299);
  and g43481 (n23566, \b[61] , n4287);
  and g43482 (n23567, \b[59] , n4532);
  and g43483 (n23568, \b[60] , n4282);
  and g43489 (n23571, n4290, n12969);
  not g43492 (n_20304, n23572);
  and g43493 (n23573, \a[35] , n_20304);
  not g43494 (n_20305, n23573);
  and g43495 (n23574, \a[35] , n_20305);
  and g43496 (n23575, n_20304, n_20305);
  not g43497 (n_20306, n23574);
  not g43498 (n_20307, n23575);
  and g43499 (n23576, n_20306, n_20307);
  not g43500 (n_20308, n23576);
  and g43501 (n23577, n23565, n_20308);
  not g43502 (n_20309, n23565);
  and g43503 (n23578, n_20309, n23576);
  not g43504 (n_20310, n23578);
  and g43505 (n23579, n23386, n_20310);
  not g43506 (n_20311, n23577);
  and g43507 (n23580, n_20311, n23579);
  not g43508 (n_20312, n23580);
  and g43509 (n23581, n23386, n_20312);
  and g43510 (n23582, n_20310, n_20312);
  and g43511 (n23583, n_20311, n23582);
  not g43512 (n_20313, n23581);
  not g43513 (n_20314, n23583);
  and g43514 (n23584, n_20313, n_20314);
  and g43515 (n23585, n_20122, n_20128);
  not g43516 (n_20315, n23584);
  not g43517 (n_20316, n23585);
  and g43518 (n23586, n_20315, n_20316);
  not g43519 (n_20317, n23586);
  and g43520 (n23587, n_20315, n_20317);
  and g43521 (n23588, n_20316, n_20317);
  not g43522 (n_20318, n23587);
  not g43523 (n_20319, n23588);
  and g43524 (n23589, n_20318, n_20319);
  and g43525 (n23590, n_20131, n_20135);
  not g43526 (n_20320, n23589);
  not g43527 (n_20321, n23590);
  and g43528 (n23591, n_20320, n_20321);
  and g43529 (n23592, n23589, n23590);
  not g43530 (n_20322, n23591);
  not g43531 (n_20323, n23592);
  and g43532 (\f[94] , n_20322, n_20323);
  and g43533 (n23594, n_20317, n_20322);
  and g43534 (n23595, n_20146, n_20312);
  and g43535 (n23596, n_20299, n_20311);
  and g43536 (n23597, \b[63] , n3843);
  and g43537 (n23598, n3641, n13797);
  not g43538 (n_20324, n23597);
  not g43539 (n_20325, n23598);
  and g43540 (n23599, n_20324, n_20325);
  not g43541 (n_20326, n23599);
  and g43542 (n23600, \a[32] , n_20326);
  not g43543 (n_20327, n23600);
  and g43544 (n23601, \a[32] , n_20327);
  and g43545 (n23602, n_20326, n_20327);
  not g43546 (n_20328, n23601);
  not g43547 (n_20329, n23602);
  and g43548 (n23603, n_20328, n_20329);
  not g43549 (n_20330, n23596);
  not g43550 (n_20331, n23603);
  and g43551 (n23604, n_20330, n_20331);
  not g43552 (n_20332, n23604);
  and g43553 (n23605, n_20330, n_20332);
  and g43554 (n23606, n_20331, n_20332);
  not g43555 (n_20333, n23605);
  not g43556 (n_20334, n23606);
  and g43557 (n23607, n_20333, n_20334);
  and g43558 (n23608, n_20272, n_20273);
  not g43559 (n_20335, n23608);
  and g43560 (n23609, n_20286, n_20335);
  and g43561 (n23610, \b[56] , n5777);
  and g43562 (n23611, \b[54] , n6059);
  and g43563 (n23612, \b[55] , n5772);
  and g43569 (n23615, n5780, n10708);
  not g43572 (n_20340, n23616);
  and g43573 (n23617, \a[41] , n_20340);
  not g43574 (n_20341, n23617);
  and g43575 (n23618, \a[41] , n_20341);
  and g43576 (n23619, n_20340, n_20341);
  not g43577 (n_20342, n23618);
  not g43578 (n_20343, n23619);
  and g43579 (n23620, n_20342, n_20343);
  and g43580 (n23621, n_20259, n_20269);
  and g43581 (n23622, \b[53] , n6595);
  and g43582 (n23623, \b[51] , n6902);
  and g43583 (n23624, \b[52] , n6590);
  and g43589 (n23627, n6598, n9972);
  not g43592 (n_20348, n23628);
  and g43593 (n23629, \a[44] , n_20348);
  not g43594 (n_20349, n23629);
  and g43595 (n23630, \a[44] , n_20349);
  and g43596 (n23631, n_20348, n_20349);
  not g43597 (n_20350, n23630);
  not g43598 (n_20351, n23631);
  and g43599 (n23632, n_20350, n_20351);
  and g43600 (n23633, n_20243, n_20253);
  and g43601 (n23634, n_20217, n_20220);
  and g43602 (n23635, \b[44] , n9339);
  and g43603 (n23636, \b[42] , n9732);
  and g43604 (n23637, \b[43] , n9334);
  and g43610 (n23640, n7072, n9342);
  not g43613 (n_20356, n23641);
  and g43614 (n23642, \a[53] , n_20356);
  not g43615 (n_20357, n23642);
  and g43616 (n23643, \a[53] , n_20357);
  and g43617 (n23644, n_20356, n_20357);
  not g43618 (n_20358, n23643);
  not g43619 (n_20359, n23644);
  and g43620 (n23645, n_20358, n_20359);
  and g43621 (n23646, n_20208, n_20213);
  and g43622 (n23647, \b[41] , n10426);
  and g43623 (n23648, \b[39] , n10796);
  and g43624 (n23649, \b[40] , n10421);
  and g43630 (n23652, n6219, n10429);
  not g43633 (n_20364, n23653);
  and g43634 (n23654, \a[56] , n_20364);
  not g43635 (n_20365, n23654);
  and g43636 (n23655, \a[56] , n_20365);
  and g43637 (n23656, n_20364, n_20365);
  not g43638 (n_20366, n23655);
  not g43639 (n_20367, n23656);
  and g43640 (n23657, n_20366, n_20367);
  and g43641 (n23658, n_20200, n_20205);
  and g43642 (n23659, n_20186, n_20198);
  and g43643 (n23660, \b[31] , n13903);
  and g43644 (n23661, \b[32] , n_11555);
  not g43645 (n_20368, n23660);
  not g43646 (n_20369, n23661);
  and g43647 (n23662, n_20368, n_20369);
  and g43648 (n23663, n_20183, n23662);
  not g43649 (n_20370, n23662);
  and g43650 (n23664, n23438, n_20370);
  not g43651 (n_20371, n23659);
  not g43652 (n_20372, n23664);
  and g43653 (n23665, n_20371, n_20372);
  not g43654 (n_20373, n23663);
  and g43655 (n23666, n_20373, n23665);
  not g43656 (n_20374, n23666);
  and g43657 (n23667, n_20371, n_20374);
  and g43658 (n23668, n_20373, n_20374);
  and g43659 (n23669, n_20372, n23668);
  not g43660 (n_20375, n23667);
  not g43661 (n_20376, n23669);
  and g43662 (n23670, n_20375, n_20376);
  and g43663 (n23671, \b[35] , n12668);
  and g43664 (n23672, \b[33] , n13047);
  and g43665 (n23673, \b[34] , n12663);
  and g43671 (n23676, n4696, n12671);
  not g43674 (n_20381, n23677);
  and g43675 (n23678, \a[62] , n_20381);
  not g43676 (n_20382, n23678);
  and g43677 (n23679, \a[62] , n_20382);
  and g43678 (n23680, n_20381, n_20382);
  not g43679 (n_20383, n23679);
  not g43680 (n_20384, n23680);
  and g43681 (n23681, n_20383, n_20384);
  not g43682 (n_20385, n23670);
  not g43683 (n_20386, n23681);
  and g43684 (n23682, n_20385, n_20386);
  not g43685 (n_20387, n23682);
  and g43686 (n23683, n_20385, n_20387);
  and g43687 (n23684, n_20386, n_20387);
  not g43688 (n_20388, n23683);
  not g43689 (n_20389, n23684);
  and g43690 (n23685, n_20388, n_20389);
  and g43691 (n23686, \b[38] , n11531);
  and g43692 (n23687, \b[36] , n11896);
  and g43693 (n23688, \b[37] , n11526);
  and g43699 (n23691, n5205, n11534);
  not g43702 (n_20394, n23692);
  and g43703 (n23693, \a[59] , n_20394);
  not g43704 (n_20395, n23693);
  and g43705 (n23694, \a[59] , n_20395);
  and g43706 (n23695, n_20394, n_20395);
  not g43707 (n_20396, n23694);
  not g43708 (n_20397, n23695);
  and g43709 (n23696, n_20396, n_20397);
  not g43710 (n_20398, n23685);
  and g43711 (n23697, n_20398, n23696);
  not g43712 (n_20399, n23696);
  and g43713 (n23698, n23685, n_20399);
  not g43714 (n_20400, n23697);
  not g43715 (n_20401, n23698);
  and g43716 (n23699, n_20400, n_20401);
  not g43717 (n_20402, n23658);
  not g43718 (n_20403, n23699);
  and g43719 (n23700, n_20402, n_20403);
  and g43720 (n23701, n23658, n23699);
  not g43721 (n_20404, n23700);
  not g43722 (n_20405, n23701);
  and g43723 (n23702, n_20404, n_20405);
  not g43724 (n_20406, n23657);
  and g43725 (n23703, n_20406, n23702);
  not g43726 (n_20407, n23702);
  and g43727 (n23704, n23657, n_20407);
  not g43728 (n_20408, n23703);
  not g43729 (n_20409, n23704);
  and g43730 (n23705, n_20408, n_20409);
  not g43731 (n_20410, n23646);
  and g43732 (n23706, n_20410, n23705);
  not g43733 (n_20411, n23705);
  and g43734 (n23707, n23646, n_20411);
  not g43735 (n_20412, n23706);
  not g43736 (n_20413, n23707);
  and g43737 (n23708, n_20412, n_20413);
  not g43738 (n_20414, n23645);
  and g43739 (n23709, n_20414, n23708);
  not g43740 (n_20415, n23708);
  and g43741 (n23710, n23645, n_20415);
  not g43742 (n_20416, n23709);
  not g43743 (n_20417, n23710);
  and g43744 (n23711, n_20416, n_20417);
  not g43745 (n_20418, n23634);
  and g43746 (n23712, n_20418, n23711);
  not g43747 (n_20419, n23711);
  and g43748 (n23713, n23634, n_20419);
  not g43749 (n_20420, n23712);
  not g43750 (n_20421, n23713);
  and g43751 (n23714, n_20420, n_20421);
  and g43752 (n23715, \b[47] , n8362);
  and g43753 (n23716, \b[45] , n8715);
  and g43754 (n23717, \b[46] , n8357);
  and g43760 (n23720, n7703, n8365);
  not g43763 (n_20426, n23721);
  and g43764 (n23722, \a[50] , n_20426);
  not g43765 (n_20427, n23722);
  and g43766 (n23723, \a[50] , n_20427);
  and g43767 (n23724, n_20426, n_20427);
  not g43768 (n_20428, n23723);
  not g43769 (n_20429, n23724);
  and g43770 (n23725, n_20428, n_20429);
  not g43771 (n_20430, n23725);
  and g43772 (n23726, n23714, n_20430);
  not g43773 (n_20431, n23726);
  and g43774 (n23727, n23714, n_20431);
  and g43775 (n23728, n_20430, n_20431);
  not g43776 (n_20432, n23727);
  not g43777 (n_20433, n23728);
  and g43778 (n23729, n_20432, n_20433);
  and g43779 (n23730, n_20227, n_20237);
  and g43780 (n23731, n23729, n23730);
  not g43781 (n_20434, n23729);
  not g43782 (n_20435, n23730);
  and g43783 (n23732, n_20434, n_20435);
  not g43784 (n_20436, n23731);
  not g43785 (n_20437, n23732);
  and g43786 (n23733, n_20436, n_20437);
  and g43787 (n23734, \b[50] , n7446);
  and g43788 (n23735, \b[48] , n7787);
  and g43789 (n23736, \b[49] , n7441);
  and g43795 (n23739, n7449, n8949);
  not g43798 (n_20442, n23740);
  and g43799 (n23741, \a[47] , n_20442);
  not g43800 (n_20443, n23741);
  and g43801 (n23742, \a[47] , n_20443);
  and g43802 (n23743, n_20442, n_20443);
  not g43803 (n_20444, n23742);
  not g43804 (n_20445, n23743);
  and g43805 (n23744, n_20444, n_20445);
  not g43806 (n_20446, n23733);
  and g43807 (n23745, n_20446, n23744);
  not g43808 (n_20447, n23744);
  and g43809 (n23746, n23733, n_20447);
  not g43810 (n_20448, n23745);
  not g43811 (n_20449, n23746);
  and g43812 (n23747, n_20448, n_20449);
  not g43813 (n_20450, n23633);
  and g43814 (n23748, n_20450, n23747);
  not g43815 (n_20451, n23748);
  and g43816 (n23749, n_20450, n_20451);
  and g43817 (n23750, n23747, n_20451);
  not g43818 (n_20452, n23749);
  not g43819 (n_20453, n23750);
  and g43820 (n23751, n_20452, n_20453);
  not g43821 (n_20454, n23632);
  not g43822 (n_20455, n23751);
  and g43823 (n23752, n_20454, n_20455);
  and g43824 (n23753, n23632, n_20453);
  and g43825 (n23754, n_20452, n23753);
  not g43826 (n_20456, n23752);
  not g43827 (n_20457, n23754);
  and g43828 (n23755, n_20456, n_20457);
  not g43829 (n_20458, n23621);
  and g43830 (n23756, n_20458, n23755);
  not g43831 (n_20459, n23755);
  and g43832 (n23757, n23621, n_20459);
  not g43833 (n_20460, n23756);
  not g43834 (n_20461, n23757);
  and g43835 (n23758, n_20460, n_20461);
  not g43836 (n_20462, n23620);
  and g43837 (n23759, n_20462, n23758);
  not g43838 (n_20463, n23758);
  and g43839 (n23760, n23620, n_20463);
  not g43840 (n_20464, n23759);
  not g43841 (n_20465, n23760);
  and g43842 (n23761, n_20464, n_20465);
  not g43843 (n_20466, n23609);
  and g43844 (n23762, n_20466, n23761);
  not g43845 (n_20467, n23761);
  and g43846 (n23763, n23609, n_20467);
  not g43847 (n_20468, n23762);
  not g43848 (n_20469, n23763);
  and g43849 (n23764, n_20468, n_20469);
  and g43850 (n23765, \b[59] , n5035);
  and g43851 (n23766, \b[57] , n5277);
  and g43852 (n23767, \b[58] , n5030);
  and g43858 (n23770, n5038, n12179);
  not g43861 (n_20474, n23771);
  and g43862 (n23772, \a[38] , n_20474);
  not g43863 (n_20475, n23772);
  and g43864 (n23773, \a[38] , n_20475);
  and g43865 (n23774, n_20474, n_20475);
  not g43866 (n_20476, n23773);
  not g43867 (n_20477, n23774);
  and g43868 (n23775, n_20476, n_20477);
  not g43869 (n_20478, n23775);
  and g43870 (n23776, n23764, n_20478);
  not g43871 (n_20479, n23776);
  and g43872 (n23777, n23764, n_20479);
  and g43873 (n23778, n_20478, n_20479);
  not g43874 (n_20480, n23777);
  not g43875 (n_20481, n23778);
  and g43876 (n23779, n_20480, n_20481);
  and g43877 (n23780, n_20290, n_20293);
  and g43878 (n23781, n23779, n23780);
  not g43879 (n_20482, n23779);
  not g43880 (n_20483, n23780);
  and g43881 (n23782, n_20482, n_20483);
  not g43882 (n_20484, n23781);
  not g43883 (n_20485, n23782);
  and g43884 (n23783, n_20484, n_20485);
  and g43885 (n23784, \b[62] , n4287);
  and g43886 (n23785, \b[60] , n4532);
  and g43887 (n23786, \b[61] , n4282);
  and g43893 (n23789, n4290, n13370);
  not g43896 (n_20490, n23790);
  and g43897 (n23791, \a[35] , n_20490);
  not g43898 (n_20491, n23791);
  and g43899 (n23792, \a[35] , n_20491);
  and g43900 (n23793, n_20490, n_20491);
  not g43901 (n_20492, n23792);
  not g43902 (n_20493, n23793);
  and g43903 (n23794, n_20492, n_20493);
  not g43904 (n_20494, n23794);
  and g43905 (n23795, n23783, n_20494);
  not g43906 (n_20495, n23795);
  and g43907 (n23796, n23783, n_20495);
  and g43908 (n23797, n_20494, n_20495);
  not g43909 (n_20496, n23796);
  not g43910 (n_20497, n23797);
  and g43911 (n23798, n_20496, n_20497);
  not g43912 (n_20498, n23607);
  and g43913 (n23799, n_20498, n23798);
  not g43914 (n_20499, n23798);
  and g43915 (n23800, n23607, n_20499);
  not g43916 (n_20500, n23799);
  not g43917 (n_20501, n23800);
  and g43918 (n23801, n_20500, n_20501);
  not g43919 (n_20502, n23595);
  not g43920 (n_20503, n23801);
  and g43921 (n23802, n_20502, n_20503);
  not g43922 (n_20504, n23802);
  and g43923 (n23803, n_20502, n_20504);
  and g43924 (n23804, n_20503, n_20504);
  not g43925 (n_20505, n23803);
  not g43926 (n_20506, n23804);
  and g43927 (n23805, n_20505, n_20506);
  not g43928 (n_20507, n23594);
  not g43929 (n_20508, n23805);
  and g43930 (n23806, n_20507, n_20508);
  and g43931 (n23807, n23594, n_20506);
  and g43932 (n23808, n_20505, n23807);
  not g43933 (n_20509, n23806);
  not g43934 (n_20510, n23808);
  and g43935 (\f[95] , n_20509, n_20510);
  and g43936 (n23810, n_20504, n_20509);
  and g43937 (n23811, n_20498, n_20499);
  not g43938 (n_20511, n23811);
  and g43939 (n23812, n_20332, n_20511);
  and g43940 (n23813, \b[57] , n5777);
  and g43941 (n23814, \b[55] , n6059);
  and g43942 (n23815, \b[56] , n5772);
  and g43948 (n23818, n5780, n11410);
  not g43951 (n_20516, n23819);
  and g43952 (n23820, \a[41] , n_20516);
  not g43953 (n_20517, n23820);
  and g43954 (n23821, \a[41] , n_20517);
  and g43955 (n23822, n_20516, n_20517);
  not g43956 (n_20518, n23821);
  not g43957 (n_20519, n23822);
  and g43958 (n23823, n_20518, n_20519);
  and g43959 (n23824, n_20451, n_20456);
  and g43960 (n23825, n_20437, n_20449);
  and g43961 (n23826, \b[42] , n10426);
  and g43962 (n23827, \b[40] , n10796);
  and g43963 (n23828, \b[41] , n10421);
  and g43969 (n23831, n6489, n10429);
  not g43972 (n_20524, n23832);
  and g43973 (n23833, \a[56] , n_20524);
  not g43974 (n_20525, n23833);
  and g43975 (n23834, \a[56] , n_20525);
  and g43976 (n23835, n_20524, n_20525);
  not g43977 (n_20526, n23834);
  not g43978 (n_20527, n23835);
  and g43979 (n23836, n_20526, n_20527);
  and g43980 (n23837, n_20398, n_20399);
  not g43981 (n_20528, n23837);
  and g43982 (n23838, n_20387, n_20528);
  and g43983 (n23839, \b[32] , n13903);
  and g43984 (n23840, \b[33] , n_11555);
  not g43985 (n_20529, n23839);
  not g43986 (n_20530, n23840);
  and g43987 (n23841, n_20529, n_20530);
  not g43988 (n_20531, n23841);
  and g43989 (n23842, n_2992, n_20531);
  and g43990 (n23843, \a[32] , n23841);
  not g43991 (n_20532, n23842);
  not g43992 (n_20533, n23843);
  and g43993 (n23844, n_20532, n_20533);
  and g43994 (n23845, n_20370, n23844);
  not g43995 (n_20534, n23845);
  and g43996 (n23846, n_20370, n_20534);
  and g43997 (n23847, n23844, n_20534);
  not g43998 (n_20535, n23846);
  not g43999 (n_20536, n23847);
  and g44000 (n23848, n_20535, n_20536);
  not g44001 (n_20537, n23668);
  not g44002 (n_20538, n23848);
  and g44003 (n23849, n_20537, n_20538);
  not g44004 (n_20539, n23849);
  and g44005 (n23850, n_20537, n_20539);
  and g44006 (n23851, n_20538, n_20539);
  not g44007 (n_20540, n23850);
  not g44008 (n_20541, n23851);
  and g44009 (n23852, n_20540, n_20541);
  and g44010 (n23853, \b[36] , n12668);
  and g44011 (n23854, \b[34] , n13047);
  and g44012 (n23855, \b[35] , n12663);
  and g44018 (n23858, n4922, n12671);
  not g44021 (n_20546, n23859);
  and g44022 (n23860, \a[62] , n_20546);
  not g44023 (n_20547, n23860);
  and g44024 (n23861, \a[62] , n_20547);
  and g44025 (n23862, n_20546, n_20547);
  not g44026 (n_20548, n23861);
  not g44027 (n_20549, n23862);
  and g44028 (n23863, n_20548, n_20549);
  not g44029 (n_20550, n23852);
  and g44030 (n23864, n_20550, n23863);
  not g44031 (n_20551, n23863);
  and g44032 (n23865, n23852, n_20551);
  not g44033 (n_20552, n23864);
  not g44034 (n_20553, n23865);
  and g44035 (n23866, n_20552, n_20553);
  and g44036 (n23867, \b[39] , n11531);
  and g44037 (n23868, \b[37] , n11896);
  and g44038 (n23869, \b[38] , n11526);
  and g44044 (n23872, n5451, n11534);
  not g44047 (n_20558, n23873);
  and g44048 (n23874, \a[59] , n_20558);
  not g44049 (n_20559, n23874);
  and g44050 (n23875, \a[59] , n_20559);
  and g44051 (n23876, n_20558, n_20559);
  not g44052 (n_20560, n23875);
  not g44053 (n_20561, n23876);
  and g44054 (n23877, n_20560, n_20561);
  not g44055 (n_20562, n23866);
  not g44056 (n_20563, n23877);
  and g44057 (n23878, n_20562, n_20563);
  and g44058 (n23879, n23866, n23877);
  not g44059 (n_20564, n23878);
  not g44060 (n_20565, n23879);
  and g44061 (n23880, n_20564, n_20565);
  not g44062 (n_20566, n23838);
  and g44063 (n23881, n_20566, n23880);
  not g44064 (n_20567, n23880);
  and g44065 (n23882, n23838, n_20567);
  not g44066 (n_20568, n23881);
  not g44067 (n_20569, n23882);
  and g44068 (n23883, n_20568, n_20569);
  not g44069 (n_20570, n23836);
  and g44070 (n23884, n_20570, n23883);
  not g44071 (n_20571, n23884);
  and g44072 (n23885, n23883, n_20571);
  and g44073 (n23886, n_20570, n_20571);
  not g44074 (n_20572, n23885);
  not g44075 (n_20573, n23886);
  and g44076 (n23887, n_20572, n_20573);
  and g44077 (n23888, n_20404, n_20408);
  and g44078 (n23889, n23887, n23888);
  not g44079 (n_20574, n23887);
  not g44080 (n_20575, n23888);
  and g44081 (n23890, n_20574, n_20575);
  not g44082 (n_20576, n23889);
  not g44083 (n_20577, n23890);
  and g44084 (n23891, n_20576, n_20577);
  and g44085 (n23892, \b[45] , n9339);
  and g44086 (n23893, \b[43] , n9732);
  and g44087 (n23894, \b[44] , n9334);
  and g44093 (n23897, n7361, n9342);
  not g44096 (n_20582, n23898);
  and g44097 (n23899, \a[53] , n_20582);
  not g44098 (n_20583, n23899);
  and g44099 (n23900, \a[53] , n_20583);
  and g44100 (n23901, n_20582, n_20583);
  not g44101 (n_20584, n23900);
  not g44102 (n_20585, n23901);
  and g44103 (n23902, n_20584, n_20585);
  not g44104 (n_20586, n23902);
  and g44105 (n23903, n23891, n_20586);
  not g44106 (n_20587, n23903);
  and g44107 (n23904, n23891, n_20587);
  and g44108 (n23905, n_20586, n_20587);
  not g44109 (n_20588, n23904);
  not g44110 (n_20589, n23905);
  and g44111 (n23906, n_20588, n_20589);
  and g44112 (n23907, n_20412, n_20416);
  and g44113 (n23908, n23906, n23907);
  not g44114 (n_20590, n23906);
  not g44115 (n_20591, n23907);
  and g44116 (n23909, n_20590, n_20591);
  not g44117 (n_20592, n23908);
  not g44118 (n_20593, n23909);
  and g44119 (n23910, n_20592, n_20593);
  and g44120 (n23911, \b[48] , n8362);
  and g44121 (n23912, \b[46] , n8715);
  and g44122 (n23913, \b[47] , n8357);
  and g44128 (n23916, n8009, n8365);
  not g44131 (n_20598, n23917);
  and g44132 (n23918, \a[50] , n_20598);
  not g44133 (n_20599, n23918);
  and g44134 (n23919, \a[50] , n_20599);
  and g44135 (n23920, n_20598, n_20599);
  not g44136 (n_20600, n23919);
  not g44137 (n_20601, n23920);
  and g44138 (n23921, n_20600, n_20601);
  not g44139 (n_20602, n23921);
  and g44140 (n23922, n23910, n_20602);
  not g44141 (n_20603, n23922);
  and g44142 (n23923, n23910, n_20603);
  and g44143 (n23924, n_20602, n_20603);
  not g44144 (n_20604, n23923);
  not g44145 (n_20605, n23924);
  and g44146 (n23925, n_20604, n_20605);
  and g44147 (n23926, n_20420, n_20431);
  and g44148 (n23927, n23925, n23926);
  not g44149 (n_20606, n23925);
  not g44150 (n_20607, n23926);
  and g44151 (n23928, n_20606, n_20607);
  not g44152 (n_20608, n23927);
  not g44153 (n_20609, n23928);
  and g44154 (n23929, n_20608, n_20609);
  and g44155 (n23930, \b[51] , n7446);
  and g44156 (n23931, \b[49] , n7787);
  and g44157 (n23932, \b[50] , n7441);
  and g44163 (n23935, n7449, n8976);
  not g44166 (n_20614, n23936);
  and g44167 (n23937, \a[47] , n_20614);
  not g44168 (n_20615, n23937);
  and g44169 (n23938, \a[47] , n_20615);
  and g44170 (n23939, n_20614, n_20615);
  not g44171 (n_20616, n23938);
  not g44172 (n_20617, n23939);
  and g44173 (n23940, n_20616, n_20617);
  not g44174 (n_20618, n23940);
  and g44175 (n23941, n23929, n_20618);
  not g44176 (n_20619, n23929);
  and g44177 (n23942, n_20619, n23940);
  not g44178 (n_20620, n23825);
  not g44179 (n_20621, n23942);
  and g44180 (n23943, n_20620, n_20621);
  not g44181 (n_20622, n23941);
  and g44182 (n23944, n_20622, n23943);
  not g44183 (n_20623, n23944);
  and g44184 (n23945, n_20620, n_20623);
  and g44185 (n23946, n_20622, n_20623);
  and g44186 (n23947, n_20621, n23946);
  not g44187 (n_20624, n23945);
  not g44188 (n_20625, n23947);
  and g44189 (n23948, n_20624, n_20625);
  and g44190 (n23949, \b[54] , n6595);
  and g44191 (n23950, \b[52] , n6902);
  and g44192 (n23951, \b[53] , n6590);
  and g44198 (n23954, n6598, n9998);
  not g44201 (n_20630, n23955);
  and g44202 (n23956, \a[44] , n_20630);
  not g44203 (n_20631, n23956);
  and g44204 (n23957, \a[44] , n_20631);
  and g44205 (n23958, n_20630, n_20631);
  not g44206 (n_20632, n23957);
  not g44207 (n_20633, n23958);
  and g44208 (n23959, n_20632, n_20633);
  and g44209 (n23960, n23948, n23959);
  not g44210 (n_20634, n23948);
  not g44211 (n_20635, n23959);
  and g44212 (n23961, n_20634, n_20635);
  not g44213 (n_20636, n23960);
  not g44214 (n_20637, n23961);
  and g44215 (n23962, n_20636, n_20637);
  not g44216 (n_20638, n23824);
  and g44217 (n23963, n_20638, n23962);
  not g44218 (n_20639, n23962);
  and g44219 (n23964, n23824, n_20639);
  not g44220 (n_20640, n23963);
  not g44221 (n_20641, n23964);
  and g44222 (n23965, n_20640, n_20641);
  not g44223 (n_20642, n23823);
  and g44224 (n23966, n_20642, n23965);
  not g44225 (n_20643, n23966);
  and g44226 (n23967, n23965, n_20643);
  and g44227 (n23968, n_20642, n_20643);
  not g44228 (n_20644, n23967);
  not g44229 (n_20645, n23968);
  and g44230 (n23969, n_20644, n_20645);
  and g44231 (n23970, n_20460, n_20464);
  and g44232 (n23971, n23969, n23970);
  not g44233 (n_20646, n23969);
  not g44234 (n_20647, n23970);
  and g44235 (n23972, n_20646, n_20647);
  not g44236 (n_20648, n23971);
  not g44237 (n_20649, n23972);
  and g44238 (n23973, n_20648, n_20649);
  and g44239 (n23974, \b[60] , n5035);
  and g44240 (n23975, \b[58] , n5277);
  and g44241 (n23976, \b[59] , n5030);
  and g44247 (n23979, n5038, n12211);
  not g44250 (n_20654, n23980);
  and g44251 (n23981, \a[38] , n_20654);
  not g44252 (n_20655, n23981);
  and g44253 (n23982, \a[38] , n_20655);
  and g44254 (n23983, n_20654, n_20655);
  not g44255 (n_20656, n23982);
  not g44256 (n_20657, n23983);
  and g44257 (n23984, n_20656, n_20657);
  not g44258 (n_20658, n23984);
  and g44259 (n23985, n23973, n_20658);
  not g44260 (n_20659, n23985);
  and g44261 (n23986, n23973, n_20659);
  and g44262 (n23987, n_20658, n_20659);
  not g44263 (n_20660, n23986);
  not g44264 (n_20661, n23987);
  and g44265 (n23988, n_20660, n_20661);
  and g44266 (n23989, n_20468, n_20479);
  and g44267 (n23990, n23988, n23989);
  not g44268 (n_20662, n23988);
  not g44269 (n_20663, n23989);
  and g44270 (n23991, n_20662, n_20663);
  not g44271 (n_20664, n23990);
  not g44272 (n_20665, n23991);
  and g44273 (n23992, n_20664, n_20665);
  and g44274 (n23993, n_20485, n_20495);
  and g44275 (n23994, \b[63] , n4287);
  and g44276 (n23995, \b[61] , n4532);
  and g44277 (n23996, \b[62] , n4282);
  and g44283 (n23999, n4290, n13771);
  not g44286 (n_20670, n24000);
  and g44287 (n24001, \a[35] , n_20670);
  not g44288 (n_20671, n24001);
  and g44289 (n24002, \a[35] , n_20671);
  and g44290 (n24003, n_20670, n_20671);
  not g44291 (n_20672, n24002);
  not g44292 (n_20673, n24003);
  and g44293 (n24004, n_20672, n_20673);
  not g44294 (n_20674, n23993);
  not g44295 (n_20675, n24004);
  and g44296 (n24005, n_20674, n_20675);
  not g44297 (n_20676, n24005);
  and g44298 (n24006, n_20674, n_20676);
  and g44299 (n24007, n_20675, n_20676);
  not g44300 (n_20677, n24006);
  not g44301 (n_20678, n24007);
  and g44302 (n24008, n_20677, n_20678);
  not g44303 (n_20679, n23992);
  and g44304 (n24009, n_20679, n24008);
  not g44305 (n_20680, n24008);
  and g44306 (n24010, n23992, n_20680);
  not g44307 (n_20681, n24009);
  not g44308 (n_20682, n24010);
  and g44309 (n24011, n_20681, n_20682);
  not g44310 (n_20683, n23812);
  and g44311 (n24012, n_20683, n24011);
  not g44312 (n_20684, n24011);
  and g44313 (n24013, n23812, n_20684);
  not g44314 (n_20685, n24012);
  not g44315 (n_20686, n24013);
  and g44316 (n24014, n_20685, n_20686);
  not g44317 (n_20687, n23810);
  and g44318 (n24015, n_20687, n24014);
  not g44319 (n_20688, n24014);
  and g44320 (n24016, n23810, n_20688);
  not g44321 (n_20689, n24015);
  not g44322 (n_20690, n24016);
  and g44323 (\f[96] , n_20689, n_20690);
  and g44324 (n24018, n_20659, n_20665);
  and g44325 (n24019, \b[62] , n4532);
  and g44326 (n24020, \b[63] , n4282);
  not g44327 (n_20691, n24019);
  not g44328 (n_20692, n24020);
  and g44329 (n24021, n_20691, n_20692);
  not g44330 (n_20693, n4290);
  and g44331 (n24022, n_20693, n24021);
  and g44332 (n24023, n13800, n24021);
  not g44333 (n_20694, n24022);
  not g44334 (n_20695, n24023);
  and g44335 (n24024, n_20694, n_20695);
  not g44336 (n_20696, n24024);
  and g44337 (n24025, \a[35] , n_20696);
  and g44338 (n24026, n_3555, n24024);
  not g44339 (n_20697, n24025);
  not g44340 (n_20698, n24026);
  and g44341 (n24027, n_20697, n_20698);
  not g44342 (n_20699, n24018);
  not g44343 (n_20700, n24027);
  and g44344 (n24028, n_20699, n_20700);
  and g44345 (n24029, n24018, n24027);
  not g44346 (n_20701, n24028);
  not g44347 (n_20702, n24029);
  and g44348 (n24030, n_20701, n_20702);
  and g44349 (n24031, \b[58] , n5777);
  and g44350 (n24032, \b[56] , n6059);
  and g44351 (n24033, \b[57] , n5772);
  and g44357 (n24036, n5780, n11436);
  not g44360 (n_20707, n24037);
  and g44361 (n24038, \a[41] , n_20707);
  not g44362 (n_20708, n24038);
  and g44363 (n24039, \a[41] , n_20708);
  and g44364 (n24040, n_20707, n_20708);
  not g44365 (n_20709, n24039);
  not g44366 (n_20710, n24040);
  and g44367 (n24041, n_20709, n_20710);
  and g44368 (n24042, n_20637, n_20640);
  and g44369 (n24043, \b[43] , n10426);
  and g44370 (n24044, \b[41] , n10796);
  and g44371 (n24045, \b[42] , n10421);
  and g44377 (n24048, n6515, n10429);
  not g44380 (n_20715, n24049);
  and g44381 (n24050, \a[56] , n_20715);
  not g44382 (n_20716, n24050);
  and g44383 (n24051, \a[56] , n_20716);
  and g44384 (n24052, n_20715, n_20716);
  not g44385 (n_20717, n24051);
  not g44386 (n_20718, n24052);
  and g44387 (n24053, n_20717, n_20718);
  and g44388 (n24054, n_20564, n_20568);
  and g44389 (n24055, \b[40] , n11531);
  and g44390 (n24056, \b[38] , n11896);
  and g44391 (n24057, \b[39] , n11526);
  and g44397 (n24060, n5955, n11534);
  not g44400 (n_20723, n24061);
  and g44401 (n24062, \a[59] , n_20723);
  not g44402 (n_20724, n24062);
  and g44403 (n24063, \a[59] , n_20724);
  and g44404 (n24064, n_20723, n_20724);
  not g44405 (n_20725, n24063);
  not g44406 (n_20726, n24064);
  and g44407 (n24065, n_20725, n_20726);
  and g44408 (n24066, n_20550, n_20551);
  not g44409 (n_20727, n24066);
  and g44410 (n24067, n_20539, n_20727);
  and g44411 (n24068, \b[33] , n13903);
  and g44412 (n24069, \b[34] , n_11555);
  not g44413 (n_20728, n24068);
  not g44414 (n_20729, n24069);
  and g44415 (n24070, n_20728, n_20729);
  and g44416 (n24071, n_20532, n_20534);
  not g44417 (n_20730, n24070);
  and g44418 (n24072, n_20730, n24071);
  not g44419 (n_20731, n24071);
  and g44420 (n24073, n24070, n_20731);
  not g44421 (n_20732, n24072);
  not g44422 (n_20733, n24073);
  and g44423 (n24074, n_20732, n_20733);
  and g44424 (n24075, \b[37] , n12668);
  and g44425 (n24076, \b[35] , n13047);
  and g44426 (n24077, \b[36] , n12663);
  and g44432 (n24080, n5181, n12671);
  not g44435 (n_20738, n24081);
  and g44436 (n24082, \a[62] , n_20738);
  not g44437 (n_20739, n24082);
  and g44438 (n24083, \a[62] , n_20739);
  and g44439 (n24084, n_20738, n_20739);
  not g44440 (n_20740, n24083);
  not g44441 (n_20741, n24084);
  and g44442 (n24085, n_20740, n_20741);
  not g44443 (n_20742, n24074);
  and g44444 (n24086, n_20742, n24085);
  not g44445 (n_20743, n24085);
  and g44446 (n24087, n24074, n_20743);
  not g44447 (n_20744, n24086);
  not g44448 (n_20745, n24087);
  and g44449 (n24088, n_20744, n_20745);
  not g44450 (n_20746, n24067);
  and g44451 (n24089, n_20746, n24088);
  not g44452 (n_20747, n24089);
  and g44453 (n24090, n_20746, n_20747);
  and g44454 (n24091, n24088, n_20747);
  not g44455 (n_20748, n24090);
  not g44456 (n_20749, n24091);
  and g44457 (n24092, n_20748, n_20749);
  not g44458 (n_20750, n24065);
  not g44459 (n_20751, n24092);
  and g44460 (n24093, n_20750, n_20751);
  and g44461 (n24094, n24065, n_20749);
  and g44462 (n24095, n_20748, n24094);
  not g44463 (n_20752, n24093);
  not g44464 (n_20753, n24095);
  and g44465 (n24096, n_20752, n_20753);
  not g44466 (n_20754, n24054);
  and g44467 (n24097, n_20754, n24096);
  not g44468 (n_20755, n24096);
  and g44469 (n24098, n24054, n_20755);
  not g44470 (n_20756, n24097);
  not g44471 (n_20757, n24098);
  and g44472 (n24099, n_20756, n_20757);
  not g44473 (n_20758, n24053);
  and g44474 (n24100, n_20758, n24099);
  not g44475 (n_20759, n24100);
  and g44476 (n24101, n24099, n_20759);
  and g44477 (n24102, n_20758, n_20759);
  not g44478 (n_20760, n24101);
  not g44479 (n_20761, n24102);
  and g44480 (n24103, n_20760, n_20761);
  and g44481 (n24104, n_20571, n_20577);
  and g44482 (n24105, n24103, n24104);
  not g44483 (n_20762, n24103);
  not g44484 (n_20763, n24104);
  and g44485 (n24106, n_20762, n_20763);
  not g44486 (n_20764, n24105);
  not g44487 (n_20765, n24106);
  and g44488 (n24107, n_20764, n_20765);
  and g44489 (n24108, \b[46] , n9339);
  and g44490 (n24109, \b[44] , n9732);
  and g44491 (n24110, \b[45] , n9334);
  and g44497 (n24113, n7677, n9342);
  not g44500 (n_20770, n24114);
  and g44501 (n24115, \a[53] , n_20770);
  not g44502 (n_20771, n24115);
  and g44503 (n24116, \a[53] , n_20771);
  and g44504 (n24117, n_20770, n_20771);
  not g44505 (n_20772, n24116);
  not g44506 (n_20773, n24117);
  and g44507 (n24118, n_20772, n_20773);
  not g44508 (n_20774, n24118);
  and g44509 (n24119, n24107, n_20774);
  not g44510 (n_20775, n24119);
  and g44511 (n24120, n24107, n_20775);
  and g44512 (n24121, n_20774, n_20775);
  not g44513 (n_20776, n24120);
  not g44514 (n_20777, n24121);
  and g44515 (n24122, n_20776, n_20777);
  and g44516 (n24123, n_20587, n_20593);
  and g44517 (n24124, n24122, n24123);
  not g44518 (n_20778, n24122);
  not g44519 (n_20779, n24123);
  and g44520 (n24125, n_20778, n_20779);
  not g44521 (n_20780, n24124);
  not g44522 (n_20781, n24125);
  and g44523 (n24126, n_20780, n_20781);
  and g44524 (n24127, \b[49] , n8362);
  and g44525 (n24128, \b[47] , n8715);
  and g44526 (n24129, \b[48] , n8357);
  and g44532 (n24132, n8365, n8625);
  not g44535 (n_20786, n24133);
  and g44536 (n24134, \a[50] , n_20786);
  not g44537 (n_20787, n24134);
  and g44538 (n24135, \a[50] , n_20787);
  and g44539 (n24136, n_20786, n_20787);
  not g44540 (n_20788, n24135);
  not g44541 (n_20789, n24136);
  and g44542 (n24137, n_20788, n_20789);
  not g44543 (n_20790, n24137);
  and g44544 (n24138, n24126, n_20790);
  not g44545 (n_20791, n24138);
  and g44546 (n24139, n24126, n_20791);
  and g44547 (n24140, n_20790, n_20791);
  not g44548 (n_20792, n24139);
  not g44549 (n_20793, n24140);
  and g44550 (n24141, n_20792, n_20793);
  and g44551 (n24142, n_20603, n_20609);
  and g44552 (n24143, n24141, n24142);
  not g44553 (n_20794, n24141);
  not g44554 (n_20795, n24142);
  and g44555 (n24144, n_20794, n_20795);
  not g44556 (n_20796, n24143);
  not g44557 (n_20797, n24144);
  and g44558 (n24145, n_20796, n_20797);
  and g44559 (n24146, \b[52] , n7446);
  and g44560 (n24147, \b[50] , n7787);
  and g44561 (n24148, \b[51] , n7441);
  and g44567 (n24151, n7449, n9628);
  not g44570 (n_20802, n24152);
  and g44571 (n24153, \a[47] , n_20802);
  not g44572 (n_20803, n24153);
  and g44573 (n24154, \a[47] , n_20803);
  and g44574 (n24155, n_20802, n_20803);
  not g44575 (n_20804, n24154);
  not g44576 (n_20805, n24155);
  and g44577 (n24156, n_20804, n_20805);
  not g44578 (n_20806, n24156);
  and g44579 (n24157, n24145, n_20806);
  not g44580 (n_20807, n24157);
  and g44581 (n24158, n24145, n_20807);
  and g44582 (n24159, n_20806, n_20807);
  not g44583 (n_20808, n24158);
  not g44584 (n_20809, n24159);
  and g44585 (n24160, n_20808, n_20809);
  not g44586 (n_20810, n23946);
  and g44587 (n24161, n_20810, n24160);
  not g44588 (n_20811, n24160);
  and g44589 (n24162, n23946, n_20811);
  not g44590 (n_20812, n24161);
  not g44591 (n_20813, n24162);
  and g44592 (n24163, n_20812, n_20813);
  and g44593 (n24164, \b[55] , n6595);
  and g44594 (n24165, \b[53] , n6902);
  and g44595 (n24166, \b[54] , n6590);
  and g44601 (n24169, n6598, n10684);
  not g44604 (n_20818, n24170);
  and g44605 (n24171, \a[44] , n_20818);
  not g44606 (n_20819, n24171);
  and g44607 (n24172, \a[44] , n_20819);
  and g44608 (n24173, n_20818, n_20819);
  not g44609 (n_20820, n24172);
  not g44610 (n_20821, n24173);
  and g44611 (n24174, n_20820, n_20821);
  not g44612 (n_20822, n24163);
  not g44613 (n_20823, n24174);
  and g44614 (n24175, n_20822, n_20823);
  and g44615 (n24176, n24163, n24174);
  not g44616 (n_20824, n24175);
  not g44617 (n_20825, n24176);
  and g44618 (n24177, n_20824, n_20825);
  not g44619 (n_20826, n24042);
  and g44620 (n24178, n_20826, n24177);
  not g44621 (n_20827, n24177);
  and g44622 (n24179, n24042, n_20827);
  not g44623 (n_20828, n24178);
  not g44624 (n_20829, n24179);
  and g44625 (n24180, n_20828, n_20829);
  not g44626 (n_20830, n24041);
  and g44627 (n24181, n_20830, n24180);
  not g44628 (n_20831, n24181);
  and g44629 (n24182, n24180, n_20831);
  and g44630 (n24183, n_20830, n_20831);
  not g44631 (n_20832, n24182);
  not g44632 (n_20833, n24183);
  and g44633 (n24184, n_20832, n_20833);
  and g44634 (n24185, n_20643, n_20649);
  and g44635 (n24186, n24184, n24185);
  not g44636 (n_20834, n24184);
  not g44637 (n_20835, n24185);
  and g44638 (n24187, n_20834, n_20835);
  not g44639 (n_20836, n24186);
  not g44640 (n_20837, n24187);
  and g44641 (n24188, n_20836, n_20837);
  and g44642 (n24189, \b[61] , n5035);
  and g44643 (n24190, \b[59] , n5277);
  and g44644 (n24191, \b[60] , n5030);
  and g44650 (n24194, n5038, n12969);
  not g44653 (n_20842, n24195);
  and g44654 (n24196, \a[38] , n_20842);
  not g44655 (n_20843, n24196);
  and g44656 (n24197, \a[38] , n_20843);
  and g44657 (n24198, n_20842, n_20843);
  not g44658 (n_20844, n24197);
  not g44659 (n_20845, n24198);
  and g44660 (n24199, n_20844, n_20845);
  not g44661 (n_20846, n24199);
  and g44662 (n24200, n24188, n_20846);
  not g44663 (n_20847, n24188);
  and g44664 (n24201, n_20847, n24199);
  not g44665 (n_20848, n24201);
  and g44666 (n24202, n24030, n_20848);
  not g44667 (n_20849, n24200);
  and g44668 (n24203, n_20849, n24202);
  not g44669 (n_20850, n24203);
  and g44670 (n24204, n24030, n_20850);
  and g44671 (n24205, n_20848, n_20850);
  and g44672 (n24206, n_20849, n24205);
  not g44673 (n_20851, n24204);
  not g44674 (n_20852, n24206);
  and g44675 (n24207, n_20851, n_20852);
  and g44676 (n24208, n_20676, n_20682);
  not g44677 (n_20853, n24207);
  not g44678 (n_20854, n24208);
  and g44679 (n24209, n_20853, n_20854);
  not g44680 (n_20855, n24209);
  and g44681 (n24210, n_20853, n_20855);
  and g44682 (n24211, n_20854, n_20855);
  not g44683 (n_20856, n24210);
  not g44684 (n_20857, n24211);
  and g44685 (n24212, n_20856, n_20857);
  and g44686 (n24213, n_20685, n_20689);
  not g44687 (n_20858, n24212);
  not g44688 (n_20859, n24213);
  and g44689 (n24214, n_20858, n_20859);
  and g44690 (n24215, n24212, n24213);
  not g44691 (n_20860, n24214);
  not g44692 (n_20861, n24215);
  and g44693 (\f[97] , n_20860, n_20861);
  and g44694 (n24217, n_20855, n_20860);
  and g44695 (n24218, n_20701, n_20850);
  and g44696 (n24219, n_20837, n_20849);
  and g44697 (n24220, \b[63] , n4532);
  and g44698 (n24221, n4290, n13797);
  not g44699 (n_20862, n24220);
  not g44700 (n_20863, n24221);
  and g44701 (n24222, n_20862, n_20863);
  not g44702 (n_20864, n24222);
  and g44703 (n24223, \a[35] , n_20864);
  not g44704 (n_20865, n24223);
  and g44705 (n24224, \a[35] , n_20865);
  and g44706 (n24225, n_20864, n_20865);
  not g44707 (n_20866, n24224);
  not g44708 (n_20867, n24225);
  and g44709 (n24226, n_20866, n_20867);
  not g44710 (n_20868, n24219);
  not g44711 (n_20869, n24226);
  and g44712 (n24227, n_20868, n_20869);
  not g44713 (n_20870, n24227);
  and g44714 (n24228, n_20868, n_20870);
  and g44715 (n24229, n_20869, n_20870);
  not g44716 (n_20871, n24228);
  not g44717 (n_20872, n24229);
  and g44718 (n24230, n_20871, n_20872);
  and g44719 (n24231, n_20810, n_20811);
  not g44720 (n_20873, n24231);
  and g44721 (n24232, n_20824, n_20873);
  and g44722 (n24233, \b[56] , n6595);
  and g44723 (n24234, \b[54] , n6902);
  and g44724 (n24235, \b[55] , n6590);
  and g44730 (n24238, n6598, n10708);
  not g44733 (n_20878, n24239);
  and g44734 (n24240, \a[44] , n_20878);
  not g44735 (n_20879, n24240);
  and g44736 (n24241, \a[44] , n_20879);
  and g44737 (n24242, n_20878, n_20879);
  not g44738 (n_20880, n24241);
  not g44739 (n_20881, n24242);
  and g44740 (n24243, n_20880, n_20881);
  and g44741 (n24244, n_20797, n_20807);
  and g44742 (n24245, \b[53] , n7446);
  and g44743 (n24246, \b[51] , n7787);
  and g44744 (n24247, \b[52] , n7441);
  and g44750 (n24250, n7449, n9972);
  not g44753 (n_20886, n24251);
  and g44754 (n24252, \a[47] , n_20886);
  not g44755 (n_20887, n24252);
  and g44756 (n24253, \a[47] , n_20887);
  and g44757 (n24254, n_20886, n_20887);
  not g44758 (n_20888, n24253);
  not g44759 (n_20889, n24254);
  and g44760 (n24255, n_20888, n_20889);
  and g44761 (n24256, n_20781, n_20791);
  and g44762 (n24257, n_20756, n_20759);
  and g44763 (n24258, \b[44] , n10426);
  and g44764 (n24259, \b[42] , n10796);
  and g44765 (n24260, \b[43] , n10421);
  and g44771 (n24263, n7072, n10429);
  not g44774 (n_20894, n24264);
  and g44775 (n24265, \a[56] , n_20894);
  not g44776 (n_20895, n24265);
  and g44777 (n24266, \a[56] , n_20895);
  and g44778 (n24267, n_20894, n_20895);
  not g44779 (n_20896, n24266);
  not g44780 (n_20897, n24267);
  and g44781 (n24268, n_20896, n_20897);
  and g44782 (n24269, n_20747, n_20752);
  and g44783 (n24270, n_20733, n_20745);
  and g44784 (n24271, \b[34] , n13903);
  and g44785 (n24272, \b[35] , n_11555);
  not g44786 (n_20898, n24271);
  not g44787 (n_20899, n24272);
  and g44788 (n24273, n_20898, n_20899);
  and g44789 (n24274, n_20730, n24273);
  not g44790 (n_20900, n24273);
  and g44791 (n24275, n24070, n_20900);
  not g44792 (n_20901, n24270);
  not g44793 (n_20902, n24275);
  and g44794 (n24276, n_20901, n_20902);
  not g44795 (n_20903, n24274);
  and g44796 (n24277, n_20903, n24276);
  not g44797 (n_20904, n24277);
  and g44798 (n24278, n_20901, n_20904);
  and g44799 (n24279, n_20903, n_20904);
  and g44800 (n24280, n_20902, n24279);
  not g44801 (n_20905, n24278);
  not g44802 (n_20906, n24280);
  and g44803 (n24281, n_20905, n_20906);
  and g44804 (n24282, \b[38] , n12668);
  and g44805 (n24283, \b[36] , n13047);
  and g44806 (n24284, \b[37] , n12663);
  and g44812 (n24287, n5205, n12671);
  not g44815 (n_20911, n24288);
  and g44816 (n24289, \a[62] , n_20911);
  not g44817 (n_20912, n24289);
  and g44818 (n24290, \a[62] , n_20912);
  and g44819 (n24291, n_20911, n_20912);
  not g44820 (n_20913, n24290);
  not g44821 (n_20914, n24291);
  and g44822 (n24292, n_20913, n_20914);
  not g44823 (n_20915, n24281);
  not g44824 (n_20916, n24292);
  and g44825 (n24293, n_20915, n_20916);
  not g44826 (n_20917, n24293);
  and g44827 (n24294, n_20915, n_20917);
  and g44828 (n24295, n_20916, n_20917);
  not g44829 (n_20918, n24294);
  not g44830 (n_20919, n24295);
  and g44831 (n24296, n_20918, n_20919);
  and g44832 (n24297, \b[41] , n11531);
  and g44833 (n24298, \b[39] , n11896);
  and g44834 (n24299, \b[40] , n11526);
  and g44840 (n24302, n6219, n11534);
  not g44843 (n_20924, n24303);
  and g44844 (n24304, \a[59] , n_20924);
  not g44845 (n_20925, n24304);
  and g44846 (n24305, \a[59] , n_20925);
  and g44847 (n24306, n_20924, n_20925);
  not g44848 (n_20926, n24305);
  not g44849 (n_20927, n24306);
  and g44850 (n24307, n_20926, n_20927);
  not g44851 (n_20928, n24296);
  and g44852 (n24308, n_20928, n24307);
  not g44853 (n_20929, n24307);
  and g44854 (n24309, n24296, n_20929);
  not g44855 (n_20930, n24308);
  not g44856 (n_20931, n24309);
  and g44857 (n24310, n_20930, n_20931);
  not g44858 (n_20932, n24269);
  not g44859 (n_20933, n24310);
  and g44860 (n24311, n_20932, n_20933);
  and g44861 (n24312, n24269, n24310);
  not g44862 (n_20934, n24311);
  not g44863 (n_20935, n24312);
  and g44864 (n24313, n_20934, n_20935);
  not g44865 (n_20936, n24268);
  and g44866 (n24314, n_20936, n24313);
  not g44867 (n_20937, n24313);
  and g44868 (n24315, n24268, n_20937);
  not g44869 (n_20938, n24314);
  not g44870 (n_20939, n24315);
  and g44871 (n24316, n_20938, n_20939);
  not g44872 (n_20940, n24257);
  and g44873 (n24317, n_20940, n24316);
  not g44874 (n_20941, n24316);
  and g44875 (n24318, n24257, n_20941);
  not g44876 (n_20942, n24317);
  not g44877 (n_20943, n24318);
  and g44878 (n24319, n_20942, n_20943);
  and g44879 (n24320, \b[47] , n9339);
  and g44880 (n24321, \b[45] , n9732);
  and g44881 (n24322, \b[46] , n9334);
  and g44887 (n24325, n7703, n9342);
  not g44890 (n_20948, n24326);
  and g44891 (n24327, \a[53] , n_20948);
  not g44892 (n_20949, n24327);
  and g44893 (n24328, \a[53] , n_20949);
  and g44894 (n24329, n_20948, n_20949);
  not g44895 (n_20950, n24328);
  not g44896 (n_20951, n24329);
  and g44897 (n24330, n_20950, n_20951);
  not g44898 (n_20952, n24330);
  and g44899 (n24331, n24319, n_20952);
  not g44900 (n_20953, n24331);
  and g44901 (n24332, n24319, n_20953);
  and g44902 (n24333, n_20952, n_20953);
  not g44903 (n_20954, n24332);
  not g44904 (n_20955, n24333);
  and g44905 (n24334, n_20954, n_20955);
  and g44906 (n24335, n_20765, n_20775);
  and g44907 (n24336, n24334, n24335);
  not g44908 (n_20956, n24334);
  not g44909 (n_20957, n24335);
  and g44910 (n24337, n_20956, n_20957);
  not g44911 (n_20958, n24336);
  not g44912 (n_20959, n24337);
  and g44913 (n24338, n_20958, n_20959);
  and g44914 (n24339, \b[50] , n8362);
  and g44915 (n24340, \b[48] , n8715);
  and g44916 (n24341, \b[49] , n8357);
  and g44922 (n24344, n8365, n8949);
  not g44925 (n_20964, n24345);
  and g44926 (n24346, \a[50] , n_20964);
  not g44927 (n_20965, n24346);
  and g44928 (n24347, \a[50] , n_20965);
  and g44929 (n24348, n_20964, n_20965);
  not g44930 (n_20966, n24347);
  not g44931 (n_20967, n24348);
  and g44932 (n24349, n_20966, n_20967);
  not g44933 (n_20968, n24338);
  and g44934 (n24350, n_20968, n24349);
  not g44935 (n_20969, n24349);
  and g44936 (n24351, n24338, n_20969);
  not g44937 (n_20970, n24350);
  not g44938 (n_20971, n24351);
  and g44939 (n24352, n_20970, n_20971);
  not g44940 (n_20972, n24256);
  and g44941 (n24353, n_20972, n24352);
  not g44942 (n_20973, n24353);
  and g44943 (n24354, n_20972, n_20973);
  and g44944 (n24355, n24352, n_20973);
  not g44945 (n_20974, n24354);
  not g44946 (n_20975, n24355);
  and g44947 (n24356, n_20974, n_20975);
  not g44948 (n_20976, n24255);
  not g44949 (n_20977, n24356);
  and g44950 (n24357, n_20976, n_20977);
  and g44951 (n24358, n24255, n_20975);
  and g44952 (n24359, n_20974, n24358);
  not g44953 (n_20978, n24357);
  not g44954 (n_20979, n24359);
  and g44955 (n24360, n_20978, n_20979);
  not g44956 (n_20980, n24244);
  and g44957 (n24361, n_20980, n24360);
  not g44958 (n_20981, n24360);
  and g44959 (n24362, n24244, n_20981);
  not g44960 (n_20982, n24361);
  not g44961 (n_20983, n24362);
  and g44962 (n24363, n_20982, n_20983);
  not g44963 (n_20984, n24243);
  and g44964 (n24364, n_20984, n24363);
  not g44965 (n_20985, n24363);
  and g44966 (n24365, n24243, n_20985);
  not g44967 (n_20986, n24364);
  not g44968 (n_20987, n24365);
  and g44969 (n24366, n_20986, n_20987);
  not g44970 (n_20988, n24232);
  and g44971 (n24367, n_20988, n24366);
  not g44972 (n_20989, n24366);
  and g44973 (n24368, n24232, n_20989);
  not g44974 (n_20990, n24367);
  not g44975 (n_20991, n24368);
  and g44976 (n24369, n_20990, n_20991);
  and g44977 (n24370, \b[59] , n5777);
  and g44978 (n24371, \b[57] , n6059);
  and g44979 (n24372, \b[58] , n5772);
  and g44985 (n24375, n5780, n12179);
  not g44988 (n_20996, n24376);
  and g44989 (n24377, \a[41] , n_20996);
  not g44990 (n_20997, n24377);
  and g44991 (n24378, \a[41] , n_20997);
  and g44992 (n24379, n_20996, n_20997);
  not g44993 (n_20998, n24378);
  not g44994 (n_20999, n24379);
  and g44995 (n24380, n_20998, n_20999);
  not g44996 (n_21000, n24380);
  and g44997 (n24381, n24369, n_21000);
  not g44998 (n_21001, n24381);
  and g44999 (n24382, n24369, n_21001);
  and g45000 (n24383, n_21000, n_21001);
  not g45001 (n_21002, n24382);
  not g45002 (n_21003, n24383);
  and g45003 (n24384, n_21002, n_21003);
  and g45004 (n24385, n_20828, n_20831);
  and g45005 (n24386, n24384, n24385);
  not g45006 (n_21004, n24384);
  not g45007 (n_21005, n24385);
  and g45008 (n24387, n_21004, n_21005);
  not g45009 (n_21006, n24386);
  not g45010 (n_21007, n24387);
  and g45011 (n24388, n_21006, n_21007);
  and g45012 (n24389, \b[62] , n5035);
  and g45013 (n24390, \b[60] , n5277);
  and g45014 (n24391, \b[61] , n5030);
  and g45020 (n24394, n5038, n13370);
  not g45023 (n_21012, n24395);
  and g45024 (n24396, \a[38] , n_21012);
  not g45025 (n_21013, n24396);
  and g45026 (n24397, \a[38] , n_21013);
  and g45027 (n24398, n_21012, n_21013);
  not g45028 (n_21014, n24397);
  not g45029 (n_21015, n24398);
  and g45030 (n24399, n_21014, n_21015);
  not g45031 (n_21016, n24399);
  and g45032 (n24400, n24388, n_21016);
  not g45033 (n_21017, n24400);
  and g45034 (n24401, n24388, n_21017);
  and g45035 (n24402, n_21016, n_21017);
  not g45036 (n_21018, n24401);
  not g45037 (n_21019, n24402);
  and g45038 (n24403, n_21018, n_21019);
  not g45039 (n_21020, n24230);
  and g45040 (n24404, n_21020, n24403);
  not g45041 (n_21021, n24403);
  and g45042 (n24405, n24230, n_21021);
  not g45043 (n_21022, n24404);
  not g45044 (n_21023, n24405);
  and g45045 (n24406, n_21022, n_21023);
  not g45046 (n_21024, n24218);
  not g45047 (n_21025, n24406);
  and g45048 (n24407, n_21024, n_21025);
  and g45049 (n24408, n24218, n24406);
  not g45050 (n_21026, n24407);
  not g45051 (n_21027, n24408);
  and g45052 (n24409, n_21026, n_21027);
  not g45053 (n_21028, n24217);
  and g45054 (n24410, n_21028, n24409);
  not g45055 (n_21029, n24409);
  and g45056 (n24411, n24217, n_21029);
  not g45057 (n_21030, n24410);
  not g45058 (n_21031, n24411);
  and g45059 (\f[98] , n_21030, n_21031);
  and g45060 (n24413, n_21026, n_21030);
  and g45061 (n24414, n_20973, n_20978);
  and g45062 (n24415, \b[54] , n7446);
  and g45063 (n24416, \b[52] , n7787);
  and g45064 (n24417, \b[53] , n7441);
  and g45070 (n24420, n7449, n9998);
  not g45073 (n_21036, n24421);
  and g45074 (n24422, \a[47] , n_21036);
  not g45075 (n_21037, n24422);
  and g45076 (n24423, \a[47] , n_21037);
  and g45077 (n24424, n_21036, n_21037);
  not g45078 (n_21038, n24423);
  not g45079 (n_21039, n24424);
  and g45080 (n24425, n_21038, n_21039);
  and g45081 (n24426, n_20959, n_20971);
  and g45082 (n24427, \b[35] , n13903);
  and g45083 (n24428, \b[36] , n_11555);
  not g45084 (n_21040, n24427);
  not g45085 (n_21041, n24428);
  and g45086 (n24429, n_21040, n_21041);
  and g45087 (n24430, \a[35] , n_20900);
  and g45088 (n24431, n_3555, n24273);
  not g45089 (n_21042, n24430);
  not g45090 (n_21043, n24431);
  and g45091 (n24432, n_21042, n_21043);
  not g45092 (n_21044, n24429);
  not g45093 (n_21045, n24432);
  and g45094 (n24433, n_21044, n_21045);
  and g45095 (n24434, n24429, n24432);
  not g45096 (n_21046, n24433);
  not g45097 (n_21047, n24434);
  and g45098 (n24435, n_21046, n_21047);
  not g45099 (n_21048, n24279);
  and g45100 (n24436, n_21048, n24435);
  not g45101 (n_21049, n24435);
  and g45102 (n24437, n24279, n_21049);
  not g45103 (n_21050, n24436);
  not g45104 (n_21051, n24437);
  and g45105 (n24438, n_21050, n_21051);
  and g45106 (n24439, \b[39] , n12668);
  and g45107 (n24440, \b[37] , n13047);
  and g45108 (n24441, \b[38] , n12663);
  and g45114 (n24444, n5451, n12671);
  not g45117 (n_21056, n24445);
  and g45118 (n24446, \a[62] , n_21056);
  not g45119 (n_21057, n24446);
  and g45120 (n24447, \a[62] , n_21057);
  and g45121 (n24448, n_21056, n_21057);
  not g45122 (n_21058, n24447);
  not g45123 (n_21059, n24448);
  and g45124 (n24449, n_21058, n_21059);
  not g45125 (n_21060, n24438);
  and g45126 (n24450, n_21060, n24449);
  not g45127 (n_21061, n24449);
  and g45128 (n24451, n24438, n_21061);
  not g45129 (n_21062, n24450);
  not g45130 (n_21063, n24451);
  and g45131 (n24452, n_21062, n_21063);
  and g45132 (n24453, \b[42] , n11531);
  and g45133 (n24454, \b[40] , n11896);
  and g45134 (n24455, \b[41] , n11526);
  and g45140 (n24458, n6489, n11534);
  not g45143 (n_21068, n24459);
  and g45144 (n24460, \a[59] , n_21068);
  not g45145 (n_21069, n24460);
  and g45146 (n24461, \a[59] , n_21069);
  and g45147 (n24462, n_21068, n_21069);
  not g45148 (n_21070, n24461);
  not g45149 (n_21071, n24462);
  and g45150 (n24463, n_21070, n_21071);
  not g45151 (n_21072, n24463);
  and g45152 (n24464, n24452, n_21072);
  not g45153 (n_21073, n24464);
  and g45154 (n24465, n24452, n_21073);
  and g45155 (n24466, n_21072, n_21073);
  not g45156 (n_21074, n24465);
  not g45157 (n_21075, n24466);
  and g45158 (n24467, n_21074, n_21075);
  and g45159 (n24468, n_20928, n_20929);
  not g45160 (n_21076, n24468);
  and g45161 (n24469, n_20917, n_21076);
  not g45162 (n_21077, n24467);
  not g45163 (n_21078, n24469);
  and g45164 (n24470, n_21077, n_21078);
  not g45165 (n_21079, n24470);
  and g45166 (n24471, n_21077, n_21079);
  and g45167 (n24472, n_21078, n_21079);
  not g45168 (n_21080, n24471);
  not g45169 (n_21081, n24472);
  and g45170 (n24473, n_21080, n_21081);
  and g45171 (n24474, \b[45] , n10426);
  and g45172 (n24475, \b[43] , n10796);
  and g45173 (n24476, \b[44] , n10421);
  and g45179 (n24479, n7361, n10429);
  not g45182 (n_21086, n24480);
  and g45183 (n24481, \a[56] , n_21086);
  not g45184 (n_21087, n24481);
  and g45185 (n24482, \a[56] , n_21087);
  and g45186 (n24483, n_21086, n_21087);
  not g45187 (n_21088, n24482);
  not g45188 (n_21089, n24483);
  and g45189 (n24484, n_21088, n_21089);
  not g45190 (n_21090, n24473);
  not g45191 (n_21091, n24484);
  and g45192 (n24485, n_21090, n_21091);
  not g45193 (n_21092, n24485);
  and g45194 (n24486, n_21090, n_21092);
  and g45195 (n24487, n_21091, n_21092);
  not g45196 (n_21093, n24486);
  not g45197 (n_21094, n24487);
  and g45198 (n24488, n_21093, n_21094);
  and g45199 (n24489, n_20934, n_20938);
  and g45200 (n24490, n24488, n24489);
  not g45201 (n_21095, n24488);
  not g45202 (n_21096, n24489);
  and g45203 (n24491, n_21095, n_21096);
  not g45204 (n_21097, n24490);
  not g45205 (n_21098, n24491);
  and g45206 (n24492, n_21097, n_21098);
  and g45207 (n24493, \b[48] , n9339);
  and g45208 (n24494, \b[46] , n9732);
  and g45209 (n24495, \b[47] , n9334);
  and g45215 (n24498, n8009, n9342);
  not g45218 (n_21103, n24499);
  and g45219 (n24500, \a[53] , n_21103);
  not g45220 (n_21104, n24500);
  and g45221 (n24501, \a[53] , n_21104);
  and g45222 (n24502, n_21103, n_21104);
  not g45223 (n_21105, n24501);
  not g45224 (n_21106, n24502);
  and g45225 (n24503, n_21105, n_21106);
  not g45226 (n_21107, n24503);
  and g45227 (n24504, n24492, n_21107);
  not g45228 (n_21108, n24504);
  and g45229 (n24505, n24492, n_21108);
  and g45230 (n24506, n_21107, n_21108);
  not g45231 (n_21109, n24505);
  not g45232 (n_21110, n24506);
  and g45233 (n24507, n_21109, n_21110);
  and g45234 (n24508, n_20942, n_20953);
  and g45235 (n24509, n24507, n24508);
  not g45236 (n_21111, n24507);
  not g45237 (n_21112, n24508);
  and g45238 (n24510, n_21111, n_21112);
  not g45239 (n_21113, n24509);
  not g45240 (n_21114, n24510);
  and g45241 (n24511, n_21113, n_21114);
  and g45242 (n24512, \b[51] , n8362);
  and g45243 (n24513, \b[49] , n8715);
  and g45244 (n24514, \b[50] , n8357);
  and g45250 (n24517, n8365, n8976);
  not g45253 (n_21119, n24518);
  and g45254 (n24519, \a[50] , n_21119);
  not g45255 (n_21120, n24519);
  and g45256 (n24520, \a[50] , n_21120);
  and g45257 (n24521, n_21119, n_21120);
  not g45258 (n_21121, n24520);
  not g45259 (n_21122, n24521);
  and g45260 (n24522, n_21121, n_21122);
  not g45261 (n_21123, n24511);
  and g45262 (n24523, n_21123, n24522);
  not g45263 (n_21124, n24522);
  and g45264 (n24524, n24511, n_21124);
  not g45265 (n_21125, n24523);
  not g45266 (n_21126, n24524);
  and g45267 (n24525, n_21125, n_21126);
  not g45268 (n_21127, n24426);
  and g45269 (n24526, n_21127, n24525);
  not g45270 (n_21128, n24525);
  and g45271 (n24527, n24426, n_21128);
  not g45272 (n_21129, n24526);
  not g45273 (n_21130, n24527);
  and g45274 (n24528, n_21129, n_21130);
  not g45275 (n_21131, n24425);
  and g45276 (n24529, n_21131, n24528);
  not g45277 (n_21132, n24528);
  and g45278 (n24530, n24425, n_21132);
  not g45279 (n_21133, n24529);
  not g45280 (n_21134, n24530);
  and g45281 (n24531, n_21133, n_21134);
  not g45282 (n_21135, n24414);
  and g45283 (n24532, n_21135, n24531);
  not g45284 (n_21136, n24531);
  and g45285 (n24533, n24414, n_21136);
  not g45286 (n_21137, n24532);
  not g45287 (n_21138, n24533);
  and g45288 (n24534, n_21137, n_21138);
  and g45289 (n24535, \b[57] , n6595);
  and g45290 (n24536, \b[55] , n6902);
  and g45291 (n24537, \b[56] , n6590);
  and g45297 (n24540, n6598, n11410);
  not g45300 (n_21143, n24541);
  and g45301 (n24542, \a[44] , n_21143);
  not g45302 (n_21144, n24542);
  and g45303 (n24543, \a[44] , n_21144);
  and g45304 (n24544, n_21143, n_21144);
  not g45305 (n_21145, n24543);
  not g45306 (n_21146, n24544);
  and g45307 (n24545, n_21145, n_21146);
  not g45308 (n_21147, n24545);
  and g45309 (n24546, n24534, n_21147);
  not g45310 (n_21148, n24546);
  and g45311 (n24547, n24534, n_21148);
  and g45312 (n24548, n_21147, n_21148);
  not g45313 (n_21149, n24547);
  not g45314 (n_21150, n24548);
  and g45315 (n24549, n_21149, n_21150);
  and g45316 (n24550, n_20982, n_20986);
  and g45317 (n24551, n24549, n24550);
  not g45318 (n_21151, n24549);
  not g45319 (n_21152, n24550);
  and g45320 (n24552, n_21151, n_21152);
  not g45321 (n_21153, n24551);
  not g45322 (n_21154, n24552);
  and g45323 (n24553, n_21153, n_21154);
  and g45324 (n24554, \b[60] , n5777);
  and g45325 (n24555, \b[58] , n6059);
  and g45326 (n24556, \b[59] , n5772);
  and g45332 (n24559, n5780, n12211);
  not g45335 (n_21159, n24560);
  and g45336 (n24561, \a[41] , n_21159);
  not g45337 (n_21160, n24561);
  and g45338 (n24562, \a[41] , n_21160);
  and g45339 (n24563, n_21159, n_21160);
  not g45340 (n_21161, n24562);
  not g45341 (n_21162, n24563);
  and g45342 (n24564, n_21161, n_21162);
  not g45343 (n_21163, n24564);
  and g45344 (n24565, n24553, n_21163);
  not g45345 (n_21164, n24565);
  and g45346 (n24566, n24553, n_21164);
  and g45347 (n24567, n_21163, n_21164);
  not g45348 (n_21165, n24566);
  not g45349 (n_21166, n24567);
  and g45350 (n24568, n_21165, n_21166);
  and g45351 (n24569, n_20990, n_21001);
  and g45352 (n24570, n24568, n24569);
  not g45353 (n_21167, n24568);
  not g45354 (n_21168, n24569);
  and g45355 (n24571, n_21167, n_21168);
  not g45356 (n_21169, n24570);
  not g45357 (n_21170, n24571);
  and g45358 (n24572, n_21169, n_21170);
  and g45359 (n24573, \b[63] , n5035);
  and g45360 (n24574, \b[61] , n5277);
  and g45361 (n24575, \b[62] , n5030);
  and g45367 (n24578, n5038, n13771);
  not g45370 (n_21175, n24579);
  and g45371 (n24580, \a[38] , n_21175);
  not g45372 (n_21176, n24580);
  and g45373 (n24581, \a[38] , n_21176);
  and g45374 (n24582, n_21175, n_21176);
  not g45375 (n_21177, n24581);
  not g45376 (n_21178, n24582);
  and g45377 (n24583, n_21177, n_21178);
  not g45378 (n_21179, n24583);
  and g45379 (n24584, n24572, n_21179);
  not g45380 (n_21180, n24584);
  and g45381 (n24585, n24572, n_21180);
  and g45382 (n24586, n_21179, n_21180);
  not g45383 (n_21181, n24585);
  not g45384 (n_21182, n24586);
  and g45385 (n24587, n_21181, n_21182);
  and g45386 (n24588, n_21007, n_21017);
  and g45387 (n24589, n24587, n24588);
  not g45388 (n_21183, n24587);
  not g45389 (n_21184, n24588);
  and g45390 (n24590, n_21183, n_21184);
  not g45391 (n_21185, n24589);
  not g45392 (n_21186, n24590);
  and g45393 (n24591, n_21185, n_21186);
  and g45394 (n24592, n_21020, n_21021);
  not g45395 (n_21187, n24592);
  and g45396 (n24593, n_20870, n_21187);
  not g45397 (n_21188, n24593);
  and g45398 (n24594, n24591, n_21188);
  not g45399 (n_21189, n24591);
  and g45400 (n24595, n_21189, n24593);
  not g45401 (n_21190, n24594);
  not g45402 (n_21191, n24595);
  and g45403 (n24596, n_21190, n_21191);
  not g45404 (n_21192, n24413);
  and g45405 (n24597, n_21192, n24596);
  not g45406 (n_21193, n24596);
  and g45407 (n24598, n24413, n_21193);
  not g45408 (n_21194, n24597);
  not g45409 (n_21195, n24598);
  and g45410 (\f[99] , n_21194, n_21195);
  and g45411 (n24600, n_21164, n_21170);
  and g45412 (n24601, \b[62] , n5277);
  and g45413 (n24602, \b[63] , n5030);
  not g45414 (n_21196, n24601);
  not g45415 (n_21197, n24602);
  and g45416 (n24603, n_21196, n_21197);
  not g45417 (n_21198, n5038);
  and g45418 (n24604, n_21198, n24603);
  and g45419 (n24605, n13800, n24603);
  not g45420 (n_21199, n24604);
  not g45421 (n_21200, n24605);
  and g45422 (n24606, n_21199, n_21200);
  not g45423 (n_21201, n24606);
  and g45424 (n24607, \a[38] , n_21201);
  and g45425 (n24608, n_4202, n24606);
  not g45426 (n_21202, n24607);
  not g45427 (n_21203, n24608);
  and g45428 (n24609, n_21202, n_21203);
  not g45429 (n_21204, n24600);
  not g45430 (n_21205, n24609);
  and g45431 (n24610, n_21204, n_21205);
  and g45432 (n24611, n24600, n24609);
  not g45433 (n_21206, n24610);
  not g45434 (n_21207, n24611);
  and g45435 (n24612, n_21206, n_21207);
  and g45436 (n24613, \b[40] , n12668);
  and g45437 (n24614, \b[38] , n13047);
  and g45438 (n24615, \b[39] , n12663);
  and g45444 (n24618, n5955, n12671);
  not g45447 (n_21212, n24619);
  and g45448 (n24620, \a[62] , n_21212);
  not g45449 (n_21213, n24620);
  and g45450 (n24621, \a[62] , n_21213);
  and g45451 (n24622, n_21212, n_21213);
  not g45452 (n_21214, n24621);
  not g45453 (n_21215, n24622);
  and g45454 (n24623, n_21214, n_21215);
  and g45455 (n24624, \b[36] , n13903);
  and g45456 (n24625, \b[37] , n_11555);
  not g45457 (n_21216, n24624);
  not g45458 (n_21217, n24625);
  and g45459 (n24626, n_21216, n_21217);
  and g45460 (n24627, n_3555, n_20900);
  not g45461 (n_21218, n24627);
  and g45462 (n24628, n_21046, n_21218);
  not g45463 (n_21219, n24628);
  and g45464 (n24629, n24626, n_21219);
  not g45465 (n_21220, n24629);
  and g45466 (n24630, n24626, n_21220);
  and g45467 (n24631, n_21219, n_21220);
  not g45468 (n_21221, n24630);
  not g45469 (n_21222, n24631);
  and g45470 (n24632, n_21221, n_21222);
  not g45471 (n_21223, n24623);
  not g45472 (n_21224, n24632);
  and g45473 (n24633, n_21223, n_21224);
  not g45474 (n_21225, n24633);
  and g45475 (n24634, n_21223, n_21225);
  and g45476 (n24635, n_21224, n_21225);
  not g45477 (n_21226, n24634);
  not g45478 (n_21227, n24635);
  and g45479 (n24636, n_21226, n_21227);
  and g45480 (n24637, n_21050, n_21063);
  and g45481 (n24638, n24636, n24637);
  not g45482 (n_21228, n24636);
  not g45483 (n_21229, n24637);
  and g45484 (n24639, n_21228, n_21229);
  not g45485 (n_21230, n24638);
  not g45486 (n_21231, n24639);
  and g45487 (n24640, n_21230, n_21231);
  and g45488 (n24641, \b[43] , n11531);
  and g45489 (n24642, \b[41] , n11896);
  and g45490 (n24643, \b[42] , n11526);
  and g45496 (n24646, n6515, n11534);
  not g45499 (n_21236, n24647);
  and g45500 (n24648, \a[59] , n_21236);
  not g45501 (n_21237, n24648);
  and g45502 (n24649, \a[59] , n_21237);
  and g45503 (n24650, n_21236, n_21237);
  not g45504 (n_21238, n24649);
  not g45505 (n_21239, n24650);
  and g45506 (n24651, n_21238, n_21239);
  not g45507 (n_21240, n24651);
  and g45508 (n24652, n24640, n_21240);
  not g45509 (n_21241, n24652);
  and g45510 (n24653, n24640, n_21241);
  and g45511 (n24654, n_21240, n_21241);
  not g45512 (n_21242, n24653);
  not g45513 (n_21243, n24654);
  and g45514 (n24655, n_21242, n_21243);
  and g45515 (n24656, n_21073, n_21079);
  and g45516 (n24657, n24655, n24656);
  not g45517 (n_21244, n24655);
  not g45518 (n_21245, n24656);
  and g45519 (n24658, n_21244, n_21245);
  not g45520 (n_21246, n24657);
  not g45521 (n_21247, n24658);
  and g45522 (n24659, n_21246, n_21247);
  and g45523 (n24660, \b[46] , n10426);
  and g45524 (n24661, \b[44] , n10796);
  and g45525 (n24662, \b[45] , n10421);
  and g45531 (n24665, n7677, n10429);
  not g45534 (n_21252, n24666);
  and g45535 (n24667, \a[56] , n_21252);
  not g45536 (n_21253, n24667);
  and g45537 (n24668, \a[56] , n_21253);
  and g45538 (n24669, n_21252, n_21253);
  not g45539 (n_21254, n24668);
  not g45540 (n_21255, n24669);
  and g45541 (n24670, n_21254, n_21255);
  not g45542 (n_21256, n24670);
  and g45543 (n24671, n24659, n_21256);
  not g45544 (n_21257, n24671);
  and g45545 (n24672, n24659, n_21257);
  and g45546 (n24673, n_21256, n_21257);
  not g45547 (n_21258, n24672);
  not g45548 (n_21259, n24673);
  and g45549 (n24674, n_21258, n_21259);
  and g45550 (n24675, n_21092, n_21098);
  and g45551 (n24676, n24674, n24675);
  not g45552 (n_21260, n24674);
  not g45553 (n_21261, n24675);
  and g45554 (n24677, n_21260, n_21261);
  not g45555 (n_21262, n24676);
  not g45556 (n_21263, n24677);
  and g45557 (n24678, n_21262, n_21263);
  and g45558 (n24679, \b[49] , n9339);
  and g45559 (n24680, \b[47] , n9732);
  and g45560 (n24681, \b[48] , n9334);
  and g45566 (n24684, n8625, n9342);
  not g45569 (n_21268, n24685);
  and g45570 (n24686, \a[53] , n_21268);
  not g45571 (n_21269, n24686);
  and g45572 (n24687, \a[53] , n_21269);
  and g45573 (n24688, n_21268, n_21269);
  not g45574 (n_21270, n24687);
  not g45575 (n_21271, n24688);
  and g45576 (n24689, n_21270, n_21271);
  not g45577 (n_21272, n24689);
  and g45578 (n24690, n24678, n_21272);
  not g45579 (n_21273, n24690);
  and g45580 (n24691, n24678, n_21273);
  and g45581 (n24692, n_21272, n_21273);
  not g45582 (n_21274, n24691);
  not g45583 (n_21275, n24692);
  and g45584 (n24693, n_21274, n_21275);
  and g45585 (n24694, n_21108, n_21114);
  and g45586 (n24695, n24693, n24694);
  not g45587 (n_21276, n24693);
  not g45588 (n_21277, n24694);
  and g45589 (n24696, n_21276, n_21277);
  not g45590 (n_21278, n24695);
  not g45591 (n_21279, n24696);
  and g45592 (n24697, n_21278, n_21279);
  and g45593 (n24698, \b[52] , n8362);
  and g45594 (n24699, \b[50] , n8715);
  and g45595 (n24700, \b[51] , n8357);
  and g45601 (n24703, n8365, n9628);
  not g45604 (n_21284, n24704);
  and g45605 (n24705, \a[50] , n_21284);
  not g45606 (n_21285, n24705);
  and g45607 (n24706, \a[50] , n_21285);
  and g45608 (n24707, n_21284, n_21285);
  not g45609 (n_21286, n24706);
  not g45610 (n_21287, n24707);
  and g45611 (n24708, n_21286, n_21287);
  not g45612 (n_21288, n24708);
  and g45613 (n24709, n24697, n_21288);
  not g45614 (n_21289, n24709);
  and g45615 (n24710, n24697, n_21289);
  and g45616 (n24711, n_21288, n_21289);
  not g45617 (n_21290, n24710);
  not g45618 (n_21291, n24711);
  and g45619 (n24712, n_21290, n_21291);
  and g45620 (n24713, n_21126, n_21129);
  not g45621 (n_21292, n24712);
  not g45622 (n_21293, n24713);
  and g45623 (n24714, n_21292, n_21293);
  not g45624 (n_21294, n24714);
  and g45625 (n24715, n_21292, n_21294);
  and g45626 (n24716, n_21293, n_21294);
  not g45627 (n_21295, n24715);
  not g45628 (n_21296, n24716);
  and g45629 (n24717, n_21295, n_21296);
  and g45630 (n24718, \b[55] , n7446);
  and g45631 (n24719, \b[53] , n7787);
  and g45632 (n24720, \b[54] , n7441);
  and g45638 (n24723, n7449, n10684);
  not g45641 (n_21301, n24724);
  and g45642 (n24725, \a[47] , n_21301);
  not g45643 (n_21302, n24725);
  and g45644 (n24726, \a[47] , n_21302);
  and g45645 (n24727, n_21301, n_21302);
  not g45646 (n_21303, n24726);
  not g45647 (n_21304, n24727);
  and g45648 (n24728, n_21303, n_21304);
  not g45649 (n_21305, n24717);
  not g45650 (n_21306, n24728);
  and g45651 (n24729, n_21305, n_21306);
  not g45652 (n_21307, n24729);
  and g45653 (n24730, n_21305, n_21307);
  and g45654 (n24731, n_21306, n_21307);
  not g45655 (n_21308, n24730);
  not g45656 (n_21309, n24731);
  and g45657 (n24732, n_21308, n_21309);
  and g45658 (n24733, n_21133, n_21137);
  and g45659 (n24734, n24732, n24733);
  not g45660 (n_21310, n24732);
  not g45661 (n_21311, n24733);
  and g45662 (n24735, n_21310, n_21311);
  not g45663 (n_21312, n24734);
  not g45664 (n_21313, n24735);
  and g45665 (n24736, n_21312, n_21313);
  and g45666 (n24737, \b[58] , n6595);
  and g45667 (n24738, \b[56] , n6902);
  and g45668 (n24739, \b[57] , n6590);
  and g45674 (n24742, n6598, n11436);
  not g45677 (n_21318, n24743);
  and g45678 (n24744, \a[44] , n_21318);
  not g45679 (n_21319, n24744);
  and g45680 (n24745, \a[44] , n_21319);
  and g45681 (n24746, n_21318, n_21319);
  not g45682 (n_21320, n24745);
  not g45683 (n_21321, n24746);
  and g45684 (n24747, n_21320, n_21321);
  not g45685 (n_21322, n24747);
  and g45686 (n24748, n24736, n_21322);
  not g45687 (n_21323, n24748);
  and g45688 (n24749, n24736, n_21323);
  and g45689 (n24750, n_21322, n_21323);
  not g45690 (n_21324, n24749);
  not g45691 (n_21325, n24750);
  and g45692 (n24751, n_21324, n_21325);
  and g45693 (n24752, n_21148, n_21154);
  and g45694 (n24753, n24751, n24752);
  not g45695 (n_21326, n24751);
  not g45696 (n_21327, n24752);
  and g45697 (n24754, n_21326, n_21327);
  not g45698 (n_21328, n24753);
  not g45699 (n_21329, n24754);
  and g45700 (n24755, n_21328, n_21329);
  and g45701 (n24756, \b[61] , n5777);
  and g45702 (n24757, \b[59] , n6059);
  and g45703 (n24758, \b[60] , n5772);
  and g45709 (n24761, n5780, n12969);
  not g45712 (n_21334, n24762);
  and g45713 (n24763, \a[41] , n_21334);
  not g45714 (n_21335, n24763);
  and g45715 (n24764, \a[41] , n_21335);
  and g45716 (n24765, n_21334, n_21335);
  not g45717 (n_21336, n24764);
  not g45718 (n_21337, n24765);
  and g45719 (n24766, n_21336, n_21337);
  not g45720 (n_21338, n24766);
  and g45721 (n24767, n24755, n_21338);
  not g45722 (n_21339, n24755);
  and g45723 (n24768, n_21339, n24766);
  not g45724 (n_21340, n24768);
  and g45725 (n24769, n24612, n_21340);
  not g45726 (n_21341, n24767);
  and g45727 (n24770, n_21341, n24769);
  not g45728 (n_21342, n24770);
  and g45729 (n24771, n24612, n_21342);
  and g45730 (n24772, n_21340, n_21342);
  and g45731 (n24773, n_21341, n24772);
  not g45732 (n_21343, n24771);
  not g45733 (n_21344, n24773);
  and g45734 (n24774, n_21343, n_21344);
  and g45735 (n24775, n_21180, n_21186);
  and g45736 (n24776, n24774, n24775);
  not g45737 (n_21345, n24774);
  not g45738 (n_21346, n24775);
  and g45739 (n24777, n_21345, n_21346);
  not g45740 (n_21347, n24776);
  not g45741 (n_21348, n24777);
  and g45742 (n24778, n_21347, n_21348);
  and g45743 (n24779, n_21190, n_21194);
  not g45744 (n_21349, n24779);
  and g45745 (n24780, n24778, n_21349);
  not g45746 (n_21350, n24778);
  and g45747 (n24781, n_21350, n24779);
  not g45748 (n_21351, n24780);
  not g45749 (n_21352, n24781);
  and g45750 (\f[100] , n_21351, n_21352);
  and g45751 (n24783, n_21348, n_21351);
  and g45752 (n24784, n_21206, n_21342);
  and g45753 (n24785, n_21329, n_21341);
  and g45754 (n24786, \b[63] , n5277);
  and g45755 (n24787, n5038, n13797);
  not g45756 (n_21353, n24786);
  not g45757 (n_21354, n24787);
  and g45758 (n24788, n_21353, n_21354);
  not g45759 (n_21355, n24788);
  and g45760 (n24789, \a[38] , n_21355);
  not g45761 (n_21356, n24789);
  and g45762 (n24790, \a[38] , n_21356);
  and g45763 (n24791, n_21355, n_21356);
  not g45764 (n_21357, n24790);
  not g45765 (n_21358, n24791);
  and g45766 (n24792, n_21357, n_21358);
  not g45767 (n_21359, n24785);
  not g45768 (n_21360, n24792);
  and g45769 (n24793, n_21359, n_21360);
  not g45770 (n_21361, n24793);
  and g45771 (n24794, n_21359, n_21361);
  and g45772 (n24795, n_21360, n_21361);
  not g45773 (n_21362, n24794);
  not g45774 (n_21363, n24795);
  and g45775 (n24796, n_21362, n_21363);
  and g45776 (n24797, n_21294, n_21307);
  and g45777 (n24798, \b[56] , n7446);
  and g45778 (n24799, \b[54] , n7787);
  and g45779 (n24800, \b[55] , n7441);
  and g45785 (n24803, n7449, n10708);
  not g45788 (n_21368, n24804);
  and g45789 (n24805, \a[47] , n_21368);
  not g45790 (n_21369, n24805);
  and g45791 (n24806, \a[47] , n_21369);
  and g45792 (n24807, n_21368, n_21369);
  not g45793 (n_21370, n24806);
  not g45794 (n_21371, n24807);
  and g45795 (n24808, n_21370, n_21371);
  and g45796 (n24809, n_21279, n_21289);
  and g45797 (n24810, \b[53] , n8362);
  and g45798 (n24811, \b[51] , n8715);
  and g45799 (n24812, \b[52] , n8357);
  and g45805 (n24815, n8365, n9972);
  not g45808 (n_21376, n24816);
  and g45809 (n24817, \a[50] , n_21376);
  not g45810 (n_21377, n24817);
  and g45811 (n24818, \a[50] , n_21377);
  and g45812 (n24819, n_21376, n_21377);
  not g45813 (n_21378, n24818);
  not g45814 (n_21379, n24819);
  and g45815 (n24820, n_21378, n_21379);
  and g45816 (n24821, n_21263, n_21273);
  and g45817 (n24822, n_21220, n_21225);
  and g45818 (n24823, \b[37] , n13903);
  and g45819 (n24824, \b[38] , n_11555);
  not g45820 (n_21380, n24823);
  not g45821 (n_21381, n24824);
  and g45822 (n24825, n_21380, n_21381);
  not g45823 (n_21382, n24825);
  and g45824 (n24826, n24626, n_21382);
  not g45825 (n_21383, n24826);
  and g45826 (n24827, n24626, n_21383);
  and g45827 (n24828, n_21382, n_21383);
  not g45828 (n_21384, n24827);
  not g45829 (n_21385, n24828);
  and g45830 (n24829, n_21384, n_21385);
  not g45831 (n_21386, n24822);
  not g45832 (n_21387, n24829);
  and g45833 (n24830, n_21386, n_21387);
  not g45834 (n_21388, n24830);
  and g45835 (n24831, n_21386, n_21388);
  and g45836 (n24832, n_21387, n_21388);
  not g45837 (n_21389, n24831);
  not g45838 (n_21390, n24832);
  and g45839 (n24833, n_21389, n_21390);
  and g45840 (n24834, \b[41] , n12668);
  and g45841 (n24835, \b[39] , n13047);
  and g45842 (n24836, \b[40] , n12663);
  and g45848 (n24839, n6219, n12671);
  not g45851 (n_21395, n24840);
  and g45852 (n24841, \a[62] , n_21395);
  not g45853 (n_21396, n24841);
  and g45854 (n24842, \a[62] , n_21396);
  and g45855 (n24843, n_21395, n_21396);
  not g45856 (n_21397, n24842);
  not g45857 (n_21398, n24843);
  and g45858 (n24844, n_21397, n_21398);
  not g45859 (n_21399, n24833);
  not g45860 (n_21400, n24844);
  and g45861 (n24845, n_21399, n_21400);
  not g45862 (n_21401, n24845);
  and g45863 (n24846, n_21399, n_21401);
  and g45864 (n24847, n_21400, n_21401);
  not g45865 (n_21402, n24846);
  not g45866 (n_21403, n24847);
  and g45867 (n24848, n_21402, n_21403);
  and g45868 (n24849, \b[44] , n11531);
  and g45869 (n24850, \b[42] , n11896);
  and g45870 (n24851, \b[43] , n11526);
  and g45876 (n24854, n7072, n11534);
  not g45879 (n_21408, n24855);
  and g45880 (n24856, \a[59] , n_21408);
  not g45881 (n_21409, n24856);
  and g45882 (n24857, \a[59] , n_21409);
  and g45883 (n24858, n_21408, n_21409);
  not g45884 (n_21410, n24857);
  not g45885 (n_21411, n24858);
  and g45886 (n24859, n_21410, n_21411);
  not g45887 (n_21412, n24848);
  and g45888 (n24860, n_21412, n24859);
  not g45889 (n_21413, n24859);
  and g45890 (n24861, n24848, n_21413);
  not g45891 (n_21414, n24860);
  not g45892 (n_21415, n24861);
  and g45893 (n24862, n_21414, n_21415);
  and g45894 (n24863, n_21231, n_21241);
  and g45895 (n24864, n24862, n24863);
  not g45896 (n_21416, n24862);
  not g45897 (n_21417, n24863);
  and g45898 (n24865, n_21416, n_21417);
  not g45899 (n_21418, n24864);
  not g45900 (n_21419, n24865);
  and g45901 (n24866, n_21418, n_21419);
  and g45902 (n24867, \b[47] , n10426);
  and g45903 (n24868, \b[45] , n10796);
  and g45904 (n24869, \b[46] , n10421);
  and g45910 (n24872, n7703, n10429);
  not g45913 (n_21424, n24873);
  and g45914 (n24874, \a[56] , n_21424);
  not g45915 (n_21425, n24874);
  and g45916 (n24875, \a[56] , n_21425);
  and g45917 (n24876, n_21424, n_21425);
  not g45918 (n_21426, n24875);
  not g45919 (n_21427, n24876);
  and g45920 (n24877, n_21426, n_21427);
  not g45921 (n_21428, n24877);
  and g45922 (n24878, n24866, n_21428);
  not g45923 (n_21429, n24878);
  and g45924 (n24879, n24866, n_21429);
  and g45925 (n24880, n_21428, n_21429);
  not g45926 (n_21430, n24879);
  not g45927 (n_21431, n24880);
  and g45928 (n24881, n_21430, n_21431);
  and g45929 (n24882, n_21247, n_21257);
  and g45930 (n24883, n24881, n24882);
  not g45931 (n_21432, n24881);
  not g45932 (n_21433, n24882);
  and g45933 (n24884, n_21432, n_21433);
  not g45934 (n_21434, n24883);
  not g45935 (n_21435, n24884);
  and g45936 (n24885, n_21434, n_21435);
  and g45937 (n24886, \b[50] , n9339);
  and g45938 (n24887, \b[48] , n9732);
  and g45939 (n24888, \b[49] , n9334);
  and g45945 (n24891, n8949, n9342);
  not g45948 (n_21440, n24892);
  and g45949 (n24893, \a[53] , n_21440);
  not g45950 (n_21441, n24893);
  and g45951 (n24894, \a[53] , n_21441);
  and g45952 (n24895, n_21440, n_21441);
  not g45953 (n_21442, n24894);
  not g45954 (n_21443, n24895);
  and g45955 (n24896, n_21442, n_21443);
  not g45956 (n_21444, n24885);
  and g45957 (n24897, n_21444, n24896);
  not g45958 (n_21445, n24896);
  and g45959 (n24898, n24885, n_21445);
  not g45960 (n_21446, n24897);
  not g45961 (n_21447, n24898);
  and g45962 (n24899, n_21446, n_21447);
  not g45963 (n_21448, n24821);
  and g45964 (n24900, n_21448, n24899);
  not g45965 (n_21449, n24900);
  and g45966 (n24901, n_21448, n_21449);
  and g45967 (n24902, n24899, n_21449);
  not g45968 (n_21450, n24901);
  not g45969 (n_21451, n24902);
  and g45970 (n24903, n_21450, n_21451);
  not g45971 (n_21452, n24820);
  not g45972 (n_21453, n24903);
  and g45973 (n24904, n_21452, n_21453);
  and g45974 (n24905, n24820, n_21451);
  and g45975 (n24906, n_21450, n24905);
  not g45976 (n_21454, n24904);
  not g45977 (n_21455, n24906);
  and g45978 (n24907, n_21454, n_21455);
  not g45979 (n_21456, n24809);
  and g45980 (n24908, n_21456, n24907);
  not g45981 (n_21457, n24907);
  and g45982 (n24909, n24809, n_21457);
  not g45983 (n_21458, n24908);
  not g45984 (n_21459, n24909);
  and g45985 (n24910, n_21458, n_21459);
  not g45986 (n_21460, n24808);
  and g45987 (n24911, n_21460, n24910);
  not g45988 (n_21461, n24910);
  and g45989 (n24912, n24808, n_21461);
  not g45990 (n_21462, n24911);
  not g45991 (n_21463, n24912);
  and g45992 (n24913, n_21462, n_21463);
  not g45993 (n_21464, n24797);
  and g45994 (n24914, n_21464, n24913);
  not g45995 (n_21465, n24913);
  and g45996 (n24915, n24797, n_21465);
  not g45997 (n_21466, n24914);
  not g45998 (n_21467, n24915);
  and g45999 (n24916, n_21466, n_21467);
  and g46000 (n24917, \b[59] , n6595);
  and g46001 (n24918, \b[57] , n6902);
  and g46002 (n24919, \b[58] , n6590);
  and g46008 (n24922, n6598, n12179);
  not g46011 (n_21472, n24923);
  and g46012 (n24924, \a[44] , n_21472);
  not g46013 (n_21473, n24924);
  and g46014 (n24925, \a[44] , n_21473);
  and g46015 (n24926, n_21472, n_21473);
  not g46016 (n_21474, n24925);
  not g46017 (n_21475, n24926);
  and g46018 (n24927, n_21474, n_21475);
  not g46019 (n_21476, n24927);
  and g46020 (n24928, n24916, n_21476);
  not g46021 (n_21477, n24928);
  and g46022 (n24929, n24916, n_21477);
  and g46023 (n24930, n_21476, n_21477);
  not g46024 (n_21478, n24929);
  not g46025 (n_21479, n24930);
  and g46026 (n24931, n_21478, n_21479);
  and g46027 (n24932, n_21313, n_21323);
  and g46028 (n24933, n24931, n24932);
  not g46029 (n_21480, n24931);
  not g46030 (n_21481, n24932);
  and g46031 (n24934, n_21480, n_21481);
  not g46032 (n_21482, n24933);
  not g46033 (n_21483, n24934);
  and g46034 (n24935, n_21482, n_21483);
  and g46035 (n24936, \b[62] , n5777);
  and g46036 (n24937, \b[60] , n6059);
  and g46037 (n24938, \b[61] , n5772);
  and g46043 (n24941, n5780, n13370);
  not g46046 (n_21488, n24942);
  and g46047 (n24943, \a[41] , n_21488);
  not g46048 (n_21489, n24943);
  and g46049 (n24944, \a[41] , n_21489);
  and g46050 (n24945, n_21488, n_21489);
  not g46051 (n_21490, n24944);
  not g46052 (n_21491, n24945);
  and g46053 (n24946, n_21490, n_21491);
  not g46054 (n_21492, n24946);
  and g46055 (n24947, n24935, n_21492);
  not g46056 (n_21493, n24947);
  and g46057 (n24948, n24935, n_21493);
  and g46058 (n24949, n_21492, n_21493);
  not g46059 (n_21494, n24948);
  not g46060 (n_21495, n24949);
  and g46061 (n24950, n_21494, n_21495);
  not g46062 (n_21496, n24796);
  and g46063 (n24951, n_21496, n24950);
  not g46064 (n_21497, n24950);
  and g46065 (n24952, n24796, n_21497);
  not g46066 (n_21498, n24951);
  not g46067 (n_21499, n24952);
  and g46068 (n24953, n_21498, n_21499);
  not g46069 (n_21500, n24784);
  not g46070 (n_21501, n24953);
  and g46071 (n24954, n_21500, n_21501);
  and g46072 (n24955, n24784, n24953);
  not g46073 (n_21502, n24954);
  not g46074 (n_21503, n24955);
  and g46075 (n24956, n_21502, n_21503);
  not g46076 (n_21504, n24783);
  and g46077 (n24957, n_21504, n24956);
  not g46078 (n_21505, n24956);
  and g46079 (n24958, n24783, n_21505);
  not g46080 (n_21506, n24957);
  not g46081 (n_21507, n24958);
  and g46082 (\f[101] , n_21506, n_21507);
  and g46083 (n24960, n_21502, n_21506);
  and g46084 (n24961, n_21449, n_21454);
  and g46085 (n24962, \b[54] , n8362);
  and g46086 (n24963, \b[52] , n8715);
  and g46087 (n24964, \b[53] , n8357);
  and g46093 (n24967, n8365, n9998);
  not g46096 (n_21512, n24968);
  and g46097 (n24969, \a[50] , n_21512);
  not g46098 (n_21513, n24969);
  and g46099 (n24970, \a[50] , n_21513);
  and g46100 (n24971, n_21512, n_21513);
  not g46101 (n_21514, n24970);
  not g46102 (n_21515, n24971);
  and g46103 (n24972, n_21514, n_21515);
  and g46104 (n24973, n_21435, n_21447);
  and g46105 (n24974, n_21383, n_21388);
  and g46106 (n24975, \b[38] , n13903);
  and g46107 (n24976, \b[39] , n_11555);
  not g46108 (n_21516, n24975);
  not g46109 (n_21517, n24976);
  and g46110 (n24977, n_21516, n_21517);
  not g46111 (n_21518, n24626);
  and g46112 (n24978, \a[38] , n_21518);
  and g46113 (n24979, n_4202, n24626);
  not g46114 (n_21519, n24978);
  not g46115 (n_21520, n24979);
  and g46116 (n24980, n_21519, n_21520);
  not g46117 (n_21521, n24977);
  not g46118 (n_21522, n24980);
  and g46119 (n24981, n_21521, n_21522);
  and g46120 (n24982, n24977, n24980);
  not g46121 (n_21523, n24981);
  not g46122 (n_21524, n24982);
  and g46123 (n24983, n_21523, n_21524);
  not g46124 (n_21525, n24974);
  and g46125 (n24984, n_21525, n24983);
  not g46126 (n_21526, n24983);
  and g46127 (n24985, n24974, n_21526);
  not g46128 (n_21527, n24984);
  not g46129 (n_21528, n24985);
  and g46130 (n24986, n_21527, n_21528);
  and g46131 (n24987, \b[42] , n12668);
  and g46132 (n24988, \b[40] , n13047);
  and g46133 (n24989, \b[41] , n12663);
  and g46139 (n24992, n6489, n12671);
  not g46142 (n_21533, n24993);
  and g46143 (n24994, \a[62] , n_21533);
  not g46144 (n_21534, n24994);
  and g46145 (n24995, \a[62] , n_21534);
  and g46146 (n24996, n_21533, n_21534);
  not g46147 (n_21535, n24995);
  not g46148 (n_21536, n24996);
  and g46149 (n24997, n_21535, n_21536);
  not g46150 (n_21537, n24997);
  and g46151 (n24998, n24986, n_21537);
  not g46152 (n_21538, n24998);
  and g46153 (n24999, n24986, n_21538);
  and g46154 (n25000, n_21537, n_21538);
  not g46155 (n_21539, n24999);
  not g46156 (n_21540, n25000);
  and g46157 (n25001, n_21539, n_21540);
  and g46158 (n25002, \b[45] , n11531);
  and g46159 (n25003, \b[43] , n11896);
  and g46160 (n25004, \b[44] , n11526);
  and g46166 (n25007, n7361, n11534);
  not g46169 (n_21545, n25008);
  and g46170 (n25009, \a[59] , n_21545);
  not g46171 (n_21546, n25009);
  and g46172 (n25010, \a[59] , n_21546);
  and g46173 (n25011, n_21545, n_21546);
  not g46174 (n_21547, n25010);
  not g46175 (n_21548, n25011);
  and g46176 (n25012, n_21547, n_21548);
  not g46177 (n_21549, n25001);
  not g46178 (n_21550, n25012);
  and g46179 (n25013, n_21549, n_21550);
  not g46180 (n_21551, n25013);
  and g46181 (n25014, n_21549, n_21551);
  and g46182 (n25015, n_21550, n_21551);
  not g46183 (n_21552, n25014);
  not g46184 (n_21553, n25015);
  and g46185 (n25016, n_21552, n_21553);
  and g46186 (n25017, n_21412, n_21413);
  not g46187 (n_21554, n25017);
  and g46188 (n25018, n_21401, n_21554);
  not g46189 (n_21555, n25016);
  not g46190 (n_21556, n25018);
  and g46191 (n25019, n_21555, n_21556);
  not g46192 (n_21557, n25019);
  and g46193 (n25020, n_21555, n_21557);
  and g46194 (n25021, n_21556, n_21557);
  not g46195 (n_21558, n25020);
  not g46196 (n_21559, n25021);
  and g46197 (n25022, n_21558, n_21559);
  and g46198 (n25023, \b[48] , n10426);
  and g46199 (n25024, \b[46] , n10796);
  and g46200 (n25025, \b[47] , n10421);
  and g46206 (n25028, n8009, n10429);
  not g46209 (n_21564, n25029);
  and g46210 (n25030, \a[56] , n_21564);
  not g46211 (n_21565, n25030);
  and g46212 (n25031, \a[56] , n_21565);
  and g46213 (n25032, n_21564, n_21565);
  not g46214 (n_21566, n25031);
  not g46215 (n_21567, n25032);
  and g46216 (n25033, n_21566, n_21567);
  not g46217 (n_21568, n25022);
  not g46218 (n_21569, n25033);
  and g46219 (n25034, n_21568, n_21569);
  not g46220 (n_21570, n25034);
  and g46221 (n25035, n_21568, n_21570);
  and g46222 (n25036, n_21569, n_21570);
  not g46223 (n_21571, n25035);
  not g46224 (n_21572, n25036);
  and g46225 (n25037, n_21571, n_21572);
  and g46226 (n25038, n_21419, n_21429);
  and g46227 (n25039, n25037, n25038);
  not g46228 (n_21573, n25037);
  not g46229 (n_21574, n25038);
  and g46230 (n25040, n_21573, n_21574);
  not g46231 (n_21575, n25039);
  not g46232 (n_21576, n25040);
  and g46233 (n25041, n_21575, n_21576);
  and g46234 (n25042, \b[51] , n9339);
  and g46235 (n25043, \b[49] , n9732);
  and g46236 (n25044, \b[50] , n9334);
  and g46242 (n25047, n8976, n9342);
  not g46245 (n_21581, n25048);
  and g46246 (n25049, \a[53] , n_21581);
  not g46247 (n_21582, n25049);
  and g46248 (n25050, \a[53] , n_21582);
  and g46249 (n25051, n_21581, n_21582);
  not g46250 (n_21583, n25050);
  not g46251 (n_21584, n25051);
  and g46252 (n25052, n_21583, n_21584);
  not g46253 (n_21585, n25041);
  and g46254 (n25053, n_21585, n25052);
  not g46255 (n_21586, n25052);
  and g46256 (n25054, n25041, n_21586);
  not g46257 (n_21587, n25053);
  not g46258 (n_21588, n25054);
  and g46259 (n25055, n_21587, n_21588);
  not g46260 (n_21589, n24973);
  and g46261 (n25056, n_21589, n25055);
  not g46262 (n_21590, n25055);
  and g46263 (n25057, n24973, n_21590);
  not g46264 (n_21591, n25056);
  not g46265 (n_21592, n25057);
  and g46266 (n25058, n_21591, n_21592);
  not g46267 (n_21593, n24972);
  and g46268 (n25059, n_21593, n25058);
  not g46269 (n_21594, n25058);
  and g46270 (n25060, n24972, n_21594);
  not g46271 (n_21595, n25059);
  not g46272 (n_21596, n25060);
  and g46273 (n25061, n_21595, n_21596);
  not g46274 (n_21597, n24961);
  and g46275 (n25062, n_21597, n25061);
  not g46276 (n_21598, n25061);
  and g46277 (n25063, n24961, n_21598);
  not g46278 (n_21599, n25062);
  not g46279 (n_21600, n25063);
  and g46280 (n25064, n_21599, n_21600);
  and g46281 (n25065, \b[57] , n7446);
  and g46282 (n25066, \b[55] , n7787);
  and g46283 (n25067, \b[56] , n7441);
  and g46289 (n25070, n7449, n11410);
  not g46292 (n_21605, n25071);
  and g46293 (n25072, \a[47] , n_21605);
  not g46294 (n_21606, n25072);
  and g46295 (n25073, \a[47] , n_21606);
  and g46296 (n25074, n_21605, n_21606);
  not g46297 (n_21607, n25073);
  not g46298 (n_21608, n25074);
  and g46299 (n25075, n_21607, n_21608);
  not g46300 (n_21609, n25075);
  and g46301 (n25076, n25064, n_21609);
  not g46302 (n_21610, n25076);
  and g46303 (n25077, n25064, n_21610);
  and g46304 (n25078, n_21609, n_21610);
  not g46305 (n_21611, n25077);
  not g46306 (n_21612, n25078);
  and g46307 (n25079, n_21611, n_21612);
  and g46308 (n25080, n_21458, n_21462);
  and g46309 (n25081, n25079, n25080);
  not g46310 (n_21613, n25079);
  not g46311 (n_21614, n25080);
  and g46312 (n25082, n_21613, n_21614);
  not g46313 (n_21615, n25081);
  not g46314 (n_21616, n25082);
  and g46315 (n25083, n_21615, n_21616);
  and g46316 (n25084, \b[60] , n6595);
  and g46317 (n25085, \b[58] , n6902);
  and g46318 (n25086, \b[59] , n6590);
  and g46324 (n25089, n6598, n12211);
  not g46327 (n_21621, n25090);
  and g46328 (n25091, \a[44] , n_21621);
  not g46329 (n_21622, n25091);
  and g46330 (n25092, \a[44] , n_21622);
  and g46331 (n25093, n_21621, n_21622);
  not g46332 (n_21623, n25092);
  not g46333 (n_21624, n25093);
  and g46334 (n25094, n_21623, n_21624);
  not g46335 (n_21625, n25094);
  and g46336 (n25095, n25083, n_21625);
  not g46337 (n_21626, n25095);
  and g46338 (n25096, n25083, n_21626);
  and g46339 (n25097, n_21625, n_21626);
  not g46340 (n_21627, n25096);
  not g46341 (n_21628, n25097);
  and g46342 (n25098, n_21627, n_21628);
  and g46343 (n25099, n_21466, n_21477);
  and g46344 (n25100, n25098, n25099);
  not g46345 (n_21629, n25098);
  not g46346 (n_21630, n25099);
  and g46347 (n25101, n_21629, n_21630);
  not g46348 (n_21631, n25100);
  not g46349 (n_21632, n25101);
  and g46350 (n25102, n_21631, n_21632);
  and g46351 (n25103, \b[63] , n5777);
  and g46352 (n25104, \b[61] , n6059);
  and g46353 (n25105, \b[62] , n5772);
  and g46359 (n25108, n5780, n13771);
  not g46362 (n_21637, n25109);
  and g46363 (n25110, \a[41] , n_21637);
  not g46364 (n_21638, n25110);
  and g46365 (n25111, \a[41] , n_21638);
  and g46366 (n25112, n_21637, n_21638);
  not g46367 (n_21639, n25111);
  not g46368 (n_21640, n25112);
  and g46369 (n25113, n_21639, n_21640);
  not g46370 (n_21641, n25113);
  and g46371 (n25114, n25102, n_21641);
  not g46372 (n_21642, n25114);
  and g46373 (n25115, n25102, n_21642);
  and g46374 (n25116, n_21641, n_21642);
  not g46375 (n_21643, n25115);
  not g46376 (n_21644, n25116);
  and g46377 (n25117, n_21643, n_21644);
  and g46378 (n25118, n_21483, n_21493);
  and g46379 (n25119, n25117, n25118);
  not g46380 (n_21645, n25117);
  not g46381 (n_21646, n25118);
  and g46382 (n25120, n_21645, n_21646);
  not g46383 (n_21647, n25119);
  not g46384 (n_21648, n25120);
  and g46385 (n25121, n_21647, n_21648);
  and g46386 (n25122, n_21496, n_21497);
  not g46387 (n_21649, n25122);
  and g46388 (n25123, n_21361, n_21649);
  not g46389 (n_21650, n25123);
  and g46390 (n25124, n25121, n_21650);
  not g46391 (n_21651, n25121);
  and g46392 (n25125, n_21651, n25123);
  not g46393 (n_21652, n25124);
  not g46394 (n_21653, n25125);
  and g46395 (n25126, n_21652, n_21653);
  not g46396 (n_21654, n24960);
  and g46397 (n25127, n_21654, n25126);
  not g46398 (n_21655, n25126);
  and g46399 (n25128, n24960, n_21655);
  not g46400 (n_21656, n25127);
  not g46401 (n_21657, n25128);
  and g46402 (\f[102] , n_21656, n_21657);
  and g46403 (n25130, n_21626, n_21632);
  and g46404 (n25131, \b[62] , n6059);
  and g46405 (n25132, \b[63] , n5772);
  not g46406 (n_21658, n25131);
  not g46407 (n_21659, n25132);
  and g46408 (n25133, n_21658, n_21659);
  not g46409 (n_21660, n5780);
  and g46410 (n25134, n_21660, n25133);
  and g46411 (n25135, n13800, n25133);
  not g46412 (n_21661, n25134);
  not g46413 (n_21662, n25135);
  and g46414 (n25136, n_21661, n_21662);
  not g46415 (n_21663, n25136);
  and g46416 (n25137, \a[41] , n_21663);
  and g46417 (n25138, n_4853, n25136);
  not g46418 (n_21664, n25137);
  not g46419 (n_21665, n25138);
  and g46420 (n25139, n_21664, n_21665);
  not g46421 (n_21666, n25130);
  not g46422 (n_21667, n25139);
  and g46423 (n25140, n_21666, n_21667);
  and g46424 (n25141, n25130, n25139);
  not g46425 (n_21668, n25140);
  not g46426 (n_21669, n25141);
  and g46427 (n25142, n_21668, n_21669);
  and g46428 (n25143, n_21527, n_21538);
  and g46429 (n25144, \b[39] , n13903);
  and g46430 (n25145, \b[40] , n_11555);
  not g46431 (n_21670, n25144);
  not g46432 (n_21671, n25145);
  and g46433 (n25146, n_21670, n_21671);
  and g46434 (n25147, n_4202, n_21518);
  not g46435 (n_21672, n25147);
  and g46436 (n25148, n_21523, n_21672);
  not g46437 (n_21673, n25148);
  and g46438 (n25149, n25146, n_21673);
  not g46439 (n_21674, n25146);
  and g46440 (n25150, n_21674, n25148);
  not g46441 (n_21675, n25149);
  not g46442 (n_21676, n25150);
  and g46443 (n25151, n_21675, n_21676);
  and g46444 (n25152, \b[43] , n12668);
  and g46445 (n25153, \b[41] , n13047);
  and g46446 (n25154, \b[42] , n12663);
  not g46447 (n_21677, n25153);
  not g46448 (n_21678, n25154);
  and g46449 (n25155, n_21677, n_21678);
  not g46450 (n_21679, n25152);
  and g46451 (n25156, n_21679, n25155);
  and g46452 (n25157, n_12644, n25156);
  not g46453 (n_21680, n6515);
  and g46454 (n25158, n_21680, n25156);
  not g46455 (n_21681, n25157);
  not g46456 (n_21682, n25158);
  and g46457 (n25159, n_21681, n_21682);
  not g46458 (n_21683, n25159);
  and g46459 (n25160, \a[62] , n_21683);
  and g46460 (n25161, n_10843, n25159);
  not g46461 (n_21684, n25160);
  not g46462 (n_21685, n25161);
  and g46463 (n25162, n_21684, n_21685);
  not g46464 (n_21686, n25162);
  and g46465 (n25163, n25151, n_21686);
  not g46466 (n_21687, n25151);
  and g46467 (n25164, n_21687, n25162);
  not g46468 (n_21688, n25163);
  not g46469 (n_21689, n25164);
  and g46470 (n25165, n_21688, n_21689);
  not g46471 (n_21690, n25143);
  and g46472 (n25166, n_21690, n25165);
  not g46473 (n_21691, n25165);
  and g46474 (n25167, n25143, n_21691);
  not g46475 (n_21692, n25166);
  not g46476 (n_21693, n25167);
  and g46477 (n25168, n_21692, n_21693);
  and g46478 (n25169, \b[46] , n11531);
  and g46479 (n25170, \b[44] , n11896);
  and g46480 (n25171, \b[45] , n11526);
  and g46486 (n25174, n7677, n11534);
  not g46489 (n_21698, n25175);
  and g46490 (n25176, \a[59] , n_21698);
  not g46491 (n_21699, n25176);
  and g46492 (n25177, \a[59] , n_21699);
  and g46493 (n25178, n_21698, n_21699);
  not g46494 (n_21700, n25177);
  not g46495 (n_21701, n25178);
  and g46496 (n25179, n_21700, n_21701);
  not g46497 (n_21702, n25179);
  and g46498 (n25180, n25168, n_21702);
  not g46499 (n_21703, n25180);
  and g46500 (n25181, n25168, n_21703);
  and g46501 (n25182, n_21702, n_21703);
  not g46502 (n_21704, n25181);
  not g46503 (n_21705, n25182);
  and g46504 (n25183, n_21704, n_21705);
  and g46505 (n25184, n_21551, n_21557);
  and g46506 (n25185, n25183, n25184);
  not g46507 (n_21706, n25183);
  not g46508 (n_21707, n25184);
  and g46509 (n25186, n_21706, n_21707);
  not g46510 (n_21708, n25185);
  not g46511 (n_21709, n25186);
  and g46512 (n25187, n_21708, n_21709);
  and g46513 (n25188, \b[49] , n10426);
  and g46514 (n25189, \b[47] , n10796);
  and g46515 (n25190, \b[48] , n10421);
  and g46521 (n25193, n8625, n10429);
  not g46524 (n_21714, n25194);
  and g46525 (n25195, \a[56] , n_21714);
  not g46526 (n_21715, n25195);
  and g46527 (n25196, \a[56] , n_21715);
  and g46528 (n25197, n_21714, n_21715);
  not g46529 (n_21716, n25196);
  not g46530 (n_21717, n25197);
  and g46531 (n25198, n_21716, n_21717);
  not g46532 (n_21718, n25198);
  and g46533 (n25199, n25187, n_21718);
  not g46534 (n_21719, n25199);
  and g46535 (n25200, n25187, n_21719);
  and g46536 (n25201, n_21718, n_21719);
  not g46537 (n_21720, n25200);
  not g46538 (n_21721, n25201);
  and g46539 (n25202, n_21720, n_21721);
  and g46540 (n25203, n_21570, n_21576);
  and g46541 (n25204, n25202, n25203);
  not g46542 (n_21722, n25202);
  not g46543 (n_21723, n25203);
  and g46544 (n25205, n_21722, n_21723);
  not g46545 (n_21724, n25204);
  not g46546 (n_21725, n25205);
  and g46547 (n25206, n_21724, n_21725);
  and g46548 (n25207, \b[52] , n9339);
  and g46549 (n25208, \b[50] , n9732);
  and g46550 (n25209, \b[51] , n9334);
  and g46556 (n25212, n9342, n9628);
  not g46559 (n_21730, n25213);
  and g46560 (n25214, \a[53] , n_21730);
  not g46561 (n_21731, n25214);
  and g46562 (n25215, \a[53] , n_21731);
  and g46563 (n25216, n_21730, n_21731);
  not g46564 (n_21732, n25215);
  not g46565 (n_21733, n25216);
  and g46566 (n25217, n_21732, n_21733);
  not g46567 (n_21734, n25217);
  and g46568 (n25218, n25206, n_21734);
  not g46569 (n_21735, n25218);
  and g46570 (n25219, n25206, n_21735);
  and g46571 (n25220, n_21734, n_21735);
  not g46572 (n_21736, n25219);
  not g46573 (n_21737, n25220);
  and g46574 (n25221, n_21736, n_21737);
  and g46575 (n25222, n_21588, n_21591);
  not g46576 (n_21738, n25221);
  not g46577 (n_21739, n25222);
  and g46578 (n25223, n_21738, n_21739);
  not g46579 (n_21740, n25223);
  and g46580 (n25224, n_21738, n_21740);
  and g46581 (n25225, n_21739, n_21740);
  not g46582 (n_21741, n25224);
  not g46583 (n_21742, n25225);
  and g46584 (n25226, n_21741, n_21742);
  and g46585 (n25227, \b[55] , n8362);
  and g46586 (n25228, \b[53] , n8715);
  and g46587 (n25229, \b[54] , n8357);
  and g46593 (n25232, n8365, n10684);
  not g46596 (n_21747, n25233);
  and g46597 (n25234, \a[50] , n_21747);
  not g46598 (n_21748, n25234);
  and g46599 (n25235, \a[50] , n_21748);
  and g46600 (n25236, n_21747, n_21748);
  not g46601 (n_21749, n25235);
  not g46602 (n_21750, n25236);
  and g46603 (n25237, n_21749, n_21750);
  not g46604 (n_21751, n25226);
  not g46605 (n_21752, n25237);
  and g46606 (n25238, n_21751, n_21752);
  not g46607 (n_21753, n25238);
  and g46608 (n25239, n_21751, n_21753);
  and g46609 (n25240, n_21752, n_21753);
  not g46610 (n_21754, n25239);
  not g46611 (n_21755, n25240);
  and g46612 (n25241, n_21754, n_21755);
  and g46613 (n25242, n_21595, n_21599);
  and g46614 (n25243, n25241, n25242);
  not g46615 (n_21756, n25241);
  not g46616 (n_21757, n25242);
  and g46617 (n25244, n_21756, n_21757);
  not g46618 (n_21758, n25243);
  not g46619 (n_21759, n25244);
  and g46620 (n25245, n_21758, n_21759);
  and g46621 (n25246, \b[58] , n7446);
  and g46622 (n25247, \b[56] , n7787);
  and g46623 (n25248, \b[57] , n7441);
  and g46629 (n25251, n7449, n11436);
  not g46632 (n_21764, n25252);
  and g46633 (n25253, \a[47] , n_21764);
  not g46634 (n_21765, n25253);
  and g46635 (n25254, \a[47] , n_21765);
  and g46636 (n25255, n_21764, n_21765);
  not g46637 (n_21766, n25254);
  not g46638 (n_21767, n25255);
  and g46639 (n25256, n_21766, n_21767);
  not g46640 (n_21768, n25256);
  and g46641 (n25257, n25245, n_21768);
  not g46642 (n_21769, n25257);
  and g46643 (n25258, n25245, n_21769);
  and g46644 (n25259, n_21768, n_21769);
  not g46645 (n_21770, n25258);
  not g46646 (n_21771, n25259);
  and g46647 (n25260, n_21770, n_21771);
  and g46648 (n25261, n_21610, n_21616);
  and g46649 (n25262, n25260, n25261);
  not g46650 (n_21772, n25260);
  not g46651 (n_21773, n25261);
  and g46652 (n25263, n_21772, n_21773);
  not g46653 (n_21774, n25262);
  not g46654 (n_21775, n25263);
  and g46655 (n25264, n_21774, n_21775);
  and g46656 (n25265, \b[61] , n6595);
  and g46657 (n25266, \b[59] , n6902);
  and g46658 (n25267, \b[60] , n6590);
  and g46664 (n25270, n6598, n12969);
  not g46667 (n_21780, n25271);
  and g46668 (n25272, \a[44] , n_21780);
  not g46669 (n_21781, n25272);
  and g46670 (n25273, \a[44] , n_21781);
  and g46671 (n25274, n_21780, n_21781);
  not g46672 (n_21782, n25273);
  not g46673 (n_21783, n25274);
  and g46674 (n25275, n_21782, n_21783);
  not g46675 (n_21784, n25275);
  and g46676 (n25276, n25264, n_21784);
  not g46677 (n_21785, n25264);
  and g46678 (n25277, n_21785, n25275);
  not g46679 (n_21786, n25277);
  and g46680 (n25278, n25142, n_21786);
  not g46681 (n_21787, n25276);
  and g46682 (n25279, n_21787, n25278);
  not g46683 (n_21788, n25279);
  and g46684 (n25280, n25142, n_21788);
  and g46685 (n25281, n_21786, n_21788);
  and g46686 (n25282, n_21787, n25281);
  not g46687 (n_21789, n25280);
  not g46688 (n_21790, n25282);
  and g46689 (n25283, n_21789, n_21790);
  and g46690 (n25284, n_21642, n_21648);
  and g46691 (n25285, n25283, n25284);
  not g46692 (n_21791, n25283);
  not g46693 (n_21792, n25284);
  and g46694 (n25286, n_21791, n_21792);
  not g46695 (n_21793, n25285);
  not g46696 (n_21794, n25286);
  and g46697 (n25287, n_21793, n_21794);
  and g46698 (n25288, n_21652, n_21656);
  not g46699 (n_21795, n25288);
  and g46700 (n25289, n25287, n_21795);
  not g46701 (n_21796, n25287);
  and g46702 (n25290, n_21796, n25288);
  not g46703 (n_21797, n25289);
  not g46704 (n_21798, n25290);
  and g46705 (\f[103] , n_21797, n_21798);
  and g46706 (n25292, n_21794, n_21797);
  and g46707 (n25293, n_21668, n_21788);
  and g46708 (n25294, n_21775, n_21787);
  and g46709 (n25295, \b[63] , n6059);
  and g46710 (n25296, n5780, n13797);
  not g46711 (n_21799, n25295);
  not g46712 (n_21800, n25296);
  and g46713 (n25297, n_21799, n_21800);
  not g46714 (n_21801, n25297);
  and g46715 (n25298, \a[41] , n_21801);
  not g46716 (n_21802, n25298);
  and g46717 (n25299, \a[41] , n_21802);
  and g46718 (n25300, n_21801, n_21802);
  not g46719 (n_21803, n25299);
  not g46720 (n_21804, n25300);
  and g46721 (n25301, n_21803, n_21804);
  not g46722 (n_21805, n25294);
  not g46723 (n_21806, n25301);
  and g46724 (n25302, n_21805, n_21806);
  not g46725 (n_21807, n25302);
  and g46726 (n25303, n_21805, n_21807);
  and g46727 (n25304, n_21806, n_21807);
  not g46728 (n_21808, n25303);
  not g46729 (n_21809, n25304);
  and g46730 (n25305, n_21808, n_21809);
  and g46731 (n25306, \b[59] , n7446);
  and g46732 (n25307, \b[57] , n7787);
  and g46733 (n25308, \b[58] , n7441);
  and g46739 (n25311, n7449, n12179);
  not g46742 (n_21814, n25312);
  and g46743 (n25313, \a[47] , n_21814);
  not g46744 (n_21815, n25313);
  and g46745 (n25314, \a[47] , n_21815);
  and g46746 (n25315, n_21814, n_21815);
  not g46747 (n_21816, n25314);
  not g46748 (n_21817, n25315);
  and g46749 (n25316, n_21816, n_21817);
  and g46750 (n25317, n_21740, n_21753);
  and g46751 (n25318, \b[56] , n8362);
  and g46752 (n25319, \b[54] , n8715);
  and g46753 (n25320, \b[55] , n8357);
  and g46759 (n25323, n8365, n10708);
  not g46762 (n_21822, n25324);
  and g46763 (n25325, \a[50] , n_21822);
  not g46764 (n_21823, n25325);
  and g46765 (n25326, \a[50] , n_21823);
  and g46766 (n25327, n_21822, n_21823);
  not g46767 (n_21824, n25326);
  not g46768 (n_21825, n25327);
  and g46769 (n25328, n_21824, n_21825);
  and g46770 (n25329, n_21725, n_21735);
  and g46771 (n25330, \b[53] , n9339);
  and g46772 (n25331, \b[51] , n9732);
  and g46773 (n25332, \b[52] , n9334);
  and g46779 (n25335, n9342, n9972);
  not g46782 (n_21830, n25336);
  and g46783 (n25337, \a[53] , n_21830);
  not g46784 (n_21831, n25337);
  and g46785 (n25338, \a[53] , n_21831);
  and g46786 (n25339, n_21830, n_21831);
  not g46787 (n_21832, n25338);
  not g46788 (n_21833, n25339);
  and g46789 (n25340, n_21832, n_21833);
  and g46790 (n25341, n_21709, n_21719);
  and g46791 (n25342, n_21692, n_21703);
  and g46792 (n25343, n_21675, n_21688);
  and g46793 (n25344, \b[40] , n13903);
  and g46794 (n25345, \b[41] , n_11555);
  not g46795 (n_21834, n25344);
  not g46796 (n_21835, n25345);
  and g46797 (n25346, n_21834, n_21835);
  not g46798 (n_21836, n25346);
  and g46799 (n25347, n25146, n_21836);
  not g46800 (n_21837, n25347);
  and g46801 (n25348, n25146, n_21837);
  and g46802 (n25349, n_21836, n_21837);
  not g46803 (n_21838, n25348);
  not g46804 (n_21839, n25349);
  and g46805 (n25350, n_21838, n_21839);
  not g46806 (n_21840, n25343);
  not g46807 (n_21841, n25350);
  and g46808 (n25351, n_21840, n_21841);
  not g46809 (n_21842, n25351);
  and g46810 (n25352, n_21840, n_21842);
  and g46811 (n25353, n_21841, n_21842);
  not g46812 (n_21843, n25352);
  not g46813 (n_21844, n25353);
  and g46814 (n25354, n_21843, n_21844);
  and g46815 (n25355, \b[44] , n12668);
  and g46816 (n25356, \b[42] , n13047);
  and g46817 (n25357, \b[43] , n12663);
  and g46823 (n25360, n7072, n12671);
  not g46826 (n_21849, n25361);
  and g46827 (n25362, \a[62] , n_21849);
  not g46828 (n_21850, n25362);
  and g46829 (n25363, \a[62] , n_21850);
  and g46830 (n25364, n_21849, n_21850);
  not g46831 (n_21851, n25363);
  not g46832 (n_21852, n25364);
  and g46833 (n25365, n_21851, n_21852);
  not g46834 (n_21853, n25354);
  and g46835 (n25366, n_21853, n25365);
  not g46836 (n_21854, n25365);
  and g46837 (n25367, n25354, n_21854);
  not g46838 (n_21855, n25366);
  not g46839 (n_21856, n25367);
  and g46840 (n25368, n_21855, n_21856);
  and g46841 (n25369, \b[47] , n11531);
  and g46842 (n25370, \b[45] , n11896);
  and g46843 (n25371, \b[46] , n11526);
  and g46849 (n25374, n7703, n11534);
  not g46852 (n_21861, n25375);
  and g46853 (n25376, \a[59] , n_21861);
  not g46854 (n_21862, n25376);
  and g46855 (n25377, \a[59] , n_21862);
  and g46856 (n25378, n_21861, n_21862);
  not g46857 (n_21863, n25377);
  not g46858 (n_21864, n25378);
  and g46859 (n25379, n_21863, n_21864);
  not g46860 (n_21865, n25368);
  not g46861 (n_21866, n25379);
  and g46862 (n25380, n_21865, n_21866);
  and g46863 (n25381, n25368, n25379);
  not g46864 (n_21867, n25380);
  not g46865 (n_21868, n25381);
  and g46866 (n25382, n_21867, n_21868);
  not g46867 (n_21869, n25382);
  and g46868 (n25383, n25342, n_21869);
  not g46869 (n_21870, n25342);
  and g46870 (n25384, n_21870, n25382);
  not g46871 (n_21871, n25383);
  not g46872 (n_21872, n25384);
  and g46873 (n25385, n_21871, n_21872);
  and g46874 (n25386, \b[50] , n10426);
  and g46875 (n25387, \b[48] , n10796);
  and g46876 (n25388, \b[49] , n10421);
  and g46882 (n25391, n8949, n10429);
  not g46885 (n_21877, n25392);
  and g46886 (n25393, \a[56] , n_21877);
  not g46887 (n_21878, n25393);
  and g46888 (n25394, \a[56] , n_21878);
  and g46889 (n25395, n_21877, n_21878);
  not g46890 (n_21879, n25394);
  not g46891 (n_21880, n25395);
  and g46892 (n25396, n_21879, n_21880);
  not g46893 (n_21881, n25385);
  and g46894 (n25397, n_21881, n25396);
  not g46895 (n_21882, n25396);
  and g46896 (n25398, n25385, n_21882);
  not g46897 (n_21883, n25397);
  not g46898 (n_21884, n25398);
  and g46899 (n25399, n_21883, n_21884);
  not g46900 (n_21885, n25341);
  and g46901 (n25400, n_21885, n25399);
  not g46902 (n_21886, n25400);
  and g46903 (n25401, n_21885, n_21886);
  and g46904 (n25402, n25399, n_21886);
  not g46905 (n_21887, n25401);
  not g46906 (n_21888, n25402);
  and g46907 (n25403, n_21887, n_21888);
  not g46908 (n_21889, n25340);
  not g46909 (n_21890, n25403);
  and g46910 (n25404, n_21889, n_21890);
  and g46911 (n25405, n25340, n_21888);
  and g46912 (n25406, n_21887, n25405);
  not g46913 (n_21891, n25404);
  not g46914 (n_21892, n25406);
  and g46915 (n25407, n_21891, n_21892);
  not g46916 (n_21893, n25329);
  and g46917 (n25408, n_21893, n25407);
  not g46918 (n_21894, n25408);
  and g46919 (n25409, n_21893, n_21894);
  and g46920 (n25410, n25407, n_21894);
  not g46921 (n_21895, n25409);
  not g46922 (n_21896, n25410);
  and g46923 (n25411, n_21895, n_21896);
  not g46924 (n_21897, n25328);
  not g46925 (n_21898, n25411);
  and g46926 (n25412, n_21897, n_21898);
  and g46927 (n25413, n25328, n_21896);
  and g46928 (n25414, n_21895, n25413);
  not g46929 (n_21899, n25412);
  not g46930 (n_21900, n25414);
  and g46931 (n25415, n_21899, n_21900);
  not g46932 (n_21901, n25317);
  and g46933 (n25416, n_21901, n25415);
  not g46934 (n_21902, n25415);
  and g46935 (n25417, n25317, n_21902);
  not g46936 (n_21903, n25416);
  not g46937 (n_21904, n25417);
  and g46938 (n25418, n_21903, n_21904);
  not g46939 (n_21905, n25316);
  and g46940 (n25419, n_21905, n25418);
  not g46941 (n_21906, n25419);
  and g46942 (n25420, n25418, n_21906);
  and g46943 (n25421, n_21905, n_21906);
  not g46944 (n_21907, n25420);
  not g46945 (n_21908, n25421);
  and g46946 (n25422, n_21907, n_21908);
  and g46947 (n25423, n_21759, n_21769);
  and g46948 (n25424, n25422, n25423);
  not g46949 (n_21909, n25422);
  not g46950 (n_21910, n25423);
  and g46951 (n25425, n_21909, n_21910);
  not g46952 (n_21911, n25424);
  not g46953 (n_21912, n25425);
  and g46954 (n25426, n_21911, n_21912);
  and g46955 (n25427, \b[62] , n6595);
  and g46956 (n25428, \b[60] , n6902);
  and g46957 (n25429, \b[61] , n6590);
  and g46963 (n25432, n6598, n13370);
  not g46966 (n_21917, n25433);
  and g46967 (n25434, \a[44] , n_21917);
  not g46968 (n_21918, n25434);
  and g46969 (n25435, \a[44] , n_21918);
  and g46970 (n25436, n_21917, n_21918);
  not g46971 (n_21919, n25435);
  not g46972 (n_21920, n25436);
  and g46973 (n25437, n_21919, n_21920);
  not g46974 (n_21921, n25437);
  and g46975 (n25438, n25426, n_21921);
  not g46976 (n_21922, n25438);
  and g46977 (n25439, n25426, n_21922);
  and g46978 (n25440, n_21921, n_21922);
  not g46979 (n_21923, n25439);
  not g46980 (n_21924, n25440);
  and g46981 (n25441, n_21923, n_21924);
  not g46982 (n_21925, n25305);
  and g46983 (n25442, n_21925, n25441);
  not g46984 (n_21926, n25441);
  and g46985 (n25443, n25305, n_21926);
  not g46986 (n_21927, n25442);
  not g46987 (n_21928, n25443);
  and g46988 (n25444, n_21927, n_21928);
  not g46989 (n_21929, n25293);
  not g46990 (n_21930, n25444);
  and g46991 (n25445, n_21929, n_21930);
  and g46992 (n25446, n25293, n25444);
  not g46993 (n_21931, n25445);
  not g46994 (n_21932, n25446);
  and g46995 (n25447, n_21931, n_21932);
  not g46996 (n_21933, n25292);
  and g46997 (n25448, n_21933, n25447);
  not g46998 (n_21934, n25447);
  and g46999 (n25449, n25292, n_21934);
  not g47000 (n_21935, n25448);
  not g47001 (n_21936, n25449);
  and g47002 (\f[104] , n_21935, n_21936);
  and g47003 (n25451, n_21931, n_21935);
  and g47004 (n25452, \b[60] , n7446);
  and g47005 (n25453, \b[58] , n7787);
  and g47006 (n25454, \b[59] , n7441);
  and g47012 (n25457, n7449, n12211);
  not g47015 (n_21941, n25458);
  and g47016 (n25459, \a[47] , n_21941);
  not g47017 (n_21942, n25459);
  and g47018 (n25460, \a[47] , n_21942);
  and g47019 (n25461, n_21941, n_21942);
  not g47020 (n_21943, n25460);
  not g47021 (n_21944, n25461);
  and g47022 (n25462, n_21943, n_21944);
  and g47023 (n25463, n_21894, n_21899);
  and g47024 (n25464, \b[57] , n8362);
  and g47025 (n25465, \b[55] , n8715);
  and g47026 (n25466, \b[56] , n8357);
  and g47032 (n25469, n8365, n11410);
  not g47035 (n_21949, n25470);
  and g47036 (n25471, \a[50] , n_21949);
  not g47037 (n_21950, n25471);
  and g47038 (n25472, \a[50] , n_21950);
  and g47039 (n25473, n_21949, n_21950);
  not g47040 (n_21951, n25472);
  not g47041 (n_21952, n25473);
  and g47042 (n25474, n_21951, n_21952);
  and g47043 (n25475, n_21886, n_21891);
  and g47044 (n25476, n_21872, n_21884);
  and g47045 (n25477, \b[51] , n10426);
  and g47046 (n25478, \b[49] , n10796);
  and g47047 (n25479, \b[50] , n10421);
  and g47053 (n25482, n8976, n10429);
  not g47056 (n_21957, n25483);
  and g47057 (n25484, \a[56] , n_21957);
  not g47058 (n_21958, n25484);
  and g47059 (n25485, \a[56] , n_21958);
  and g47060 (n25486, n_21957, n_21958);
  not g47061 (n_21959, n25485);
  not g47062 (n_21960, n25486);
  and g47063 (n25487, n_21959, n_21960);
  and g47064 (n25488, \a[41] , n_21674);
  and g47065 (n25489, n_4853, n25146);
  not g47066 (n_21961, n25488);
  not g47067 (n_21962, n25489);
  and g47068 (n25490, n_21961, n_21962);
  and g47069 (n25491, \b[41] , n13903);
  and g47070 (n25492, \b[42] , n_11555);
  not g47071 (n_21963, n25491);
  not g47072 (n_21964, n25492);
  and g47073 (n25493, n_21963, n_21964);
  and g47074 (n25494, n25490, n25493);
  not g47075 (n_21965, n25490);
  not g47076 (n_21966, n25493);
  and g47077 (n25495, n_21965, n_21966);
  not g47078 (n_21967, n25494);
  not g47079 (n_21968, n25495);
  and g47080 (n25496, n_21967, n_21968);
  and g47081 (n25497, \b[45] , n12668);
  and g47082 (n25498, \b[43] , n13047);
  and g47083 (n25499, \b[44] , n12663);
  and g47089 (n25502, n7361, n12671);
  not g47092 (n_21973, n25503);
  and g47093 (n25504, \a[62] , n_21973);
  not g47094 (n_21974, n25504);
  and g47095 (n25505, \a[62] , n_21974);
  and g47096 (n25506, n_21973, n_21974);
  not g47097 (n_21975, n25505);
  not g47098 (n_21976, n25506);
  and g47099 (n25507, n_21975, n_21976);
  not g47100 (n_21977, n25507);
  and g47101 (n25508, n25496, n_21977);
  not g47102 (n_21978, n25508);
  and g47103 (n25509, n25496, n_21978);
  and g47104 (n25510, n_21977, n_21978);
  not g47105 (n_21979, n25509);
  not g47106 (n_21980, n25510);
  and g47107 (n25511, n_21979, n_21980);
  and g47108 (n25512, n_21837, n_21842);
  and g47109 (n25513, n25511, n25512);
  not g47110 (n_21981, n25511);
  not g47111 (n_21982, n25512);
  and g47112 (n25514, n_21981, n_21982);
  not g47113 (n_21983, n25513);
  not g47114 (n_21984, n25514);
  and g47115 (n25515, n_21983, n_21984);
  and g47116 (n25516, \b[48] , n11531);
  and g47117 (n25517, \b[46] , n11896);
  and g47118 (n25518, \b[47] , n11526);
  and g47124 (n25521, n8009, n11534);
  not g47127 (n_21989, n25522);
  and g47128 (n25523, \a[59] , n_21989);
  not g47129 (n_21990, n25523);
  and g47130 (n25524, \a[59] , n_21990);
  and g47131 (n25525, n_21989, n_21990);
  not g47132 (n_21991, n25524);
  not g47133 (n_21992, n25525);
  and g47134 (n25526, n_21991, n_21992);
  not g47135 (n_21993, n25526);
  and g47136 (n25527, n25515, n_21993);
  not g47137 (n_21994, n25527);
  and g47138 (n25528, n25515, n_21994);
  and g47139 (n25529, n_21993, n_21994);
  not g47140 (n_21995, n25528);
  not g47141 (n_21996, n25529);
  and g47142 (n25530, n_21995, n_21996);
  and g47143 (n25531, n_21853, n_21854);
  not g47144 (n_21997, n25531);
  and g47145 (n25532, n_21867, n_21997);
  not g47146 (n_21998, n25530);
  not g47147 (n_21999, n25532);
  and g47148 (n25533, n_21998, n_21999);
  and g47149 (n25534, n25530, n25532);
  not g47150 (n_22000, n25533);
  not g47151 (n_22001, n25534);
  and g47152 (n25535, n_22000, n_22001);
  not g47153 (n_22002, n25487);
  and g47154 (n25536, n_22002, n25535);
  not g47155 (n_22003, n25536);
  and g47156 (n25537, n_22002, n_22003);
  and g47157 (n25538, n25535, n_22003);
  not g47158 (n_22004, n25537);
  not g47159 (n_22005, n25538);
  and g47160 (n25539, n_22004, n_22005);
  not g47161 (n_22006, n25476);
  not g47162 (n_22007, n25539);
  and g47163 (n25540, n_22006, n_22007);
  not g47164 (n_22008, n25540);
  and g47165 (n25541, n_22006, n_22008);
  and g47166 (n25542, n_22007, n_22008);
  not g47167 (n_22009, n25541);
  not g47168 (n_22010, n25542);
  and g47169 (n25543, n_22009, n_22010);
  and g47170 (n25544, \b[54] , n9339);
  and g47171 (n25545, \b[52] , n9732);
  and g47172 (n25546, \b[53] , n9334);
  and g47178 (n25549, n9342, n9998);
  not g47181 (n_22015, n25550);
  and g47182 (n25551, \a[53] , n_22015);
  not g47183 (n_22016, n25551);
  and g47184 (n25552, \a[53] , n_22016);
  and g47185 (n25553, n_22015, n_22016);
  not g47186 (n_22017, n25552);
  not g47187 (n_22018, n25553);
  and g47188 (n25554, n_22017, n_22018);
  and g47189 (n25555, n25543, n25554);
  not g47190 (n_22019, n25543);
  not g47191 (n_22020, n25554);
  and g47192 (n25556, n_22019, n_22020);
  not g47193 (n_22021, n25555);
  not g47194 (n_22022, n25556);
  and g47195 (n25557, n_22021, n_22022);
  not g47196 (n_22023, n25475);
  and g47197 (n25558, n_22023, n25557);
  not g47198 (n_22024, n25557);
  and g47199 (n25559, n25475, n_22024);
  not g47200 (n_22025, n25558);
  not g47201 (n_22026, n25559);
  and g47202 (n25560, n_22025, n_22026);
  not g47203 (n_22027, n25560);
  and g47204 (n25561, n25474, n_22027);
  not g47205 (n_22028, n25474);
  and g47206 (n25562, n_22028, n25560);
  not g47207 (n_22029, n25561);
  not g47208 (n_22030, n25562);
  and g47209 (n25563, n_22029, n_22030);
  not g47210 (n_22031, n25463);
  and g47211 (n25564, n_22031, n25563);
  not g47212 (n_22032, n25563);
  and g47213 (n25565, n25463, n_22032);
  not g47214 (n_22033, n25564);
  not g47215 (n_22034, n25565);
  and g47216 (n25566, n_22033, n_22034);
  not g47217 (n_22035, n25462);
  and g47218 (n25567, n_22035, n25566);
  not g47219 (n_22036, n25567);
  and g47220 (n25568, n25566, n_22036);
  and g47221 (n25569, n_22035, n_22036);
  not g47222 (n_22037, n25568);
  not g47223 (n_22038, n25569);
  and g47224 (n25570, n_22037, n_22038);
  and g47225 (n25571, n_21903, n_21906);
  and g47226 (n25572, n25570, n25571);
  not g47227 (n_22039, n25570);
  not g47228 (n_22040, n25571);
  and g47229 (n25573, n_22039, n_22040);
  not g47230 (n_22041, n25572);
  not g47231 (n_22042, n25573);
  and g47232 (n25574, n_22041, n_22042);
  and g47233 (n25575, \b[63] , n6595);
  and g47234 (n25576, \b[61] , n6902);
  and g47235 (n25577, \b[62] , n6590);
  and g47241 (n25580, n6598, n13771);
  not g47244 (n_22047, n25581);
  and g47245 (n25582, \a[44] , n_22047);
  not g47246 (n_22048, n25582);
  and g47247 (n25583, \a[44] , n_22048);
  and g47248 (n25584, n_22047, n_22048);
  not g47249 (n_22049, n25583);
  not g47250 (n_22050, n25584);
  and g47251 (n25585, n_22049, n_22050);
  not g47252 (n_22051, n25585);
  and g47253 (n25586, n25574, n_22051);
  not g47254 (n_22052, n25586);
  and g47255 (n25587, n25574, n_22052);
  and g47256 (n25588, n_22051, n_22052);
  not g47257 (n_22053, n25587);
  not g47258 (n_22054, n25588);
  and g47259 (n25589, n_22053, n_22054);
  and g47260 (n25590, n_21912, n_21922);
  and g47261 (n25591, n25589, n25590);
  not g47262 (n_22055, n25589);
  not g47263 (n_22056, n25590);
  and g47264 (n25592, n_22055, n_22056);
  not g47265 (n_22057, n25591);
  not g47266 (n_22058, n25592);
  and g47267 (n25593, n_22057, n_22058);
  and g47268 (n25594, n_21925, n_21926);
  not g47269 (n_22059, n25594);
  and g47270 (n25595, n_21807, n_22059);
  not g47271 (n_22060, n25595);
  and g47272 (n25596, n25593, n_22060);
  not g47273 (n_22061, n25593);
  and g47274 (n25597, n_22061, n25595);
  not g47275 (n_22062, n25596);
  not g47276 (n_22063, n25597);
  and g47277 (n25598, n_22062, n_22063);
  not g47278 (n_22064, n25451);
  and g47279 (n25599, n_22064, n25598);
  not g47280 (n_22065, n25598);
  and g47281 (n25600, n25451, n_22065);
  not g47282 (n_22066, n25599);
  not g47283 (n_22067, n25600);
  and g47284 (\f[105] , n_22066, n_22067);
  and g47285 (n25602, n_22036, n_22042);
  and g47286 (n25603, \b[62] , n6902);
  and g47287 (n25604, \b[63] , n6590);
  not g47288 (n_22068, n25603);
  not g47289 (n_22069, n25604);
  and g47290 (n25605, n_22068, n_22069);
  not g47291 (n_22070, n6598);
  and g47292 (n25606, n_22070, n25605);
  and g47293 (n25607, n13800, n25605);
  not g47294 (n_22071, n25606);
  not g47295 (n_22072, n25607);
  and g47296 (n25608, n_22071, n_22072);
  not g47297 (n_22073, n25608);
  and g47298 (n25609, \a[44] , n_22073);
  and g47299 (n25610, n_5572, n25608);
  not g47300 (n_22074, n25609);
  not g47301 (n_22075, n25610);
  and g47302 (n25611, n_22074, n_22075);
  not g47303 (n_22076, n25602);
  not g47304 (n_22077, n25611);
  and g47305 (n25612, n_22076, n_22077);
  and g47306 (n25613, n25602, n25611);
  not g47307 (n_22078, n25612);
  not g47308 (n_22079, n25613);
  and g47309 (n25614, n_22078, n_22079);
  and g47310 (n25615, \b[61] , n7446);
  and g47311 (n25616, \b[59] , n7787);
  and g47312 (n25617, \b[60] , n7441);
  and g47318 (n25620, n7449, n12969);
  not g47321 (n_22084, n25621);
  and g47322 (n25622, \a[47] , n_22084);
  not g47323 (n_22085, n25622);
  and g47324 (n25623, \a[47] , n_22085);
  and g47325 (n25624, n_22084, n_22085);
  not g47326 (n_22086, n25623);
  not g47327 (n_22087, n25624);
  and g47328 (n25625, n_22086, n_22087);
  and g47329 (n25626, n_22030, n_22033);
  and g47330 (n25627, n_22022, n_22025);
  and g47331 (n25628, n_21978, n_21984);
  and g47332 (n25629, \b[42] , n13903);
  and g47333 (n25630, \b[43] , n_11555);
  not g47334 (n_22088, n25629);
  not g47335 (n_22089, n25630);
  and g47336 (n25631, n_22088, n_22089);
  and g47337 (n25632, n_4853, n_21674);
  not g47338 (n_22090, n25632);
  and g47339 (n25633, n_21968, n_22090);
  not g47340 (n_22091, n25633);
  and g47341 (n25634, n25631, n_22091);
  not g47342 (n_22092, n25634);
  and g47343 (n25635, n25631, n_22092);
  and g47344 (n25636, n_22091, n_22092);
  not g47345 (n_22093, n25635);
  not g47346 (n_22094, n25636);
  and g47347 (n25637, n_22093, n_22094);
  and g47348 (n25638, \b[46] , n12668);
  and g47349 (n25639, \b[44] , n13047);
  and g47350 (n25640, \b[45] , n12663);
  not g47351 (n_22095, n25639);
  not g47352 (n_22096, n25640);
  and g47353 (n25641, n_22095, n_22096);
  not g47354 (n_22097, n25638);
  and g47355 (n25642, n_22097, n25641);
  and g47356 (n25643, n_12644, n25642);
  and g47357 (n25644, n_13970, n25642);
  not g47358 (n_22098, n25643);
  not g47359 (n_22099, n25644);
  and g47360 (n25645, n_22098, n_22099);
  not g47361 (n_22100, n25645);
  and g47362 (n25646, \a[62] , n_22100);
  and g47363 (n25647, n_10843, n25645);
  not g47364 (n_22101, n25646);
  not g47365 (n_22102, n25647);
  and g47366 (n25648, n_22101, n_22102);
  not g47367 (n_22103, n25637);
  not g47368 (n_22104, n25648);
  and g47369 (n25649, n_22103, n_22104);
  and g47370 (n25650, n25637, n25648);
  not g47371 (n_22105, n25649);
  not g47372 (n_22106, n25650);
  and g47373 (n25651, n_22105, n_22106);
  not g47374 (n_22107, n25628);
  and g47375 (n25652, n_22107, n25651);
  not g47376 (n_22108, n25651);
  and g47377 (n25653, n25628, n_22108);
  not g47378 (n_22109, n25652);
  not g47379 (n_22110, n25653);
  and g47380 (n25654, n_22109, n_22110);
  and g47381 (n25655, \b[49] , n11531);
  and g47382 (n25656, \b[47] , n11896);
  and g47383 (n25657, \b[48] , n11526);
  and g47389 (n25660, n8625, n11534);
  not g47392 (n_22115, n25661);
  and g47393 (n25662, \a[59] , n_22115);
  not g47394 (n_22116, n25662);
  and g47395 (n25663, \a[59] , n_22116);
  and g47396 (n25664, n_22115, n_22116);
  not g47397 (n_22117, n25663);
  not g47398 (n_22118, n25664);
  and g47399 (n25665, n_22117, n_22118);
  not g47400 (n_22119, n25665);
  and g47401 (n25666, n25654, n_22119);
  not g47402 (n_22120, n25666);
  and g47403 (n25667, n25654, n_22120);
  and g47404 (n25668, n_22119, n_22120);
  not g47405 (n_22121, n25667);
  not g47406 (n_22122, n25668);
  and g47407 (n25669, n_22121, n_22122);
  and g47408 (n25670, n_21994, n_22000);
  and g47409 (n25671, n25669, n25670);
  not g47410 (n_22123, n25669);
  not g47411 (n_22124, n25670);
  and g47412 (n25672, n_22123, n_22124);
  not g47413 (n_22125, n25671);
  not g47414 (n_22126, n25672);
  and g47415 (n25673, n_22125, n_22126);
  and g47416 (n25674, \b[52] , n10426);
  and g47417 (n25675, \b[50] , n10796);
  and g47418 (n25676, \b[51] , n10421);
  and g47424 (n25679, n9628, n10429);
  not g47427 (n_22131, n25680);
  and g47428 (n25681, \a[56] , n_22131);
  not g47429 (n_22132, n25681);
  and g47430 (n25682, \a[56] , n_22132);
  and g47431 (n25683, n_22131, n_22132);
  not g47432 (n_22133, n25682);
  not g47433 (n_22134, n25683);
  and g47434 (n25684, n_22133, n_22134);
  not g47435 (n_22135, n25684);
  and g47436 (n25685, n25673, n_22135);
  not g47437 (n_22136, n25685);
  and g47438 (n25686, n25673, n_22136);
  and g47439 (n25687, n_22135, n_22136);
  not g47440 (n_22137, n25686);
  not g47441 (n_22138, n25687);
  and g47442 (n25688, n_22137, n_22138);
  and g47443 (n25689, n_22003, n_22008);
  and g47444 (n25690, n25688, n25689);
  not g47445 (n_22139, n25688);
  not g47446 (n_22140, n25689);
  and g47447 (n25691, n_22139, n_22140);
  not g47448 (n_22141, n25690);
  not g47449 (n_22142, n25691);
  and g47450 (n25692, n_22141, n_22142);
  and g47451 (n25693, \b[55] , n9339);
  and g47452 (n25694, \b[53] , n9732);
  and g47453 (n25695, \b[54] , n9334);
  and g47459 (n25698, n9342, n10684);
  not g47462 (n_22147, n25699);
  and g47463 (n25700, \a[53] , n_22147);
  not g47464 (n_22148, n25700);
  and g47465 (n25701, \a[53] , n_22148);
  and g47466 (n25702, n_22147, n_22148);
  not g47467 (n_22149, n25701);
  not g47468 (n_22150, n25702);
  and g47469 (n25703, n_22149, n_22150);
  not g47470 (n_22151, n25703);
  and g47471 (n25704, n25692, n_22151);
  not g47472 (n_22152, n25704);
  and g47473 (n25705, n25692, n_22152);
  and g47474 (n25706, n_22151, n_22152);
  not g47475 (n_22153, n25705);
  not g47476 (n_22154, n25706);
  and g47477 (n25707, n_22153, n_22154);
  not g47478 (n_22155, n25627);
  and g47479 (n25708, n_22155, n25707);
  not g47480 (n_22156, n25707);
  and g47481 (n25709, n25627, n_22156);
  not g47482 (n_22157, n25708);
  not g47483 (n_22158, n25709);
  and g47484 (n25710, n_22157, n_22158);
  and g47485 (n25711, \b[58] , n8362);
  and g47486 (n25712, \b[56] , n8715);
  and g47487 (n25713, \b[57] , n8357);
  and g47493 (n25716, n8365, n11436);
  not g47496 (n_22163, n25717);
  and g47497 (n25718, \a[50] , n_22163);
  not g47498 (n_22164, n25718);
  and g47499 (n25719, \a[50] , n_22164);
  and g47500 (n25720, n_22163, n_22164);
  not g47501 (n_22165, n25719);
  not g47502 (n_22166, n25720);
  and g47503 (n25721, n_22165, n_22166);
  and g47504 (n25722, n25710, n25721);
  not g47505 (n_22167, n25710);
  not g47506 (n_22168, n25721);
  and g47507 (n25723, n_22167, n_22168);
  not g47508 (n_22169, n25722);
  not g47509 (n_22170, n25723);
  and g47510 (n25724, n_22169, n_22170);
  not g47511 (n_22171, n25626);
  and g47512 (n25725, n_22171, n25724);
  not g47513 (n_22172, n25725);
  and g47514 (n25726, n_22171, n_22172);
  and g47515 (n25727, n25724, n_22172);
  not g47516 (n_22173, n25726);
  not g47517 (n_22174, n25727);
  and g47518 (n25728, n_22173, n_22174);
  not g47519 (n_22175, n25625);
  not g47520 (n_22176, n25728);
  and g47521 (n25729, n_22175, n_22176);
  not g47522 (n_22177, n25729);
  and g47523 (n25730, n_22175, n_22177);
  and g47524 (n25731, n_22176, n_22177);
  not g47525 (n_22178, n25730);
  not g47526 (n_22179, n25731);
  and g47527 (n25732, n_22178, n_22179);
  not g47528 (n_22180, n25732);
  and g47529 (n25733, n25614, n_22180);
  not g47530 (n_22181, n25733);
  and g47531 (n25734, n25614, n_22181);
  and g47532 (n25735, n_22180, n_22181);
  not g47533 (n_22182, n25734);
  not g47534 (n_22183, n25735);
  and g47535 (n25736, n_22182, n_22183);
  and g47536 (n25737, n_22052, n_22058);
  and g47537 (n25738, n25736, n25737);
  not g47538 (n_22184, n25736);
  not g47539 (n_22185, n25737);
  and g47540 (n25739, n_22184, n_22185);
  not g47541 (n_22186, n25738);
  not g47542 (n_22187, n25739);
  and g47543 (n25740, n_22186, n_22187);
  and g47544 (n25741, n_22062, n_22066);
  not g47545 (n_22188, n25741);
  and g47546 (n25742, n25740, n_22188);
  not g47547 (n_22189, n25740);
  and g47548 (n25743, n_22189, n25741);
  not g47549 (n_22190, n25742);
  not g47550 (n_22191, n25743);
  and g47551 (\f[106] , n_22190, n_22191);
  and g47552 (n25745, n_22187, n_22190);
  and g47553 (n25746, n_22078, n_22181);
  and g47554 (n25747, n_22172, n_22177);
  and g47555 (n25748, \b[63] , n6902);
  and g47556 (n25749, n6598, n13797);
  not g47557 (n_22192, n25748);
  not g47558 (n_22193, n25749);
  and g47559 (n25750, n_22192, n_22193);
  not g47560 (n_22194, n25750);
  and g47561 (n25751, \a[44] , n_22194);
  not g47562 (n_22195, n25751);
  and g47563 (n25752, \a[44] , n_22195);
  and g47564 (n25753, n_22194, n_22195);
  not g47565 (n_22196, n25752);
  not g47566 (n_22197, n25753);
  and g47567 (n25754, n_22196, n_22197);
  not g47568 (n_22198, n25747);
  not g47569 (n_22199, n25754);
  and g47570 (n25755, n_22198, n_22199);
  not g47571 (n_22200, n25755);
  and g47572 (n25756, n_22198, n_22200);
  and g47573 (n25757, n_22199, n_22200);
  not g47574 (n_22201, n25756);
  not g47575 (n_22202, n25757);
  and g47576 (n25758, n_22201, n_22202);
  and g47577 (n25759, \b[59] , n8362);
  and g47578 (n25760, \b[57] , n8715);
  and g47579 (n25761, \b[58] , n8357);
  and g47585 (n25764, n8365, n12179);
  not g47588 (n_22207, n25765);
  and g47589 (n25766, \a[50] , n_22207);
  not g47590 (n_22208, n25766);
  and g47591 (n25767, \a[50] , n_22208);
  and g47592 (n25768, n_22207, n_22208);
  not g47593 (n_22209, n25767);
  not g47594 (n_22210, n25768);
  and g47595 (n25769, n_22209, n_22210);
  and g47596 (n25770, n_22142, n_22152);
  and g47597 (n25771, \b[56] , n9339);
  and g47598 (n25772, \b[54] , n9732);
  and g47599 (n25773, \b[55] , n9334);
  and g47605 (n25776, n9342, n10708);
  not g47608 (n_22215, n25777);
  and g47609 (n25778, \a[53] , n_22215);
  not g47610 (n_22216, n25778);
  and g47611 (n25779, \a[53] , n_22216);
  and g47612 (n25780, n_22215, n_22216);
  not g47613 (n_22217, n25779);
  not g47614 (n_22218, n25780);
  and g47615 (n25781, n_22217, n_22218);
  and g47616 (n25782, n_22126, n_22136);
  and g47617 (n25783, \b[53] , n10426);
  and g47618 (n25784, \b[51] , n10796);
  and g47619 (n25785, \b[52] , n10421);
  and g47625 (n25788, n9972, n10429);
  not g47628 (n_22223, n25789);
  and g47629 (n25790, \a[56] , n_22223);
  not g47630 (n_22224, n25790);
  and g47631 (n25791, \a[56] , n_22224);
  and g47632 (n25792, n_22223, n_22224);
  not g47633 (n_22225, n25791);
  not g47634 (n_22226, n25792);
  and g47635 (n25793, n_22225, n_22226);
  and g47636 (n25794, n_22109, n_22120);
  and g47637 (n25795, \b[50] , n11531);
  and g47638 (n25796, \b[48] , n11896);
  and g47639 (n25797, \b[49] , n11526);
  and g47645 (n25800, n8949, n11534);
  not g47648 (n_22231, n25801);
  and g47649 (n25802, \a[59] , n_22231);
  not g47650 (n_22232, n25802);
  and g47651 (n25803, \a[59] , n_22232);
  and g47652 (n25804, n_22231, n_22232);
  not g47653 (n_22233, n25803);
  not g47654 (n_22234, n25804);
  and g47655 (n25805, n_22233, n_22234);
  and g47656 (n25806, n_22092, n_22105);
  and g47657 (n25807, \b[43] , n13903);
  and g47658 (n25808, \b[44] , n_11555);
  not g47659 (n_22235, n25807);
  not g47660 (n_22236, n25808);
  and g47661 (n25809, n_22235, n_22236);
  not g47662 (n_22237, n25809);
  and g47663 (n25810, n25631, n_22237);
  not g47664 (n_22238, n25631);
  and g47665 (n25811, n_22238, n25809);
  not g47666 (n_22239, n25810);
  not g47667 (n_22240, n25811);
  and g47668 (n25812, n_22239, n_22240);
  and g47669 (n25813, \b[47] , n12668);
  and g47670 (n25814, \b[45] , n13047);
  and g47671 (n25815, \b[46] , n12663);
  not g47672 (n_22241, n25814);
  not g47673 (n_22242, n25815);
  and g47674 (n25816, n_22241, n_22242);
  not g47675 (n_22243, n25813);
  and g47676 (n25817, n_22243, n25816);
  and g47677 (n25818, n_12644, n25817);
  and g47678 (n25819, n_16121, n25817);
  not g47679 (n_22244, n25818);
  not g47680 (n_22245, n25819);
  and g47681 (n25820, n_22244, n_22245);
  not g47682 (n_22246, n25820);
  and g47683 (n25821, \a[62] , n_22246);
  and g47684 (n25822, n_10843, n25820);
  not g47685 (n_22247, n25821);
  not g47686 (n_22248, n25822);
  and g47687 (n25823, n_22247, n_22248);
  not g47688 (n_22249, n25823);
  and g47689 (n25824, n25812, n_22249);
  not g47690 (n_22250, n25812);
  and g47691 (n25825, n_22250, n25823);
  not g47692 (n_22251, n25824);
  not g47693 (n_22252, n25825);
  and g47694 (n25826, n_22251, n_22252);
  not g47695 (n_22253, n25806);
  and g47696 (n25827, n_22253, n25826);
  not g47697 (n_22254, n25827);
  and g47698 (n25828, n_22253, n_22254);
  and g47699 (n25829, n25826, n_22254);
  not g47700 (n_22255, n25828);
  not g47701 (n_22256, n25829);
  and g47702 (n25830, n_22255, n_22256);
  not g47703 (n_22257, n25805);
  not g47704 (n_22258, n25830);
  and g47705 (n25831, n_22257, n_22258);
  and g47706 (n25832, n25805, n_22256);
  and g47707 (n25833, n_22255, n25832);
  not g47708 (n_22259, n25831);
  not g47709 (n_22260, n25833);
  and g47710 (n25834, n_22259, n_22260);
  not g47711 (n_22261, n25794);
  and g47712 (n25835, n_22261, n25834);
  not g47713 (n_22262, n25835);
  and g47714 (n25836, n_22261, n_22262);
  and g47715 (n25837, n25834, n_22262);
  not g47716 (n_22263, n25836);
  not g47717 (n_22264, n25837);
  and g47718 (n25838, n_22263, n_22264);
  not g47719 (n_22265, n25793);
  not g47720 (n_22266, n25838);
  and g47721 (n25839, n_22265, n_22266);
  and g47722 (n25840, n25793, n_22264);
  and g47723 (n25841, n_22263, n25840);
  not g47724 (n_22267, n25839);
  not g47725 (n_22268, n25841);
  and g47726 (n25842, n_22267, n_22268);
  not g47727 (n_22269, n25782);
  and g47728 (n25843, n_22269, n25842);
  not g47729 (n_22270, n25843);
  and g47730 (n25844, n_22269, n_22270);
  and g47731 (n25845, n25842, n_22270);
  not g47732 (n_22271, n25844);
  not g47733 (n_22272, n25845);
  and g47734 (n25846, n_22271, n_22272);
  not g47735 (n_22273, n25781);
  not g47736 (n_22274, n25846);
  and g47737 (n25847, n_22273, n_22274);
  and g47738 (n25848, n25781, n_22272);
  and g47739 (n25849, n_22271, n25848);
  not g47740 (n_22275, n25847);
  not g47741 (n_22276, n25849);
  and g47742 (n25850, n_22275, n_22276);
  not g47743 (n_22277, n25770);
  and g47744 (n25851, n_22277, n25850);
  not g47745 (n_22278, n25850);
  and g47746 (n25852, n25770, n_22278);
  not g47747 (n_22279, n25851);
  not g47748 (n_22280, n25852);
  and g47749 (n25853, n_22279, n_22280);
  not g47750 (n_22281, n25769);
  and g47751 (n25854, n_22281, n25853);
  not g47752 (n_22282, n25854);
  and g47753 (n25855, n25853, n_22282);
  and g47754 (n25856, n_22281, n_22282);
  not g47755 (n_22283, n25855);
  not g47756 (n_22284, n25856);
  and g47757 (n25857, n_22283, n_22284);
  and g47758 (n25858, n_22155, n_22156);
  not g47759 (n_22285, n25858);
  and g47760 (n25859, n_22170, n_22285);
  not g47761 (n_22286, n25857);
  not g47762 (n_22287, n25859);
  and g47763 (n25860, n_22286, n_22287);
  not g47764 (n_22288, n25860);
  and g47765 (n25861, n_22286, n_22288);
  and g47766 (n25862, n_22287, n_22288);
  not g47767 (n_22289, n25861);
  not g47768 (n_22290, n25862);
  and g47769 (n25863, n_22289, n_22290);
  and g47770 (n25864, \b[62] , n7446);
  and g47771 (n25865, \b[60] , n7787);
  and g47772 (n25866, \b[61] , n7441);
  and g47778 (n25869, n7449, n13370);
  not g47781 (n_22295, n25870);
  and g47782 (n25871, \a[47] , n_22295);
  not g47783 (n_22296, n25871);
  and g47784 (n25872, \a[47] , n_22296);
  and g47785 (n25873, n_22295, n_22296);
  not g47786 (n_22297, n25872);
  not g47787 (n_22298, n25873);
  and g47788 (n25874, n_22297, n_22298);
  not g47789 (n_22299, n25863);
  not g47790 (n_22300, n25874);
  and g47791 (n25875, n_22299, n_22300);
  not g47792 (n_22301, n25875);
  and g47793 (n25876, n_22299, n_22301);
  and g47794 (n25877, n_22300, n_22301);
  not g47795 (n_22302, n25876);
  not g47796 (n_22303, n25877);
  and g47797 (n25878, n_22302, n_22303);
  not g47798 (n_22304, n25758);
  and g47799 (n25879, n_22304, n25878);
  not g47800 (n_22305, n25878);
  and g47801 (n25880, n25758, n_22305);
  not g47802 (n_22306, n25879);
  not g47803 (n_22307, n25880);
  and g47804 (n25881, n_22306, n_22307);
  not g47805 (n_22308, n25746);
  not g47806 (n_22309, n25881);
  and g47807 (n25882, n_22308, n_22309);
  and g47808 (n25883, n25746, n25881);
  not g47809 (n_22310, n25882);
  not g47810 (n_22311, n25883);
  and g47811 (n25884, n_22310, n_22311);
  not g47812 (n_22312, n25745);
  and g47813 (n25885, n_22312, n25884);
  not g47814 (n_22313, n25884);
  and g47815 (n25886, n25745, n_22313);
  not g47816 (n_22314, n25885);
  not g47817 (n_22315, n25886);
  and g47818 (\f[107] , n_22314, n_22315);
  and g47819 (n25888, n_22310, n_22314);
  and g47820 (n25889, \b[63] , n7446);
  and g47821 (n25890, \b[61] , n7787);
  and g47822 (n25891, \b[62] , n7441);
  and g47828 (n25894, n7449, n13771);
  not g47831 (n_22320, n25895);
  and g47832 (n25896, \a[47] , n_22320);
  not g47833 (n_22321, n25896);
  and g47834 (n25897, \a[47] , n_22321);
  and g47835 (n25898, n_22320, n_22321);
  not g47836 (n_22322, n25897);
  not g47837 (n_22323, n25898);
  and g47838 (n25899, n_22322, n_22323);
  and g47839 (n25900, n_22279, n_22282);
  and g47840 (n25901, \b[60] , n8362);
  and g47841 (n25902, \b[58] , n8715);
  and g47842 (n25903, \b[59] , n8357);
  and g47848 (n25906, n8365, n12211);
  not g47851 (n_22328, n25907);
  and g47852 (n25908, \a[50] , n_22328);
  not g47853 (n_22329, n25908);
  and g47854 (n25909, \a[50] , n_22329);
  and g47855 (n25910, n_22328, n_22329);
  not g47856 (n_22330, n25909);
  not g47857 (n_22331, n25910);
  and g47858 (n25911, n_22330, n_22331);
  and g47859 (n25912, n_22270, n_22275);
  and g47860 (n25913, \b[57] , n9339);
  and g47861 (n25914, \b[55] , n9732);
  and g47862 (n25915, \b[56] , n9334);
  and g47868 (n25918, n9342, n11410);
  not g47871 (n_22336, n25919);
  and g47872 (n25920, \a[53] , n_22336);
  not g47873 (n_22337, n25920);
  and g47874 (n25921, \a[53] , n_22337);
  and g47875 (n25922, n_22336, n_22337);
  not g47876 (n_22338, n25921);
  not g47877 (n_22339, n25922);
  and g47878 (n25923, n_22338, n_22339);
  and g47879 (n25924, n_22262, n_22267);
  and g47880 (n25925, \b[54] , n10426);
  and g47881 (n25926, \b[52] , n10796);
  and g47882 (n25927, \b[53] , n10421);
  and g47888 (n25930, n9998, n10429);
  not g47891 (n_22344, n25931);
  and g47892 (n25932, \a[56] , n_22344);
  not g47893 (n_22345, n25932);
  and g47894 (n25933, \a[56] , n_22345);
  and g47895 (n25934, n_22344, n_22345);
  not g47896 (n_22346, n25933);
  not g47897 (n_22347, n25934);
  and g47898 (n25935, n_22346, n_22347);
  and g47899 (n25936, n_22254, n_22259);
  and g47900 (n25937, n_22239, n_22251);
  and g47901 (n25938, \b[44] , n13903);
  and g47902 (n25939, \b[45] , n_11555);
  not g47903 (n_22348, n25938);
  not g47904 (n_22349, n25939);
  and g47905 (n25940, n_22348, n_22349);
  not g47906 (n_22350, n25940);
  and g47907 (n25941, n_5572, n_22350);
  and g47908 (n25942, \a[44] , n25940);
  not g47909 (n_22351, n25941);
  not g47910 (n_22352, n25942);
  and g47911 (n25943, n_22351, n_22352);
  and g47912 (n25944, n_22238, n25943);
  not g47913 (n_22353, n25944);
  and g47914 (n25945, n_22238, n_22353);
  and g47915 (n25946, n25943, n_22353);
  not g47916 (n_22354, n25945);
  not g47917 (n_22355, n25946);
  and g47918 (n25947, n_22354, n_22355);
  not g47919 (n_22356, n25937);
  not g47920 (n_22357, n25947);
  and g47921 (n25948, n_22356, n_22357);
  not g47922 (n_22358, n25948);
  and g47923 (n25949, n_22356, n_22358);
  and g47924 (n25950, n_22357, n_22358);
  not g47925 (n_22359, n25949);
  not g47926 (n_22360, n25950);
  and g47927 (n25951, n_22359, n_22360);
  and g47928 (n25952, \b[48] , n12668);
  and g47929 (n25953, \b[46] , n13047);
  and g47930 (n25954, \b[47] , n12663);
  and g47936 (n25957, n8009, n12671);
  not g47939 (n_22365, n25958);
  and g47940 (n25959, \a[62] , n_22365);
  not g47941 (n_22366, n25959);
  and g47942 (n25960, \a[62] , n_22366);
  and g47943 (n25961, n_22365, n_22366);
  not g47944 (n_22367, n25960);
  not g47945 (n_22368, n25961);
  and g47946 (n25962, n_22367, n_22368);
  not g47947 (n_22369, n25951);
  not g47948 (n_22370, n25962);
  and g47949 (n25963, n_22369, n_22370);
  not g47950 (n_22371, n25963);
  and g47951 (n25964, n_22369, n_22371);
  and g47952 (n25965, n_22370, n_22371);
  not g47953 (n_22372, n25964);
  not g47954 (n_22373, n25965);
  and g47955 (n25966, n_22372, n_22373);
  and g47956 (n25967, \b[51] , n11531);
  and g47957 (n25968, \b[49] , n11896);
  and g47958 (n25969, \b[50] , n11526);
  and g47964 (n25972, n8976, n11534);
  not g47967 (n_22378, n25973);
  and g47968 (n25974, \a[59] , n_22378);
  not g47969 (n_22379, n25974);
  and g47970 (n25975, \a[59] , n_22379);
  and g47971 (n25976, n_22378, n_22379);
  not g47972 (n_22380, n25975);
  not g47973 (n_22381, n25976);
  and g47974 (n25977, n_22380, n_22381);
  and g47975 (n25978, n25966, n25977);
  not g47976 (n_22382, n25966);
  not g47977 (n_22383, n25977);
  and g47978 (n25979, n_22382, n_22383);
  not g47979 (n_22384, n25978);
  not g47980 (n_22385, n25979);
  and g47981 (n25980, n_22384, n_22385);
  not g47982 (n_22386, n25936);
  and g47983 (n25981, n_22386, n25980);
  not g47984 (n_22387, n25980);
  and g47985 (n25982, n25936, n_22387);
  not g47986 (n_22388, n25981);
  not g47987 (n_22389, n25982);
  and g47988 (n25983, n_22388, n_22389);
  not g47989 (n_22390, n25983);
  and g47990 (n25984, n25935, n_22390);
  not g47991 (n_22391, n25935);
  and g47992 (n25985, n_22391, n25983);
  not g47993 (n_22392, n25984);
  not g47994 (n_22393, n25985);
  and g47995 (n25986, n_22392, n_22393);
  not g47996 (n_22394, n25924);
  and g47997 (n25987, n_22394, n25986);
  not g47998 (n_22395, n25986);
  and g47999 (n25988, n25924, n_22395);
  not g48000 (n_22396, n25987);
  not g48001 (n_22397, n25988);
  and g48002 (n25989, n_22396, n_22397);
  not g48003 (n_22398, n25989);
  and g48004 (n25990, n25923, n_22398);
  not g48005 (n_22399, n25923);
  and g48006 (n25991, n_22399, n25989);
  not g48007 (n_22400, n25990);
  not g48008 (n_22401, n25991);
  and g48009 (n25992, n_22400, n_22401);
  not g48010 (n_22402, n25912);
  and g48011 (n25993, n_22402, n25992);
  not g48012 (n_22403, n25992);
  and g48013 (n25994, n25912, n_22403);
  not g48014 (n_22404, n25993);
  not g48015 (n_22405, n25994);
  and g48016 (n25995, n_22404, n_22405);
  not g48017 (n_22406, n25995);
  and g48018 (n25996, n25911, n_22406);
  not g48019 (n_22407, n25911);
  and g48020 (n25997, n_22407, n25995);
  not g48021 (n_22408, n25996);
  not g48022 (n_22409, n25997);
  and g48023 (n25998, n_22408, n_22409);
  not g48024 (n_22410, n25900);
  and g48025 (n25999, n_22410, n25998);
  not g48026 (n_22411, n25998);
  and g48027 (n26000, n25900, n_22411);
  not g48028 (n_22412, n25999);
  not g48029 (n_22413, n26000);
  and g48030 (n26001, n_22412, n_22413);
  not g48031 (n_22414, n25899);
  and g48032 (n26002, n_22414, n26001);
  not g48033 (n_22415, n26002);
  and g48034 (n26003, n26001, n_22415);
  and g48035 (n26004, n_22414, n_22415);
  not g48036 (n_22416, n26003);
  not g48037 (n_22417, n26004);
  and g48038 (n26005, n_22416, n_22417);
  and g48039 (n26006, n_22288, n_22301);
  and g48040 (n26007, n26005, n26006);
  not g48041 (n_22418, n26005);
  not g48042 (n_22419, n26006);
  and g48043 (n26008, n_22418, n_22419);
  not g48044 (n_22420, n26007);
  not g48045 (n_22421, n26008);
  and g48046 (n26009, n_22420, n_22421);
  and g48047 (n26010, n_22304, n_22305);
  not g48048 (n_22422, n26010);
  and g48049 (n26011, n_22200, n_22422);
  not g48050 (n_22423, n26011);
  and g48051 (n26012, n26009, n_22423);
  not g48052 (n_22424, n26009);
  and g48053 (n26013, n_22424, n26011);
  not g48054 (n_22425, n26012);
  not g48055 (n_22426, n26013);
  and g48056 (n26014, n_22425, n_22426);
  not g48057 (n_22427, n25888);
  and g48058 (n26015, n_22427, n26014);
  not g48059 (n_22428, n26014);
  and g48060 (n26016, n25888, n_22428);
  not g48061 (n_22429, n26015);
  not g48062 (n_22430, n26016);
  and g48063 (\f[108] , n_22429, n_22430);
  and g48064 (n26018, n_22409, n_22412);
  and g48065 (n26019, \b[62] , n7787);
  and g48066 (n26020, \b[63] , n7441);
  not g48067 (n_22431, n26019);
  not g48068 (n_22432, n26020);
  and g48069 (n26021, n_22431, n_22432);
  not g48070 (n_22433, n7449);
  and g48071 (n26022, n_22433, n26021);
  and g48072 (n26023, n13800, n26021);
  not g48073 (n_22434, n26022);
  not g48074 (n_22435, n26023);
  and g48075 (n26024, n_22434, n_22435);
  not g48076 (n_22436, n26024);
  and g48077 (n26025, \a[47] , n_22436);
  and g48078 (n26026, n_6314, n26024);
  not g48079 (n_22437, n26025);
  not g48080 (n_22438, n26026);
  and g48081 (n26027, n_22437, n_22438);
  not g48082 (n_22439, n26018);
  not g48083 (n_22440, n26027);
  and g48084 (n26028, n_22439, n_22440);
  and g48085 (n26029, n26018, n26027);
  not g48086 (n_22441, n26028);
  not g48087 (n_22442, n26029);
  and g48088 (n26030, n_22441, n_22442);
  and g48089 (n26031, \b[61] , n8362);
  and g48090 (n26032, \b[59] , n8715);
  and g48091 (n26033, \b[60] , n8357);
  and g48097 (n26036, n8365, n12969);
  not g48100 (n_22447, n26037);
  and g48101 (n26038, \a[50] , n_22447);
  not g48102 (n_22448, n26038);
  and g48103 (n26039, \a[50] , n_22448);
  and g48104 (n26040, n_22447, n_22448);
  not g48105 (n_22449, n26039);
  not g48106 (n_22450, n26040);
  and g48107 (n26041, n_22449, n_22450);
  and g48108 (n26042, n_22401, n_22404);
  and g48109 (n26043, n_22393, n_22396);
  and g48110 (n26044, \b[55] , n10426);
  and g48111 (n26045, \b[53] , n10796);
  and g48112 (n26046, \b[54] , n10421);
  and g48118 (n26049, n10429, n10684);
  not g48121 (n_22455, n26050);
  and g48122 (n26051, \a[56] , n_22455);
  not g48123 (n_22456, n26051);
  and g48124 (n26052, \a[56] , n_22456);
  and g48125 (n26053, n_22455, n_22456);
  not g48126 (n_22457, n26052);
  not g48127 (n_22458, n26053);
  and g48128 (n26054, n_22457, n_22458);
  and g48129 (n26055, n_22385, n_22388);
  and g48130 (n26056, \b[52] , n11531);
  and g48131 (n26057, \b[50] , n11896);
  and g48132 (n26058, \b[51] , n11526);
  and g48138 (n26061, n9628, n11534);
  not g48141 (n_22463, n26062);
  and g48142 (n26063, \a[59] , n_22463);
  not g48143 (n_22464, n26063);
  and g48144 (n26064, \a[59] , n_22464);
  and g48145 (n26065, n_22463, n_22464);
  not g48146 (n_22465, n26064);
  not g48147 (n_22466, n26065);
  and g48148 (n26066, n_22465, n_22466);
  and g48149 (n26067, n_22358, n_22371);
  and g48150 (n26068, \b[45] , n13903);
  and g48151 (n26069, \b[46] , n_11555);
  not g48152 (n_22467, n26068);
  not g48153 (n_22468, n26069);
  and g48154 (n26070, n_22467, n_22468);
  and g48155 (n26071, n_22351, n_22353);
  not g48156 (n_22469, n26070);
  and g48157 (n26072, n_22469, n26071);
  not g48158 (n_22470, n26071);
  and g48159 (n26073, n26070, n_22470);
  not g48160 (n_22471, n26072);
  not g48161 (n_22472, n26073);
  and g48162 (n26074, n_22471, n_22472);
  and g48163 (n26075, \b[49] , n12668);
  and g48164 (n26076, \b[47] , n13047);
  and g48165 (n26077, \b[48] , n12663);
  and g48171 (n26080, n8625, n12671);
  not g48174 (n_22477, n26081);
  and g48175 (n26082, \a[62] , n_22477);
  not g48176 (n_22478, n26082);
  and g48177 (n26083, \a[62] , n_22478);
  and g48178 (n26084, n_22477, n_22478);
  not g48179 (n_22479, n26083);
  not g48180 (n_22480, n26084);
  and g48181 (n26085, n_22479, n_22480);
  not g48182 (n_22481, n26074);
  and g48183 (n26086, n_22481, n26085);
  not g48184 (n_22482, n26085);
  and g48185 (n26087, n26074, n_22482);
  not g48186 (n_22483, n26086);
  not g48187 (n_22484, n26087);
  and g48188 (n26088, n_22483, n_22484);
  not g48189 (n_22485, n26067);
  and g48190 (n26089, n_22485, n26088);
  not g48191 (n_22486, n26089);
  and g48192 (n26090, n_22485, n_22486);
  and g48193 (n26091, n26088, n_22486);
  not g48194 (n_22487, n26090);
  not g48195 (n_22488, n26091);
  and g48196 (n26092, n_22487, n_22488);
  not g48197 (n_22489, n26066);
  not g48198 (n_22490, n26092);
  and g48199 (n26093, n_22489, n_22490);
  and g48200 (n26094, n26066, n_22488);
  and g48201 (n26095, n_22487, n26094);
  not g48202 (n_22491, n26093);
  not g48203 (n_22492, n26095);
  and g48204 (n26096, n_22491, n_22492);
  not g48205 (n_22493, n26055);
  and g48206 (n26097, n_22493, n26096);
  not g48207 (n_22494, n26096);
  and g48208 (n26098, n26055, n_22494);
  not g48209 (n_22495, n26097);
  not g48210 (n_22496, n26098);
  and g48211 (n26099, n_22495, n_22496);
  not g48212 (n_22497, n26054);
  and g48213 (n26100, n_22497, n26099);
  not g48214 (n_22498, n26100);
  and g48215 (n26101, n26099, n_22498);
  and g48216 (n26102, n_22497, n_22498);
  not g48217 (n_22499, n26101);
  not g48218 (n_22500, n26102);
  and g48219 (n26103, n_22499, n_22500);
  not g48220 (n_22501, n26043);
  and g48221 (n26104, n_22501, n26103);
  not g48222 (n_22502, n26103);
  and g48223 (n26105, n26043, n_22502);
  not g48224 (n_22503, n26104);
  not g48225 (n_22504, n26105);
  and g48226 (n26106, n_22503, n_22504);
  and g48227 (n26107, \b[58] , n9339);
  and g48228 (n26108, \b[56] , n9732);
  and g48229 (n26109, \b[57] , n9334);
  and g48235 (n26112, n9342, n11436);
  not g48238 (n_22509, n26113);
  and g48239 (n26114, \a[53] , n_22509);
  not g48240 (n_22510, n26114);
  and g48241 (n26115, \a[53] , n_22510);
  and g48242 (n26116, n_22509, n_22510);
  not g48243 (n_22511, n26115);
  not g48244 (n_22512, n26116);
  and g48245 (n26117, n_22511, n_22512);
  and g48246 (n26118, n26106, n26117);
  not g48247 (n_22513, n26106);
  not g48248 (n_22514, n26117);
  and g48249 (n26119, n_22513, n_22514);
  not g48250 (n_22515, n26118);
  not g48251 (n_22516, n26119);
  and g48252 (n26120, n_22515, n_22516);
  not g48253 (n_22517, n26042);
  and g48254 (n26121, n_22517, n26120);
  not g48255 (n_22518, n26121);
  and g48256 (n26122, n_22517, n_22518);
  and g48257 (n26123, n26120, n_22518);
  not g48258 (n_22519, n26122);
  not g48259 (n_22520, n26123);
  and g48260 (n26124, n_22519, n_22520);
  not g48261 (n_22521, n26041);
  not g48262 (n_22522, n26124);
  and g48263 (n26125, n_22521, n_22522);
  not g48264 (n_22523, n26125);
  and g48265 (n26126, n_22521, n_22523);
  and g48266 (n26127, n_22522, n_22523);
  not g48267 (n_22524, n26126);
  not g48268 (n_22525, n26127);
  and g48269 (n26128, n_22524, n_22525);
  not g48270 (n_22526, n26128);
  and g48271 (n26129, n26030, n_22526);
  not g48272 (n_22527, n26129);
  and g48273 (n26130, n26030, n_22527);
  and g48274 (n26131, n_22526, n_22527);
  not g48275 (n_22528, n26130);
  not g48276 (n_22529, n26131);
  and g48277 (n26132, n_22528, n_22529);
  and g48278 (n26133, n_22415, n_22421);
  and g48279 (n26134, n26132, n26133);
  not g48280 (n_22530, n26132);
  not g48281 (n_22531, n26133);
  and g48282 (n26135, n_22530, n_22531);
  not g48283 (n_22532, n26134);
  not g48284 (n_22533, n26135);
  and g48285 (n26136, n_22532, n_22533);
  and g48286 (n26137, n_22425, n_22429);
  not g48287 (n_22534, n26137);
  and g48288 (n26138, n26136, n_22534);
  not g48289 (n_22535, n26136);
  and g48290 (n26139, n_22535, n26137);
  not g48291 (n_22536, n26138);
  not g48292 (n_22537, n26139);
  and g48293 (\f[109] , n_22536, n_22537);
  and g48294 (n26141, \b[59] , n9339);
  and g48295 (n26142, \b[57] , n9732);
  and g48296 (n26143, \b[58] , n9334);
  and g48302 (n26146, n9342, n12179);
  not g48305 (n_22542, n26147);
  and g48306 (n26148, \a[53] , n_22542);
  not g48307 (n_22543, n26148);
  and g48308 (n26149, \a[53] , n_22543);
  and g48309 (n26150, n_22542, n_22543);
  not g48310 (n_22544, n26149);
  not g48311 (n_22545, n26150);
  and g48312 (n26151, n_22544, n_22545);
  and g48313 (n26152, n_22495, n_22498);
  and g48314 (n26153, \b[56] , n10426);
  and g48315 (n26154, \b[54] , n10796);
  and g48316 (n26155, \b[55] , n10421);
  and g48322 (n26158, n10429, n10708);
  not g48325 (n_22550, n26159);
  and g48326 (n26160, \a[56] , n_22550);
  not g48327 (n_22551, n26160);
  and g48328 (n26161, \a[56] , n_22551);
  and g48329 (n26162, n_22550, n_22551);
  not g48330 (n_22552, n26161);
  not g48331 (n_22553, n26162);
  and g48332 (n26163, n_22552, n_22553);
  and g48333 (n26164, n_22486, n_22491);
  and g48334 (n26165, \b[53] , n11531);
  and g48335 (n26166, \b[51] , n11896);
  and g48336 (n26167, \b[52] , n11526);
  and g48342 (n26170, n9972, n11534);
  not g48345 (n_22558, n26171);
  and g48346 (n26172, \a[59] , n_22558);
  not g48347 (n_22559, n26172);
  and g48348 (n26173, \a[59] , n_22559);
  and g48349 (n26174, n_22558, n_22559);
  not g48350 (n_22560, n26173);
  not g48351 (n_22561, n26174);
  and g48352 (n26175, n_22560, n_22561);
  and g48353 (n26176, n_22472, n_22484);
  and g48354 (n26177, \b[46] , n13903);
  and g48355 (n26178, \b[47] , n_11555);
  not g48356 (n_22562, n26177);
  not g48357 (n_22563, n26178);
  and g48358 (n26179, n_22562, n_22563);
  not g48359 (n_22564, n26179);
  and g48360 (n26180, n26070, n_22564);
  and g48361 (n26181, n_22469, n26179);
  not g48362 (n_22565, n26176);
  not g48363 (n_22566, n26181);
  and g48364 (n26182, n_22565, n_22566);
  not g48365 (n_22567, n26180);
  and g48366 (n26183, n_22567, n26182);
  not g48367 (n_22568, n26183);
  and g48368 (n26184, n_22565, n_22568);
  and g48369 (n26185, n_22566, n_22568);
  and g48370 (n26186, n_22567, n26185);
  not g48371 (n_22569, n26184);
  not g48372 (n_22570, n26186);
  and g48373 (n26187, n_22569, n_22570);
  and g48374 (n26188, \b[50] , n12668);
  and g48375 (n26189, \b[48] , n13047);
  and g48376 (n26190, \b[49] , n12663);
  and g48382 (n26193, n8949, n12671);
  not g48385 (n_22575, n26194);
  and g48386 (n26195, \a[62] , n_22575);
  not g48387 (n_22576, n26195);
  and g48388 (n26196, \a[62] , n_22576);
  and g48389 (n26197, n_22575, n_22576);
  not g48390 (n_22577, n26196);
  not g48391 (n_22578, n26197);
  and g48392 (n26198, n_22577, n_22578);
  not g48393 (n_22579, n26187);
  and g48394 (n26199, n_22579, n26198);
  not g48395 (n_22580, n26198);
  and g48396 (n26200, n26187, n_22580);
  not g48397 (n_22581, n26199);
  not g48398 (n_22582, n26200);
  and g48399 (n26201, n_22581, n_22582);
  not g48400 (n_22583, n26175);
  not g48401 (n_22584, n26201);
  and g48402 (n26202, n_22583, n_22584);
  and g48403 (n26203, n26175, n26201);
  not g48404 (n_22585, n26202);
  not g48405 (n_22586, n26203);
  and g48406 (n26204, n_22585, n_22586);
  not g48407 (n_22587, n26164);
  and g48408 (n26205, n_22587, n26204);
  not g48409 (n_22588, n26205);
  and g48410 (n26206, n_22587, n_22588);
  and g48411 (n26207, n26204, n_22588);
  not g48412 (n_22589, n26206);
  not g48413 (n_22590, n26207);
  and g48414 (n26208, n_22589, n_22590);
  not g48415 (n_22591, n26163);
  not g48416 (n_22592, n26208);
  and g48417 (n26209, n_22591, n_22592);
  and g48418 (n26210, n26163, n_22590);
  and g48419 (n26211, n_22589, n26210);
  not g48420 (n_22593, n26209);
  not g48421 (n_22594, n26211);
  and g48422 (n26212, n_22593, n_22594);
  not g48423 (n_22595, n26152);
  and g48424 (n26213, n_22595, n26212);
  not g48425 (n_22596, n26212);
  and g48426 (n26214, n26152, n_22596);
  not g48427 (n_22597, n26213);
  not g48428 (n_22598, n26214);
  and g48429 (n26215, n_22597, n_22598);
  not g48430 (n_22599, n26151);
  and g48431 (n26216, n_22599, n26215);
  not g48432 (n_22600, n26216);
  and g48433 (n26217, n26215, n_22600);
  and g48434 (n26218, n_22599, n_22600);
  not g48435 (n_22601, n26217);
  not g48436 (n_22602, n26218);
  and g48437 (n26219, n_22601, n_22602);
  and g48438 (n26220, n_22501, n_22502);
  not g48439 (n_22603, n26220);
  and g48440 (n26221, n_22516, n_22603);
  not g48441 (n_22604, n26219);
  not g48442 (n_22605, n26221);
  and g48443 (n26222, n_22604, n_22605);
  not g48444 (n_22606, n26222);
  and g48445 (n26223, n_22604, n_22606);
  and g48446 (n26224, n_22605, n_22606);
  not g48447 (n_22607, n26223);
  not g48448 (n_22608, n26224);
  and g48449 (n26225, n_22607, n_22608);
  and g48450 (n26226, \b[62] , n8362);
  and g48451 (n26227, \b[60] , n8715);
  and g48452 (n26228, \b[61] , n8357);
  and g48458 (n26231, n8365, n13370);
  not g48461 (n_22613, n26232);
  and g48462 (n26233, \a[50] , n_22613);
  not g48463 (n_22614, n26233);
  and g48464 (n26234, \a[50] , n_22614);
  and g48465 (n26235, n_22613, n_22614);
  not g48466 (n_22615, n26234);
  not g48467 (n_22616, n26235);
  and g48468 (n26236, n_22615, n_22616);
  not g48469 (n_22617, n26225);
  not g48470 (n_22618, n26236);
  and g48471 (n26237, n_22617, n_22618);
  not g48472 (n_22619, n26237);
  and g48473 (n26238, n_22617, n_22619);
  and g48474 (n26239, n_22618, n_22619);
  not g48475 (n_22620, n26238);
  not g48476 (n_22621, n26239);
  and g48477 (n26240, n_22620, n_22621);
  and g48478 (n26241, n_22518, n_22523);
  and g48479 (n26242, \b[63] , n7787);
  not g48480 (n_22622, n26242);
  and g48481 (n26243, n_22433, n_22622);
  and g48482 (n26244, n_11840, n_22622);
  not g48483 (n_22623, n26243);
  not g48484 (n_22624, n26244);
  and g48485 (n26245, n_22623, n_22624);
  not g48486 (n_22625, n26245);
  and g48487 (n26246, \a[47] , n_22625);
  and g48488 (n26247, n_6314, n26245);
  not g48489 (n_22626, n26246);
  not g48490 (n_22627, n26247);
  and g48491 (n26248, n_22626, n_22627);
  not g48492 (n_22628, n26241);
  not g48493 (n_22629, n26248);
  and g48494 (n26249, n_22628, n_22629);
  and g48495 (n26250, n26241, n26248);
  not g48496 (n_22630, n26249);
  not g48497 (n_22631, n26250);
  and g48498 (n26251, n_22630, n_22631);
  not g48499 (n_22632, n26240);
  and g48500 (n26252, n_22632, n26251);
  not g48501 (n_22633, n26252);
  and g48502 (n26253, n_22632, n_22633);
  and g48503 (n26254, n26251, n_22633);
  not g48504 (n_22634, n26253);
  not g48505 (n_22635, n26254);
  and g48506 (n26255, n_22634, n_22635);
  and g48507 (n26256, n_22441, n_22527);
  and g48508 (n26257, n26255, n26256);
  not g48509 (n_22636, n26255);
  not g48510 (n_22637, n26256);
  and g48511 (n26258, n_22636, n_22637);
  not g48512 (n_22638, n26257);
  not g48513 (n_22639, n26258);
  and g48514 (n26259, n_22638, n_22639);
  and g48515 (n26260, n_22533, n_22536);
  not g48516 (n_22640, n26260);
  and g48517 (n26261, n26259, n_22640);
  not g48518 (n_22641, n26259);
  and g48519 (n26262, n_22641, n26260);
  not g48520 (n_22642, n26261);
  not g48521 (n_22643, n26262);
  and g48522 (\f[110] , n_22642, n_22643);
  and g48523 (n26264, \b[63] , n8362);
  and g48524 (n26265, \b[61] , n8715);
  and g48525 (n26266, \b[62] , n8357);
  and g48531 (n26269, n8365, n13771);
  not g48534 (n_22648, n26270);
  and g48535 (n26271, \a[50] , n_22648);
  not g48536 (n_22649, n26271);
  and g48537 (n26272, \a[50] , n_22649);
  and g48538 (n26273, n_22648, n_22649);
  not g48539 (n_22650, n26272);
  not g48540 (n_22651, n26273);
  and g48541 (n26274, n_22650, n_22651);
  and g48542 (n26275, n_22597, n_22600);
  and g48543 (n26276, \b[60] , n9339);
  and g48544 (n26277, \b[58] , n9732);
  and g48545 (n26278, \b[59] , n9334);
  and g48551 (n26281, n9342, n12211);
  not g48554 (n_22656, n26282);
  and g48555 (n26283, \a[53] , n_22656);
  not g48556 (n_22657, n26283);
  and g48557 (n26284, \a[53] , n_22657);
  and g48558 (n26285, n_22656, n_22657);
  not g48559 (n_22658, n26284);
  not g48560 (n_22659, n26285);
  and g48561 (n26286, n_22658, n_22659);
  and g48562 (n26287, n_22588, n_22593);
  and g48563 (n26288, \b[57] , n10426);
  and g48564 (n26289, \b[55] , n10796);
  and g48565 (n26290, \b[56] , n10421);
  and g48571 (n26293, n10429, n11410);
  not g48574 (n_22664, n26294);
  and g48575 (n26295, \a[56] , n_22664);
  not g48576 (n_22665, n26295);
  and g48577 (n26296, \a[56] , n_22665);
  and g48578 (n26297, n_22664, n_22665);
  not g48579 (n_22666, n26296);
  not g48580 (n_22667, n26297);
  and g48581 (n26298, n_22666, n_22667);
  and g48582 (n26299, n_22579, n_22580);
  not g48583 (n_22668, n26299);
  and g48584 (n26300, n_22585, n_22668);
  and g48585 (n26301, \b[51] , n12668);
  and g48586 (n26302, \b[49] , n13047);
  and g48587 (n26303, \b[50] , n12663);
  and g48593 (n26306, n8976, n12671);
  not g48596 (n_22673, n26307);
  and g48597 (n26308, \a[62] , n_22673);
  not g48598 (n_22674, n26308);
  and g48599 (n26309, \a[62] , n_22674);
  and g48600 (n26310, n_22673, n_22674);
  not g48601 (n_22675, n26309);
  not g48602 (n_22676, n26310);
  and g48603 (n26311, n_22675, n_22676);
  and g48604 (n26312, \b[47] , n13903);
  and g48605 (n26313, \b[48] , n_11555);
  not g48606 (n_22677, n26312);
  not g48607 (n_22678, n26313);
  and g48608 (n26314, n_22677, n_22678);
  and g48609 (n26315, \a[47] , n_22564);
  and g48610 (n26316, n_6314, n26179);
  not g48611 (n_22679, n26315);
  not g48612 (n_22680, n26316);
  and g48613 (n26317, n_22679, n_22680);
  not g48614 (n_22681, n26314);
  not g48615 (n_22682, n26317);
  and g48616 (n26318, n_22681, n_22682);
  and g48617 (n26319, n26314, n26317);
  not g48618 (n_22683, n26318);
  not g48619 (n_22684, n26319);
  and g48620 (n26320, n_22683, n_22684);
  not g48621 (n_22685, n26311);
  and g48622 (n26321, n_22685, n26320);
  not g48623 (n_22686, n26321);
  and g48624 (n26322, n_22685, n_22686);
  and g48625 (n26323, n26320, n_22686);
  not g48626 (n_22687, n26322);
  not g48627 (n_22688, n26323);
  and g48628 (n26324, n_22687, n_22688);
  not g48629 (n_22689, n26185);
  not g48630 (n_22690, n26324);
  and g48631 (n26325, n_22689, n_22690);
  not g48632 (n_22691, n26325);
  and g48633 (n26326, n_22689, n_22691);
  and g48634 (n26327, n_22690, n_22691);
  not g48635 (n_22692, n26326);
  not g48636 (n_22693, n26327);
  and g48637 (n26328, n_22692, n_22693);
  and g48638 (n26329, \b[54] , n11531);
  and g48639 (n26330, \b[52] , n11896);
  and g48640 (n26331, \b[53] , n11526);
  and g48646 (n26334, n9998, n11534);
  not g48649 (n_22698, n26335);
  and g48650 (n26336, \a[59] , n_22698);
  not g48651 (n_22699, n26336);
  and g48652 (n26337, \a[59] , n_22699);
  and g48653 (n26338, n_22698, n_22699);
  not g48654 (n_22700, n26337);
  not g48655 (n_22701, n26338);
  and g48656 (n26339, n_22700, n_22701);
  and g48657 (n26340, n26328, n26339);
  not g48658 (n_22702, n26328);
  not g48659 (n_22703, n26339);
  and g48660 (n26341, n_22702, n_22703);
  not g48661 (n_22704, n26340);
  not g48662 (n_22705, n26341);
  and g48663 (n26342, n_22704, n_22705);
  not g48664 (n_22706, n26300);
  and g48665 (n26343, n_22706, n26342);
  not g48666 (n_22707, n26342);
  and g48667 (n26344, n26300, n_22707);
  not g48668 (n_22708, n26343);
  not g48669 (n_22709, n26344);
  and g48670 (n26345, n_22708, n_22709);
  not g48671 (n_22710, n26345);
  and g48672 (n26346, n26298, n_22710);
  not g48673 (n_22711, n26298);
  and g48674 (n26347, n_22711, n26345);
  not g48675 (n_22712, n26346);
  not g48676 (n_22713, n26347);
  and g48677 (n26348, n_22712, n_22713);
  not g48678 (n_22714, n26287);
  and g48679 (n26349, n_22714, n26348);
  not g48680 (n_22715, n26348);
  and g48681 (n26350, n26287, n_22715);
  not g48682 (n_22716, n26349);
  not g48683 (n_22717, n26350);
  and g48684 (n26351, n_22716, n_22717);
  not g48685 (n_22718, n26351);
  and g48686 (n26352, n26286, n_22718);
  not g48687 (n_22719, n26286);
  and g48688 (n26353, n_22719, n26351);
  not g48689 (n_22720, n26352);
  not g48690 (n_22721, n26353);
  and g48691 (n26354, n_22720, n_22721);
  not g48692 (n_22722, n26275);
  and g48693 (n26355, n_22722, n26354);
  not g48694 (n_22723, n26354);
  and g48695 (n26356, n26275, n_22723);
  not g48696 (n_22724, n26355);
  not g48697 (n_22725, n26356);
  and g48698 (n26357, n_22724, n_22725);
  not g48699 (n_22726, n26274);
  and g48700 (n26358, n_22726, n26357);
  not g48701 (n_22727, n26358);
  and g48702 (n26359, n26357, n_22727);
  and g48703 (n26360, n_22726, n_22727);
  not g48704 (n_22728, n26359);
  not g48705 (n_22729, n26360);
  and g48706 (n26361, n_22728, n_22729);
  and g48707 (n26362, n_22606, n_22619);
  and g48708 (n26363, n26361, n26362);
  not g48709 (n_22730, n26361);
  not g48710 (n_22731, n26362);
  and g48711 (n26364, n_22730, n_22731);
  not g48712 (n_22732, n26363);
  not g48713 (n_22733, n26364);
  and g48714 (n26365, n_22732, n_22733);
  and g48715 (n26366, n_22630, n_22633);
  not g48716 (n_22734, n26365);
  and g48717 (n26367, n_22734, n26366);
  not g48718 (n_22735, n26366);
  and g48719 (n26368, n26365, n_22735);
  not g48720 (n_22736, n26367);
  not g48721 (n_22737, n26368);
  and g48722 (n26369, n_22736, n_22737);
  and g48723 (n26370, n_22639, n_22642);
  not g48724 (n_22738, n26370);
  and g48725 (n26371, n26369, n_22738);
  not g48726 (n_22739, n26369);
  and g48727 (n26372, n_22739, n26370);
  not g48728 (n_22740, n26371);
  not g48729 (n_22741, n26372);
  and g48730 (\f[111] , n_22740, n_22741);
  and g48731 (n26374, \b[62] , n8715);
  and g48732 (n26375, \b[63] , n8357);
  not g48733 (n_22742, n26374);
  not g48734 (n_22743, n26375);
  and g48735 (n26376, n_22742, n_22743);
  and g48736 (n26377, n8365, n_11843);
  not g48737 (n_22744, n26377);
  and g48738 (n26378, n26376, n_22744);
  not g48739 (n_22745, n26378);
  and g48740 (n26379, \a[50] , n_22745);
  not g48741 (n_22746, n26379);
  and g48742 (n26380, \a[50] , n_22746);
  and g48743 (n26381, n_22745, n_22746);
  not g48744 (n_22747, n26380);
  not g48745 (n_22748, n26381);
  and g48746 (n26382, n_22747, n_22748);
  and g48747 (n26383, n_22721, n_22724);
  and g48748 (n26384, \b[61] , n9339);
  and g48749 (n26385, \b[59] , n9732);
  and g48750 (n26386, \b[60] , n9334);
  and g48756 (n26389, n9342, n12969);
  not g48759 (n_22753, n26390);
  and g48760 (n26391, \a[53] , n_22753);
  not g48761 (n_22754, n26391);
  and g48762 (n26392, \a[53] , n_22754);
  and g48763 (n26393, n_22753, n_22754);
  not g48764 (n_22755, n26392);
  not g48765 (n_22756, n26393);
  and g48766 (n26394, n_22755, n_22756);
  and g48767 (n26395, n_22713, n_22716);
  and g48768 (n26396, \b[58] , n10426);
  and g48769 (n26397, \b[56] , n10796);
  and g48770 (n26398, \b[57] , n10421);
  and g48776 (n26401, n10429, n11436);
  not g48779 (n_22761, n26402);
  and g48780 (n26403, \a[56] , n_22761);
  not g48781 (n_22762, n26403);
  and g48782 (n26404, \a[56] , n_22762);
  and g48783 (n26405, n_22761, n_22762);
  not g48784 (n_22763, n26404);
  not g48785 (n_22764, n26405);
  and g48786 (n26406, n_22763, n_22764);
  and g48787 (n26407, n_22705, n_22708);
  and g48788 (n26408, \b[55] , n11531);
  and g48789 (n26409, \b[53] , n11896);
  and g48790 (n26410, \b[54] , n11526);
  and g48796 (n26413, n10684, n11534);
  not g48799 (n_22769, n26414);
  and g48800 (n26415, \a[59] , n_22769);
  not g48801 (n_22770, n26415);
  and g48802 (n26416, \a[59] , n_22770);
  and g48803 (n26417, n_22769, n_22770);
  not g48804 (n_22771, n26416);
  not g48805 (n_22772, n26417);
  and g48806 (n26418, n_22771, n_22772);
  and g48807 (n26419, n_22686, n_22691);
  and g48808 (n26420, \b[48] , n13903);
  and g48809 (n26421, \b[49] , n_11555);
  not g48810 (n_22773, n26420);
  not g48811 (n_22774, n26421);
  and g48812 (n26422, n_22773, n_22774);
  and g48813 (n26423, n_6314, n_22564);
  not g48814 (n_22775, n26423);
  and g48815 (n26424, n_22683, n_22775);
  not g48816 (n_22776, n26424);
  and g48817 (n26425, n26422, n_22776);
  not g48818 (n_22777, n26422);
  and g48819 (n26426, n_22777, n26424);
  not g48820 (n_22778, n26425);
  not g48821 (n_22779, n26426);
  and g48822 (n26427, n_22778, n_22779);
  and g48823 (n26428, \b[52] , n12668);
  and g48824 (n26429, \b[50] , n13047);
  and g48825 (n26430, \b[51] , n12663);
  not g48826 (n_22780, n26429);
  not g48827 (n_22781, n26430);
  and g48828 (n26431, n_22780, n_22781);
  not g48829 (n_22782, n26428);
  and g48830 (n26432, n_22782, n26431);
  and g48831 (n26433, n_12644, n26432);
  and g48832 (n26434, n_16004, n26432);
  not g48833 (n_22783, n26433);
  not g48834 (n_22784, n26434);
  and g48835 (n26435, n_22783, n_22784);
  not g48836 (n_22785, n26435);
  and g48837 (n26436, \a[62] , n_22785);
  and g48838 (n26437, n_10843, n26435);
  not g48839 (n_22786, n26436);
  not g48840 (n_22787, n26437);
  and g48841 (n26438, n_22786, n_22787);
  not g48842 (n_22788, n26438);
  and g48843 (n26439, n26427, n_22788);
  not g48844 (n_22789, n26427);
  and g48845 (n26440, n_22789, n26438);
  not g48846 (n_22790, n26439);
  not g48847 (n_22791, n26440);
  and g48848 (n26441, n_22790, n_22791);
  not g48849 (n_22792, n26419);
  and g48850 (n26442, n_22792, n26441);
  not g48851 (n_22793, n26442);
  and g48852 (n26443, n_22792, n_22793);
  and g48853 (n26444, n26441, n_22793);
  not g48854 (n_22794, n26443);
  not g48855 (n_22795, n26444);
  and g48856 (n26445, n_22794, n_22795);
  not g48857 (n_22796, n26418);
  not g48858 (n_22797, n26445);
  and g48859 (n26446, n_22796, n_22797);
  and g48860 (n26447, n26418, n_22795);
  and g48861 (n26448, n_22794, n26447);
  not g48862 (n_22798, n26446);
  not g48863 (n_22799, n26448);
  and g48864 (n26449, n_22798, n_22799);
  not g48865 (n_22800, n26407);
  and g48866 (n26450, n_22800, n26449);
  not g48867 (n_22801, n26449);
  and g48868 (n26451, n26407, n_22801);
  not g48869 (n_22802, n26450);
  not g48870 (n_22803, n26451);
  and g48871 (n26452, n_22802, n_22803);
  not g48872 (n_22804, n26406);
  and g48873 (n26453, n_22804, n26452);
  not g48874 (n_22805, n26452);
  and g48875 (n26454, n26406, n_22805);
  not g48876 (n_22806, n26453);
  not g48877 (n_22807, n26454);
  and g48878 (n26455, n_22806, n_22807);
  not g48879 (n_22808, n26395);
  and g48880 (n26456, n_22808, n26455);
  not g48881 (n_22809, n26456);
  and g48882 (n26457, n_22808, n_22809);
  and g48883 (n26458, n26455, n_22809);
  not g48884 (n_22810, n26457);
  not g48885 (n_22811, n26458);
  and g48886 (n26459, n_22810, n_22811);
  not g48887 (n_22812, n26394);
  not g48888 (n_22813, n26459);
  and g48889 (n26460, n_22812, n_22813);
  and g48890 (n26461, n26394, n_22811);
  and g48891 (n26462, n_22810, n26461);
  not g48892 (n_22814, n26460);
  not g48893 (n_22815, n26462);
  and g48894 (n26463, n_22814, n_22815);
  not g48895 (n_22816, n26383);
  and g48896 (n26464, n_22816, n26463);
  not g48897 (n_22817, n26463);
  and g48898 (n26465, n26383, n_22817);
  not g48899 (n_22818, n26464);
  not g48900 (n_22819, n26465);
  and g48901 (n26466, n_22818, n_22819);
  not g48902 (n_22820, n26382);
  and g48903 (n26467, n_22820, n26466);
  not g48904 (n_22821, n26467);
  and g48905 (n26468, n26466, n_22821);
  and g48906 (n26469, n_22820, n_22821);
  not g48907 (n_22822, n26468);
  not g48908 (n_22823, n26469);
  and g48909 (n26470, n_22822, n_22823);
  and g48910 (n26471, n_22727, n_22733);
  and g48911 (n26472, n26470, n26471);
  not g48912 (n_22824, n26470);
  not g48913 (n_22825, n26471);
  and g48914 (n26473, n_22824, n_22825);
  not g48915 (n_22826, n26472);
  not g48916 (n_22827, n26473);
  and g48917 (n26474, n_22826, n_22827);
  and g48918 (n26475, n_22737, n_22740);
  not g48919 (n_22828, n26475);
  and g48920 (n26476, n26474, n_22828);
  not g48921 (n_22829, n26474);
  and g48922 (n26477, n_22829, n26475);
  not g48923 (n_22830, n26476);
  not g48924 (n_22831, n26477);
  and g48925 (\f[112] , n_22830, n_22831);
  and g48926 (n26479, \b[59] , n10426);
  and g48927 (n26480, \b[57] , n10796);
  and g48928 (n26481, \b[58] , n10421);
  and g48934 (n26484, n10429, n12179);
  not g48937 (n_22836, n26485);
  and g48938 (n26486, \a[56] , n_22836);
  not g48939 (n_22837, n26486);
  and g48940 (n26487, \a[56] , n_22837);
  and g48941 (n26488, n_22836, n_22837);
  not g48942 (n_22838, n26487);
  not g48943 (n_22839, n26488);
  and g48944 (n26489, n_22838, n_22839);
  and g48945 (n26490, n_22793, n_22798);
  and g48946 (n26491, \b[53] , n12668);
  and g48947 (n26492, \b[51] , n13047);
  and g48948 (n26493, \b[52] , n12663);
  and g48954 (n26496, n9972, n12671);
  not g48957 (n_22844, n26497);
  and g48958 (n26498, \a[62] , n_22844);
  not g48959 (n_22845, n26498);
  and g48960 (n26499, \a[62] , n_22845);
  and g48961 (n26500, n_22844, n_22845);
  not g48962 (n_22846, n26499);
  not g48963 (n_22847, n26500);
  and g48964 (n26501, n_22846, n_22847);
  and g48965 (n26502, \b[49] , n13903);
  and g48966 (n26503, \b[50] , n_11555);
  not g48967 (n_22848, n26502);
  not g48968 (n_22849, n26503);
  and g48969 (n26504, n_22848, n_22849);
  not g48970 (n_22850, n26504);
  and g48971 (n26505, n26422, n_22850);
  not g48972 (n_22851, n26505);
  and g48973 (n26506, n26422, n_22851);
  and g48974 (n26507, n_22850, n_22851);
  not g48975 (n_22852, n26506);
  not g48976 (n_22853, n26507);
  and g48977 (n26508, n_22852, n_22853);
  not g48978 (n_22854, n26501);
  not g48979 (n_22855, n26508);
  and g48980 (n26509, n_22854, n_22855);
  not g48981 (n_22856, n26509);
  and g48982 (n26510, n_22854, n_22856);
  and g48983 (n26511, n_22855, n_22856);
  not g48984 (n_22857, n26510);
  not g48985 (n_22858, n26511);
  and g48986 (n26512, n_22857, n_22858);
  and g48987 (n26513, n_22778, n_22790);
  and g48988 (n26514, n26512, n26513);
  not g48989 (n_22859, n26512);
  not g48990 (n_22860, n26513);
  and g48991 (n26515, n_22859, n_22860);
  not g48992 (n_22861, n26514);
  not g48993 (n_22862, n26515);
  and g48994 (n26516, n_22861, n_22862);
  and g48995 (n26517, \b[56] , n11531);
  and g48996 (n26518, \b[54] , n11896);
  and g48997 (n26519, \b[55] , n11526);
  and g49003 (n26522, n10708, n11534);
  not g49006 (n_22867, n26523);
  and g49007 (n26524, \a[59] , n_22867);
  not g49008 (n_22868, n26524);
  and g49009 (n26525, \a[59] , n_22868);
  and g49010 (n26526, n_22867, n_22868);
  not g49011 (n_22869, n26525);
  not g49012 (n_22870, n26526);
  and g49013 (n26527, n_22869, n_22870);
  not g49014 (n_22871, n26516);
  and g49015 (n26528, n_22871, n26527);
  not g49016 (n_22872, n26527);
  and g49017 (n26529, n26516, n_22872);
  not g49018 (n_22873, n26528);
  not g49019 (n_22874, n26529);
  and g49020 (n26530, n_22873, n_22874);
  not g49021 (n_22875, n26490);
  and g49022 (n26531, n_22875, n26530);
  not g49023 (n_22876, n26530);
  and g49024 (n26532, n26490, n_22876);
  not g49025 (n_22877, n26531);
  not g49026 (n_22878, n26532);
  and g49027 (n26533, n_22877, n_22878);
  not g49028 (n_22879, n26489);
  and g49029 (n26534, n_22879, n26533);
  not g49030 (n_22880, n26534);
  and g49031 (n26535, n26533, n_22880);
  and g49032 (n26536, n_22879, n_22880);
  not g49033 (n_22881, n26535);
  not g49034 (n_22882, n26536);
  and g49035 (n26537, n_22881, n_22882);
  and g49036 (n26538, n_22802, n_22806);
  and g49037 (n26539, n26537, n26538);
  not g49038 (n_22883, n26537);
  not g49039 (n_22884, n26538);
  and g49040 (n26540, n_22883, n_22884);
  not g49041 (n_22885, n26539);
  not g49042 (n_22886, n26540);
  and g49043 (n26541, n_22885, n_22886);
  and g49044 (n26542, \b[62] , n9339);
  and g49045 (n26543, \b[60] , n9732);
  and g49046 (n26544, \b[61] , n9334);
  and g49052 (n26547, n9342, n13370);
  not g49055 (n_22891, n26548);
  and g49056 (n26549, \a[53] , n_22891);
  not g49057 (n_22892, n26549);
  and g49058 (n26550, \a[53] , n_22892);
  and g49059 (n26551, n_22891, n_22892);
  not g49060 (n_22893, n26550);
  not g49061 (n_22894, n26551);
  and g49062 (n26552, n_22893, n_22894);
  not g49063 (n_22895, n26552);
  and g49064 (n26553, n26541, n_22895);
  not g49065 (n_22896, n26553);
  and g49066 (n26554, n26541, n_22896);
  and g49067 (n26555, n_22895, n_22896);
  not g49068 (n_22897, n26554);
  not g49069 (n_22898, n26555);
  and g49070 (n26556, n_22897, n_22898);
  and g49071 (n26557, n_22809, n_22814);
  and g49072 (n26558, \b[63] , n8715);
  not g49073 (n_22899, n8365);
  not g49074 (n_22900, n26558);
  and g49075 (n26559, n_22899, n_22900);
  and g49076 (n26560, n_11840, n_22900);
  not g49077 (n_22901, n26559);
  not g49078 (n_22902, n26560);
  and g49079 (n26561, n_22901, n_22902);
  not g49080 (n_22903, n26561);
  and g49081 (n26562, \a[50] , n_22903);
  and g49082 (n26563, n_7111, n26561);
  not g49083 (n_22904, n26562);
  not g49084 (n_22905, n26563);
  and g49085 (n26564, n_22904, n_22905);
  not g49086 (n_22906, n26557);
  not g49087 (n_22907, n26564);
  and g49088 (n26565, n_22906, n_22907);
  and g49089 (n26566, n26557, n26564);
  not g49090 (n_22908, n26565);
  not g49091 (n_22909, n26566);
  and g49092 (n26567, n_22908, n_22909);
  not g49093 (n_22910, n26556);
  and g49094 (n26568, n_22910, n26567);
  not g49095 (n_22911, n26568);
  and g49096 (n26569, n_22910, n_22911);
  and g49097 (n26570, n26567, n_22911);
  not g49098 (n_22912, n26569);
  not g49099 (n_22913, n26570);
  and g49100 (n26571, n_22912, n_22913);
  and g49101 (n26572, n_22818, n_22821);
  and g49102 (n26573, n26571, n26572);
  not g49103 (n_22914, n26571);
  not g49104 (n_22915, n26572);
  and g49105 (n26574, n_22914, n_22915);
  not g49106 (n_22916, n26573);
  not g49107 (n_22917, n26574);
  and g49108 (n26575, n_22916, n_22917);
  and g49109 (n26576, n_22827, n_22830);
  not g49110 (n_22918, n26576);
  and g49111 (n26577, n26575, n_22918);
  not g49112 (n_22919, n26575);
  and g49113 (n26578, n_22919, n26576);
  not g49114 (n_22920, n26577);
  not g49115 (n_22921, n26578);
  and g49116 (\f[113] , n_22920, n_22921);
  and g49117 (n26580, n_22877, n_22880);
  and g49118 (n26581, \b[60] , n10426);
  and g49119 (n26582, \b[58] , n10796);
  and g49120 (n26583, \b[59] , n10421);
  and g49126 (n26586, n10429, n12211);
  not g49129 (n_22926, n26587);
  and g49130 (n26588, \a[56] , n_22926);
  not g49131 (n_22927, n26588);
  and g49132 (n26589, \a[56] , n_22927);
  and g49133 (n26590, n_22926, n_22927);
  not g49134 (n_22928, n26589);
  not g49135 (n_22929, n26590);
  and g49136 (n26591, n_22928, n_22929);
  and g49137 (n26592, n_22862, n_22874);
  and g49138 (n26593, \b[57] , n11531);
  and g49139 (n26594, \b[55] , n11896);
  and g49140 (n26595, \b[56] , n11526);
  and g49146 (n26598, n11410, n11534);
  not g49149 (n_22934, n26599);
  and g49150 (n26600, \a[59] , n_22934);
  not g49151 (n_22935, n26600);
  and g49152 (n26601, \a[59] , n_22935);
  and g49153 (n26602, n_22934, n_22935);
  not g49154 (n_22936, n26601);
  not g49155 (n_22937, n26602);
  and g49156 (n26603, n_22936, n_22937);
  and g49157 (n26604, \b[54] , n12668);
  and g49158 (n26605, \b[52] , n13047);
  and g49159 (n26606, \b[53] , n12663);
  and g49165 (n26609, n9998, n12671);
  not g49168 (n_22942, n26610);
  and g49169 (n26611, \a[62] , n_22942);
  not g49170 (n_22943, n26611);
  and g49171 (n26612, \a[62] , n_22943);
  and g49172 (n26613, n_22942, n_22943);
  not g49173 (n_22944, n26612);
  not g49174 (n_22945, n26613);
  and g49175 (n26614, n_22944, n_22945);
  and g49176 (n26615, n_22851, n_22856);
  and g49177 (n26616, \b[50] , n13903);
  and g49178 (n26617, \b[51] , n_11555);
  not g49179 (n_22946, n26616);
  not g49180 (n_22947, n26617);
  and g49181 (n26618, n_22946, n_22947);
  not g49182 (n_22948, n26618);
  and g49183 (n26619, n_7111, n_22948);
  and g49184 (n26620, \a[50] , n26618);
  not g49185 (n_22949, n26619);
  not g49186 (n_22950, n26620);
  and g49187 (n26621, n_22949, n_22950);
  and g49188 (n26622, n_22777, n26621);
  not g49189 (n_22951, n26621);
  and g49190 (n26623, n26422, n_22951);
  not g49191 (n_22952, n26622);
  not g49192 (n_22953, n26623);
  and g49193 (n26624, n_22952, n_22953);
  not g49194 (n_22954, n26615);
  and g49195 (n26625, n_22954, n26624);
  not g49196 (n_22955, n26625);
  and g49197 (n26626, n_22954, n_22955);
  and g49198 (n26627, n26624, n_22955);
  not g49199 (n_22956, n26626);
  not g49200 (n_22957, n26627);
  and g49201 (n26628, n_22956, n_22957);
  not g49202 (n_22958, n26614);
  not g49203 (n_22959, n26628);
  and g49204 (n26629, n_22958, n_22959);
  and g49205 (n26630, n26614, n_22957);
  and g49206 (n26631, n_22956, n26630);
  not g49207 (n_22960, n26629);
  not g49208 (n_22961, n26631);
  and g49209 (n26632, n_22960, n_22961);
  not g49210 (n_22962, n26603);
  and g49211 (n26633, n_22962, n26632);
  not g49212 (n_22963, n26633);
  and g49213 (n26634, n_22962, n_22963);
  and g49214 (n26635, n26632, n_22963);
  not g49215 (n_22964, n26634);
  not g49216 (n_22965, n26635);
  and g49217 (n26636, n_22964, n_22965);
  not g49218 (n_22966, n26592);
  not g49219 (n_22967, n26636);
  and g49220 (n26637, n_22966, n_22967);
  and g49221 (n26638, n26592, n_22965);
  and g49222 (n26639, n_22964, n26638);
  not g49223 (n_22968, n26637);
  not g49224 (n_22969, n26639);
  and g49225 (n26640, n_22968, n_22969);
  not g49226 (n_22970, n26591);
  and g49227 (n26641, n_22970, n26640);
  not g49228 (n_22971, n26640);
  and g49229 (n26642, n26591, n_22971);
  not g49230 (n_22972, n26641);
  not g49231 (n_22973, n26642);
  and g49232 (n26643, n_22972, n_22973);
  not g49233 (n_22974, n26580);
  and g49234 (n26644, n_22974, n26643);
  not g49235 (n_22975, n26643);
  and g49236 (n26645, n26580, n_22975);
  not g49237 (n_22976, n26644);
  not g49238 (n_22977, n26645);
  and g49239 (n26646, n_22976, n_22977);
  and g49240 (n26647, \b[63] , n9339);
  and g49241 (n26648, \b[61] , n9732);
  and g49242 (n26649, \b[62] , n9334);
  and g49248 (n26652, n9342, n13771);
  not g49251 (n_22982, n26653);
  and g49252 (n26654, \a[53] , n_22982);
  not g49253 (n_22983, n26654);
  and g49254 (n26655, \a[53] , n_22983);
  and g49255 (n26656, n_22982, n_22983);
  not g49256 (n_22984, n26655);
  not g49257 (n_22985, n26656);
  and g49258 (n26657, n_22984, n_22985);
  not g49259 (n_22986, n26657);
  and g49260 (n26658, n26646, n_22986);
  not g49261 (n_22987, n26658);
  and g49262 (n26659, n26646, n_22987);
  and g49263 (n26660, n_22986, n_22987);
  not g49264 (n_22988, n26659);
  not g49265 (n_22989, n26660);
  and g49266 (n26661, n_22988, n_22989);
  and g49267 (n26662, n_22886, n_22896);
  and g49268 (n26663, n26661, n26662);
  not g49269 (n_22990, n26661);
  not g49270 (n_22991, n26662);
  and g49271 (n26664, n_22990, n_22991);
  not g49272 (n_22992, n26663);
  not g49273 (n_22993, n26664);
  and g49274 (n26665, n_22992, n_22993);
  and g49275 (n26666, n_22908, n_22911);
  not g49276 (n_22994, n26665);
  and g49277 (n26667, n_22994, n26666);
  not g49278 (n_22995, n26666);
  and g49279 (n26668, n26665, n_22995);
  not g49280 (n_22996, n26667);
  not g49281 (n_22997, n26668);
  and g49282 (n26669, n_22996, n_22997);
  and g49283 (n26670, n_22917, n_22920);
  not g49284 (n_22998, n26670);
  and g49285 (n26671, n26669, n_22998);
  not g49286 (n_22999, n26669);
  and g49287 (n26672, n_22999, n26670);
  not g49288 (n_23000, n26671);
  not g49289 (n_23001, n26672);
  and g49290 (\f[114] , n_23000, n_23001);
  and g49291 (n26674, \b[62] , n9732);
  and g49292 (n26675, \b[63] , n9334);
  not g49293 (n_23002, n26674);
  not g49294 (n_23003, n26675);
  and g49295 (n26676, n_23002, n_23003);
  and g49296 (n26677, n9342, n_11843);
  not g49297 (n_23004, n26677);
  and g49298 (n26678, n26676, n_23004);
  not g49299 (n_23005, n26678);
  and g49300 (n26679, \a[53] , n_23005);
  not g49301 (n_23006, n26679);
  and g49302 (n26680, \a[53] , n_23006);
  and g49303 (n26681, n_23005, n_23006);
  not g49304 (n_23007, n26680);
  not g49305 (n_23008, n26681);
  and g49306 (n26682, n_23007, n_23008);
  and g49307 (n26683, n_22972, n_22976);
  and g49308 (n26684, \b[61] , n10426);
  and g49309 (n26685, \b[59] , n10796);
  and g49310 (n26686, \b[60] , n10421);
  and g49316 (n26689, n10429, n12969);
  not g49319 (n_23013, n26690);
  and g49320 (n26691, \a[56] , n_23013);
  not g49321 (n_23014, n26691);
  and g49322 (n26692, \a[56] , n_23014);
  and g49323 (n26693, n_23013, n_23014);
  not g49324 (n_23015, n26692);
  not g49325 (n_23016, n26693);
  and g49326 (n26694, n_23015, n_23016);
  and g49327 (n26695, n_22963, n_22968);
  and g49328 (n26696, \b[58] , n11531);
  and g49329 (n26697, \b[56] , n11896);
  and g49330 (n26698, \b[57] , n11526);
  and g49336 (n26701, n11436, n11534);
  not g49339 (n_23021, n26702);
  and g49340 (n26703, \a[59] , n_23021);
  not g49341 (n_23022, n26703);
  and g49342 (n26704, \a[59] , n_23022);
  and g49343 (n26705, n_23021, n_23022);
  not g49344 (n_23023, n26704);
  not g49345 (n_23024, n26705);
  and g49346 (n26706, n_23023, n_23024);
  and g49347 (n26707, n_22955, n_22960);
  and g49348 (n26708, \b[51] , n13903);
  and g49349 (n26709, \b[52] , n_11555);
  not g49350 (n_23025, n26708);
  not g49351 (n_23026, n26709);
  and g49352 (n26710, n_23025, n_23026);
  and g49353 (n26711, n_22949, n_22952);
  not g49354 (n_23027, n26710);
  and g49355 (n26712, n_23027, n26711);
  not g49356 (n_23028, n26711);
  and g49357 (n26713, n26710, n_23028);
  not g49358 (n_23029, n26712);
  not g49359 (n_23030, n26713);
  and g49360 (n26714, n_23029, n_23030);
  and g49361 (n26715, \b[55] , n12668);
  and g49362 (n26716, \b[53] , n13047);
  and g49363 (n26717, \b[54] , n12663);
  and g49369 (n26720, n10684, n12671);
  not g49372 (n_23035, n26721);
  and g49373 (n26722, \a[62] , n_23035);
  not g49374 (n_23036, n26722);
  and g49375 (n26723, \a[62] , n_23036);
  and g49376 (n26724, n_23035, n_23036);
  not g49377 (n_23037, n26723);
  not g49378 (n_23038, n26724);
  and g49379 (n26725, n_23037, n_23038);
  not g49380 (n_23039, n26714);
  and g49381 (n26726, n_23039, n26725);
  not g49382 (n_23040, n26725);
  and g49383 (n26727, n26714, n_23040);
  not g49384 (n_23041, n26726);
  not g49385 (n_23042, n26727);
  and g49386 (n26728, n_23041, n_23042);
  not g49387 (n_23043, n26707);
  and g49388 (n26729, n_23043, n26728);
  not g49389 (n_23044, n26728);
  and g49390 (n26730, n26707, n_23044);
  not g49391 (n_23045, n26729);
  not g49392 (n_23046, n26730);
  and g49393 (n26731, n_23045, n_23046);
  not g49394 (n_23047, n26706);
  and g49395 (n26732, n_23047, n26731);
  not g49396 (n_23048, n26731);
  and g49397 (n26733, n26706, n_23048);
  not g49398 (n_23049, n26732);
  not g49399 (n_23050, n26733);
  and g49400 (n26734, n_23049, n_23050);
  not g49401 (n_23051, n26695);
  and g49402 (n26735, n_23051, n26734);
  not g49403 (n_23052, n26735);
  and g49404 (n26736, n_23051, n_23052);
  and g49405 (n26737, n26734, n_23052);
  not g49406 (n_23053, n26736);
  not g49407 (n_23054, n26737);
  and g49408 (n26738, n_23053, n_23054);
  not g49409 (n_23055, n26694);
  not g49410 (n_23056, n26738);
  and g49411 (n26739, n_23055, n_23056);
  and g49412 (n26740, n26694, n_23054);
  and g49413 (n26741, n_23053, n26740);
  not g49414 (n_23057, n26739);
  not g49415 (n_23058, n26741);
  and g49416 (n26742, n_23057, n_23058);
  not g49417 (n_23059, n26683);
  and g49418 (n26743, n_23059, n26742);
  not g49419 (n_23060, n26742);
  and g49420 (n26744, n26683, n_23060);
  not g49421 (n_23061, n26743);
  not g49422 (n_23062, n26744);
  and g49423 (n26745, n_23061, n_23062);
  not g49424 (n_23063, n26682);
  and g49425 (n26746, n_23063, n26745);
  not g49426 (n_23064, n26746);
  and g49427 (n26747, n26745, n_23064);
  and g49428 (n26748, n_23063, n_23064);
  not g49429 (n_23065, n26747);
  not g49430 (n_23066, n26748);
  and g49431 (n26749, n_23065, n_23066);
  and g49432 (n26750, n_22987, n_22993);
  and g49433 (n26751, n26749, n26750);
  not g49434 (n_23067, n26749);
  not g49435 (n_23068, n26750);
  and g49436 (n26752, n_23067, n_23068);
  not g49437 (n_23069, n26751);
  not g49438 (n_23070, n26752);
  and g49439 (n26753, n_23069, n_23070);
  and g49440 (n26754, n_22997, n_23000);
  not g49441 (n_23071, n26754);
  and g49442 (n26755, n26753, n_23071);
  not g49443 (n_23072, n26753);
  and g49444 (n26756, n_23072, n26754);
  not g49445 (n_23073, n26755);
  not g49446 (n_23074, n26756);
  and g49447 (\f[115] , n_23073, n_23074);
  and g49448 (n26758, n_23045, n_23049);
  and g49449 (n26759, n_23030, n_23042);
  and g49450 (n26760, \b[52] , n13903);
  and g49451 (n26761, \b[53] , n_11555);
  not g49452 (n_23075, n26760);
  not g49453 (n_23076, n26761);
  and g49454 (n26762, n_23075, n_23076);
  not g49455 (n_23077, n26762);
  and g49456 (n26763, n26710, n_23077);
  and g49457 (n26764, n_23027, n26762);
  not g49458 (n_23078, n26759);
  not g49459 (n_23079, n26764);
  and g49460 (n26765, n_23078, n_23079);
  not g49461 (n_23080, n26763);
  and g49462 (n26766, n_23080, n26765);
  not g49463 (n_23081, n26766);
  and g49464 (n26767, n_23078, n_23081);
  and g49465 (n26768, n_23079, n_23081);
  and g49466 (n26769, n_23080, n26768);
  not g49467 (n_23082, n26767);
  not g49468 (n_23083, n26769);
  and g49469 (n26770, n_23082, n_23083);
  and g49470 (n26771, \b[56] , n12668);
  and g49471 (n26772, \b[54] , n13047);
  and g49472 (n26773, \b[55] , n12663);
  and g49478 (n26776, n10708, n12671);
  not g49481 (n_23088, n26777);
  and g49482 (n26778, \a[62] , n_23088);
  not g49483 (n_23089, n26778);
  and g49484 (n26779, \a[62] , n_23089);
  and g49485 (n26780, n_23088, n_23089);
  not g49486 (n_23090, n26779);
  not g49487 (n_23091, n26780);
  and g49488 (n26781, n_23090, n_23091);
  not g49489 (n_23092, n26770);
  and g49490 (n26782, n_23092, n26781);
  not g49491 (n_23093, n26781);
  and g49492 (n26783, n26770, n_23093);
  not g49493 (n_23094, n26782);
  not g49494 (n_23095, n26783);
  and g49495 (n26784, n_23094, n_23095);
  and g49496 (n26785, \b[59] , n11531);
  and g49497 (n26786, \b[57] , n11896);
  and g49498 (n26787, \b[58] , n11526);
  and g49504 (n26790, n11534, n12179);
  not g49507 (n_23100, n26791);
  and g49508 (n26792, \a[59] , n_23100);
  not g49509 (n_23101, n26792);
  and g49510 (n26793, \a[59] , n_23101);
  and g49511 (n26794, n_23100, n_23101);
  not g49512 (n_23102, n26793);
  not g49513 (n_23103, n26794);
  and g49514 (n26795, n_23102, n_23103);
  not g49515 (n_23104, n26784);
  not g49516 (n_23105, n26795);
  and g49517 (n26796, n_23104, n_23105);
  and g49518 (n26797, n26784, n26795);
  not g49519 (n_23106, n26796);
  not g49520 (n_23107, n26797);
  and g49521 (n26798, n_23106, n_23107);
  not g49522 (n_23108, n26798);
  and g49523 (n26799, n26758, n_23108);
  not g49524 (n_23109, n26758);
  and g49525 (n26800, n_23109, n26798);
  not g49526 (n_23110, n26799);
  not g49527 (n_23111, n26800);
  and g49528 (n26801, n_23110, n_23111);
  and g49529 (n26802, \b[62] , n10426);
  and g49530 (n26803, \b[60] , n10796);
  and g49531 (n26804, \b[61] , n10421);
  and g49537 (n26807, n10429, n13370);
  not g49540 (n_23116, n26808);
  and g49541 (n26809, \a[56] , n_23116);
  not g49542 (n_23117, n26809);
  and g49543 (n26810, \a[56] , n_23117);
  and g49544 (n26811, n_23116, n_23117);
  not g49545 (n_23118, n26810);
  not g49546 (n_23119, n26811);
  and g49547 (n26812, n_23118, n_23119);
  not g49548 (n_23120, n26812);
  and g49549 (n26813, n26801, n_23120);
  not g49550 (n_23121, n26813);
  and g49551 (n26814, n26801, n_23121);
  and g49552 (n26815, n_23120, n_23121);
  not g49553 (n_23122, n26814);
  not g49554 (n_23123, n26815);
  and g49555 (n26816, n_23122, n_23123);
  and g49556 (n26817, n_23052, n_23057);
  and g49557 (n26818, \b[63] , n9732);
  not g49558 (n_23124, n9342);
  not g49559 (n_23125, n26818);
  and g49560 (n26819, n_23124, n_23125);
  and g49561 (n26820, n_11840, n_23125);
  not g49562 (n_23126, n26819);
  not g49563 (n_23127, n26820);
  and g49564 (n26821, n_23126, n_23127);
  not g49565 (n_23128, n26821);
  and g49566 (n26822, \a[53] , n_23128);
  and g49567 (n26823, n_7957, n26821);
  not g49568 (n_23129, n26822);
  not g49569 (n_23130, n26823);
  and g49570 (n26824, n_23129, n_23130);
  not g49571 (n_23131, n26817);
  not g49572 (n_23132, n26824);
  and g49573 (n26825, n_23131, n_23132);
  and g49574 (n26826, n26817, n26824);
  not g49575 (n_23133, n26825);
  not g49576 (n_23134, n26826);
  and g49577 (n26827, n_23133, n_23134);
  not g49578 (n_23135, n26816);
  and g49579 (n26828, n_23135, n26827);
  not g49580 (n_23136, n26828);
  and g49581 (n26829, n_23135, n_23136);
  and g49582 (n26830, n26827, n_23136);
  not g49583 (n_23137, n26829);
  not g49584 (n_23138, n26830);
  and g49585 (n26831, n_23137, n_23138);
  and g49586 (n26832, n_23061, n_23064);
  and g49587 (n26833, n26831, n26832);
  not g49588 (n_23139, n26831);
  not g49589 (n_23140, n26832);
  and g49590 (n26834, n_23139, n_23140);
  not g49591 (n_23141, n26833);
  not g49592 (n_23142, n26834);
  and g49593 (n26835, n_23141, n_23142);
  and g49594 (n26836, n_23070, n_23073);
  not g49595 (n_23143, n26836);
  and g49596 (n26837, n26835, n_23143);
  not g49597 (n_23144, n26835);
  and g49598 (n26838, n_23144, n26836);
  not g49599 (n_23145, n26837);
  not g49600 (n_23146, n26838);
  and g49601 (\f[116] , n_23145, n_23146);
  and g49602 (n26840, n_23142, n_23145);
  and g49603 (n26841, n_23133, n_23136);
  and g49604 (n26842, n_23111, n_23121);
  and g49605 (n26843, \b[63] , n10426);
  and g49606 (n26844, \b[61] , n10796);
  and g49607 (n26845, \b[62] , n10421);
  and g49613 (n26848, n10429, n13771);
  not g49616 (n_23151, n26849);
  and g49617 (n26850, \a[56] , n_23151);
  not g49618 (n_23152, n26850);
  and g49619 (n26851, \a[56] , n_23152);
  and g49620 (n26852, n_23151, n_23152);
  not g49621 (n_23153, n26851);
  not g49622 (n_23154, n26852);
  and g49623 (n26853, n_23153, n_23154);
  not g49624 (n_23155, n26842);
  not g49625 (n_23156, n26853);
  and g49626 (n26854, n_23155, n_23156);
  not g49627 (n_23157, n26854);
  and g49628 (n26855, n_23155, n_23157);
  and g49629 (n26856, n_23156, n_23157);
  not g49630 (n_23158, n26855);
  not g49631 (n_23159, n26856);
  and g49632 (n26857, n_23158, n_23159);
  and g49633 (n26858, n_23092, n_23093);
  not g49634 (n_23160, n26858);
  and g49635 (n26859, n_23106, n_23160);
  and g49636 (n26860, \b[60] , n11531);
  and g49637 (n26861, \b[58] , n11896);
  and g49638 (n26862, \b[59] , n11526);
  and g49644 (n26865, n11534, n12211);
  not g49647 (n_23165, n26866);
  and g49648 (n26867, \a[59] , n_23165);
  not g49649 (n_23166, n26867);
  and g49650 (n26868, \a[59] , n_23166);
  and g49651 (n26869, n_23165, n_23166);
  not g49652 (n_23167, n26868);
  not g49653 (n_23168, n26869);
  and g49654 (n26870, n_23167, n_23168);
  and g49655 (n26871, \a[53] , n_23077);
  and g49656 (n26872, n_7957, n26762);
  not g49657 (n_23169, n26871);
  not g49658 (n_23170, n26872);
  and g49659 (n26873, n_23169, n_23170);
  and g49660 (n26874, \b[53] , n13903);
  and g49661 (n26875, \b[54] , n_11555);
  not g49662 (n_23171, n26874);
  not g49663 (n_23172, n26875);
  and g49664 (n26876, n_23171, n_23172);
  and g49665 (n26877, n26873, n26876);
  not g49666 (n_23173, n26873);
  not g49667 (n_23174, n26876);
  and g49668 (n26878, n_23173, n_23174);
  not g49669 (n_23175, n26877);
  not g49670 (n_23176, n26878);
  and g49671 (n26879, n_23175, n_23176);
  and g49672 (n26880, \b[57] , n12668);
  and g49673 (n26881, \b[55] , n13047);
  and g49674 (n26882, \b[56] , n12663);
  and g49680 (n26885, n11410, n12671);
  not g49683 (n_23181, n26886);
  and g49684 (n26887, \a[62] , n_23181);
  not g49685 (n_23182, n26887);
  and g49686 (n26888, \a[62] , n_23182);
  and g49687 (n26889, n_23181, n_23182);
  not g49688 (n_23183, n26888);
  not g49689 (n_23184, n26889);
  and g49690 (n26890, n_23183, n_23184);
  not g49691 (n_23185, n26890);
  and g49692 (n26891, n26879, n_23185);
  not g49693 (n_23186, n26891);
  and g49694 (n26892, n26879, n_23186);
  and g49695 (n26893, n_23185, n_23186);
  not g49696 (n_23187, n26892);
  not g49697 (n_23188, n26893);
  and g49698 (n26894, n_23187, n_23188);
  not g49699 (n_23189, n26768);
  not g49700 (n_23190, n26894);
  and g49701 (n26895, n_23189, n_23190);
  and g49702 (n26896, n26768, n26894);
  not g49703 (n_23191, n26895);
  not g49704 (n_23192, n26896);
  and g49705 (n26897, n_23191, n_23192);
  not g49706 (n_23193, n26870);
  and g49707 (n26898, n_23193, n26897);
  not g49708 (n_23194, n26898);
  and g49709 (n26899, n_23193, n_23194);
  and g49710 (n26900, n26897, n_23194);
  not g49711 (n_23195, n26899);
  not g49712 (n_23196, n26900);
  and g49713 (n26901, n_23195, n_23196);
  not g49714 (n_23197, n26859);
  not g49715 (n_23198, n26901);
  and g49716 (n26902, n_23197, n_23198);
  not g49717 (n_23199, n26902);
  and g49718 (n26903, n_23197, n_23199);
  and g49719 (n26904, n_23198, n_23199);
  not g49720 (n_23200, n26903);
  not g49721 (n_23201, n26904);
  and g49722 (n26905, n_23200, n_23201);
  not g49723 (n_23202, n26857);
  and g49724 (n26906, n_23202, n26905);
  not g49725 (n_23203, n26905);
  and g49726 (n26907, n26857, n_23203);
  not g49727 (n_23204, n26906);
  not g49728 (n_23205, n26907);
  and g49729 (n26908, n_23204, n_23205);
  not g49730 (n_23206, n26841);
  not g49731 (n_23207, n26908);
  and g49732 (n26909, n_23206, n_23207);
  and g49733 (n26910, n26841, n26908);
  not g49734 (n_23208, n26909);
  not g49735 (n_23209, n26910);
  and g49736 (n26911, n_23208, n_23209);
  not g49737 (n_23210, n26840);
  and g49738 (n26912, n_23210, n26911);
  not g49739 (n_23211, n26911);
  and g49740 (n26913, n26840, n_23211);
  not g49741 (n_23212, n26912);
  not g49742 (n_23213, n26913);
  and g49743 (\f[117] , n_23212, n_23213);
  and g49744 (n26915, \b[62] , n10796);
  and g49745 (n26916, \b[63] , n10421);
  not g49746 (n_23214, n26915);
  not g49747 (n_23215, n26916);
  and g49748 (n26917, n_23214, n_23215);
  and g49749 (n26918, n10429, n_11843);
  not g49750 (n_23216, n26918);
  and g49751 (n26919, n26917, n_23216);
  not g49752 (n_23217, n26919);
  and g49753 (n26920, \a[56] , n_23217);
  not g49754 (n_23218, n26920);
  and g49755 (n26921, \a[56] , n_23218);
  and g49756 (n26922, n_23217, n_23218);
  not g49757 (n_23219, n26921);
  not g49758 (n_23220, n26922);
  and g49759 (n26923, n_23219, n_23220);
  and g49760 (n26924, n_23194, n_23199);
  and g49761 (n26925, \b[61] , n11531);
  and g49762 (n26926, \b[59] , n11896);
  and g49763 (n26927, \b[60] , n11526);
  and g49769 (n26930, n11534, n12969);
  not g49772 (n_23225, n26931);
  and g49773 (n26932, \a[59] , n_23225);
  not g49774 (n_23226, n26932);
  and g49775 (n26933, \a[59] , n_23226);
  and g49776 (n26934, n_23225, n_23226);
  not g49777 (n_23227, n26933);
  not g49778 (n_23228, n26934);
  and g49779 (n26935, n_23227, n_23228);
  and g49780 (n26936, n_23186, n_23191);
  and g49781 (n26937, \b[54] , n13903);
  and g49782 (n26938, \b[55] , n_11555);
  not g49783 (n_23229, n26937);
  not g49784 (n_23230, n26938);
  and g49785 (n26939, n_23229, n_23230);
  and g49786 (n26940, n_7957, n_23077);
  not g49787 (n_23231, n26940);
  and g49788 (n26941, n_23176, n_23231);
  not g49789 (n_23232, n26941);
  and g49790 (n26942, n26939, n_23232);
  not g49791 (n_23233, n26939);
  and g49792 (n26943, n_23233, n26941);
  not g49793 (n_23234, n26942);
  not g49794 (n_23235, n26943);
  and g49795 (n26944, n_23234, n_23235);
  and g49796 (n26945, \b[58] , n12668);
  and g49797 (n26946, \b[56] , n13047);
  and g49798 (n26947, \b[57] , n12663);
  not g49799 (n_23236, n26946);
  not g49800 (n_23237, n26947);
  and g49801 (n26948, n_23236, n_23237);
  not g49802 (n_23238, n26945);
  and g49803 (n26949, n_23238, n26948);
  and g49804 (n26950, n_12644, n26949);
  and g49805 (n26951, n_13160, n26949);
  not g49806 (n_23239, n26950);
  not g49807 (n_23240, n26951);
  and g49808 (n26952, n_23239, n_23240);
  not g49809 (n_23241, n26952);
  and g49810 (n26953, \a[62] , n_23241);
  and g49811 (n26954, n_10843, n26952);
  not g49812 (n_23242, n26953);
  not g49813 (n_23243, n26954);
  and g49814 (n26955, n_23242, n_23243);
  not g49815 (n_23244, n26955);
  and g49816 (n26956, n26944, n_23244);
  not g49817 (n_23245, n26944);
  and g49818 (n26957, n_23245, n26955);
  not g49819 (n_23246, n26956);
  not g49820 (n_23247, n26957);
  and g49821 (n26958, n_23246, n_23247);
  not g49822 (n_23248, n26936);
  and g49823 (n26959, n_23248, n26958);
  not g49824 (n_23249, n26959);
  and g49825 (n26960, n_23248, n_23249);
  and g49826 (n26961, n26958, n_23249);
  not g49827 (n_23250, n26960);
  not g49828 (n_23251, n26961);
  and g49829 (n26962, n_23250, n_23251);
  not g49830 (n_23252, n26935);
  not g49831 (n_23253, n26962);
  and g49832 (n26963, n_23252, n_23253);
  and g49833 (n26964, n26935, n_23251);
  and g49834 (n26965, n_23250, n26964);
  not g49835 (n_23254, n26963);
  not g49836 (n_23255, n26965);
  and g49837 (n26966, n_23254, n_23255);
  not g49838 (n_23256, n26924);
  and g49839 (n26967, n_23256, n26966);
  not g49840 (n_23257, n26966);
  and g49841 (n26968, n26924, n_23257);
  not g49842 (n_23258, n26967);
  not g49843 (n_23259, n26968);
  and g49844 (n26969, n_23258, n_23259);
  not g49845 (n_23260, n26923);
  and g49846 (n26970, n_23260, n26969);
  not g49847 (n_23261, n26970);
  and g49848 (n26971, n26969, n_23261);
  and g49849 (n26972, n_23260, n_23261);
  not g49850 (n_23262, n26971);
  not g49851 (n_23263, n26972);
  and g49852 (n26973, n_23262, n_23263);
  and g49853 (n26974, n_23202, n_23203);
  not g49854 (n_23264, n26974);
  and g49855 (n26975, n_23157, n_23264);
  not g49856 (n_23265, n26973);
  not g49857 (n_23266, n26975);
  and g49858 (n26976, n_23265, n_23266);
  not g49859 (n_23267, n26976);
  and g49860 (n26977, n_23265, n_23267);
  and g49861 (n26978, n_23266, n_23267);
  not g49862 (n_23268, n26977);
  not g49863 (n_23269, n26978);
  and g49864 (n26979, n_23268, n_23269);
  and g49865 (n26980, n_23208, n_23212);
  not g49866 (n_23270, n26979);
  not g49867 (n_23271, n26980);
  and g49868 (n26981, n_23270, n_23271);
  and g49869 (n26982, n26979, n26980);
  not g49870 (n_23272, n26981);
  not g49871 (n_23273, n26982);
  and g49872 (\f[118] , n_23272, n_23273);
  and g49873 (n26984, \b[59] , n12668);
  and g49874 (n26985, \b[57] , n13047);
  and g49875 (n26986, \b[58] , n12663);
  and g49881 (n26989, n12179, n12671);
  not g49884 (n_23278, n26990);
  and g49885 (n26991, \a[62] , n_23278);
  not g49886 (n_23279, n26991);
  and g49887 (n26992, \a[62] , n_23279);
  and g49888 (n26993, n_23278, n_23279);
  not g49889 (n_23280, n26992);
  not g49890 (n_23281, n26993);
  and g49891 (n26994, n_23280, n_23281);
  and g49892 (n26995, \b[55] , n13903);
  and g49893 (n26996, \b[56] , n_11555);
  not g49894 (n_23282, n26995);
  not g49895 (n_23283, n26996);
  and g49896 (n26997, n_23282, n_23283);
  not g49897 (n_23284, n26997);
  and g49898 (n26998, n26939, n_23284);
  not g49899 (n_23285, n26998);
  and g49900 (n26999, n26939, n_23285);
  and g49901 (n27000, n_23284, n_23285);
  not g49902 (n_23286, n26999);
  not g49903 (n_23287, n27000);
  and g49904 (n27001, n_23286, n_23287);
  not g49905 (n_23288, n26994);
  not g49906 (n_23289, n27001);
  and g49907 (n27002, n_23288, n_23289);
  not g49908 (n_23290, n27002);
  and g49909 (n27003, n_23288, n_23290);
  and g49910 (n27004, n_23289, n_23290);
  not g49911 (n_23291, n27003);
  not g49912 (n_23292, n27004);
  and g49913 (n27005, n_23291, n_23292);
  and g49914 (n27006, n_23234, n_23246);
  and g49915 (n27007, n27005, n27006);
  not g49916 (n_23293, n27005);
  not g49917 (n_23294, n27006);
  and g49918 (n27008, n_23293, n_23294);
  not g49919 (n_23295, n27007);
  not g49920 (n_23296, n27008);
  and g49921 (n27009, n_23295, n_23296);
  and g49922 (n27010, \b[62] , n11531);
  and g49923 (n27011, \b[60] , n11896);
  and g49924 (n27012, \b[61] , n11526);
  and g49930 (n27015, n11534, n13370);
  not g49933 (n_23301, n27016);
  and g49934 (n27017, \a[59] , n_23301);
  not g49935 (n_23302, n27017);
  and g49936 (n27018, \a[59] , n_23302);
  and g49937 (n27019, n_23301, n_23302);
  not g49938 (n_23303, n27018);
  not g49939 (n_23304, n27019);
  and g49940 (n27020, n_23303, n_23304);
  not g49941 (n_23305, n27020);
  and g49942 (n27021, n27009, n_23305);
  not g49943 (n_23306, n27021);
  and g49944 (n27022, n27009, n_23306);
  and g49945 (n27023, n_23305, n_23306);
  not g49946 (n_23307, n27022);
  not g49947 (n_23308, n27023);
  and g49948 (n27024, n_23307, n_23308);
  and g49949 (n27025, n_23249, n_23254);
  and g49950 (n27026, \b[63] , n10796);
  not g49951 (n_23309, n10429);
  not g49952 (n_23310, n27026);
  and g49953 (n27027, n_23309, n_23310);
  and g49954 (n27028, n_11840, n_23310);
  not g49955 (n_23311, n27027);
  not g49956 (n_23312, n27028);
  and g49957 (n27029, n_23311, n_23312);
  not g49958 (n_23313, n27029);
  and g49959 (n27030, \a[56] , n_23313);
  and g49960 (n27031, n_8895, n27029);
  not g49961 (n_23314, n27030);
  not g49962 (n_23315, n27031);
  and g49963 (n27032, n_23314, n_23315);
  not g49964 (n_23316, n27025);
  not g49965 (n_23317, n27032);
  and g49966 (n27033, n_23316, n_23317);
  and g49967 (n27034, n27025, n27032);
  not g49968 (n_23318, n27033);
  not g49969 (n_23319, n27034);
  and g49970 (n27035, n_23318, n_23319);
  not g49971 (n_23320, n27024);
  and g49972 (n27036, n_23320, n27035);
  not g49973 (n_23321, n27036);
  and g49974 (n27037, n_23320, n_23321);
  and g49975 (n27038, n27035, n_23321);
  not g49976 (n_23322, n27037);
  not g49977 (n_23323, n27038);
  and g49978 (n27039, n_23322, n_23323);
  and g49979 (n27040, n_23258, n_23261);
  and g49980 (n27041, n27039, n27040);
  not g49981 (n_23324, n27039);
  not g49982 (n_23325, n27040);
  and g49983 (n27042, n_23324, n_23325);
  not g49984 (n_23326, n27041);
  not g49985 (n_23327, n27042);
  and g49986 (n27043, n_23326, n_23327);
  and g49987 (n27044, n_23267, n_23272);
  not g49988 (n_23328, n27044);
  and g49989 (n27045, n27043, n_23328);
  not g49990 (n_23329, n27043);
  and g49991 (n27046, n_23329, n27044);
  not g49992 (n_23330, n27045);
  not g49993 (n_23331, n27046);
  and g49994 (\f[119] , n_23330, n_23331);
  and g49995 (n27048, n_23296, n_23306);
  and g49996 (n27049, \b[63] , n11531);
  and g49997 (n27050, \b[61] , n11896);
  and g49998 (n27051, \b[62] , n11526);
  and g50004 (n27054, n11534, n13771);
  not g50007 (n_23336, n27055);
  and g50008 (n27056, \a[59] , n_23336);
  not g50009 (n_23337, n27056);
  and g50010 (n27057, \a[59] , n_23337);
  and g50011 (n27058, n_23336, n_23337);
  not g50012 (n_23338, n27057);
  not g50013 (n_23339, n27058);
  and g50014 (n27059, n_23338, n_23339);
  not g50015 (n_23340, n27048);
  not g50016 (n_23341, n27059);
  and g50017 (n27060, n_23340, n_23341);
  not g50018 (n_23342, n27060);
  and g50019 (n27061, n_23340, n_23342);
  and g50020 (n27062, n_23341, n_23342);
  not g50021 (n_23343, n27061);
  not g50022 (n_23344, n27062);
  and g50023 (n27063, n_23343, n_23344);
  and g50024 (n27064, \b[56] , n13903);
  and g50025 (n27065, \b[57] , n_11555);
  not g50026 (n_23345, n27064);
  not g50027 (n_23346, n27065);
  and g50028 (n27066, n_23345, n_23346);
  not g50029 (n_23347, n27066);
  and g50030 (n27067, n_8895, n_23347);
  not g50031 (n_23348, n27067);
  and g50032 (n27068, n_8895, n_23348);
  and g50033 (n27069, n_23347, n_23348);
  not g50034 (n_23349, n27068);
  not g50035 (n_23350, n27069);
  and g50036 (n27070, n_23349, n_23350);
  not g50037 (n_23351, n27070);
  and g50038 (n27071, n_23233, n_23351);
  not g50039 (n_23352, n27071);
  and g50040 (n27072, n_23233, n_23352);
  and g50041 (n27073, n_23351, n_23352);
  not g50042 (n_23353, n27072);
  not g50043 (n_23354, n27073);
  and g50044 (n27074, n_23353, n_23354);
  and g50045 (n27075, n_23285, n_23290);
  and g50046 (n27076, n27074, n27075);
  not g50047 (n_23355, n27074);
  not g50048 (n_23356, n27075);
  and g50049 (n27077, n_23355, n_23356);
  not g50050 (n_23357, n27076);
  not g50051 (n_23358, n27077);
  and g50052 (n27078, n_23357, n_23358);
  and g50053 (n27079, \b[60] , n12668);
  and g50054 (n27080, \b[58] , n13047);
  and g50055 (n27081, \b[59] , n12663);
  and g50061 (n27084, n12211, n12671);
  not g50064 (n_23363, n27085);
  and g50065 (n27086, \a[62] , n_23363);
  not g50066 (n_23364, n27086);
  and g50067 (n27087, \a[62] , n_23364);
  and g50068 (n27088, n_23363, n_23364);
  not g50069 (n_23365, n27087);
  not g50070 (n_23366, n27088);
  and g50071 (n27089, n_23365, n_23366);
  not g50072 (n_23367, n27089);
  and g50073 (n27090, n27078, n_23367);
  not g50074 (n_23368, n27078);
  and g50075 (n27091, n_23368, n27089);
  not g50076 (n_23369, n27063);
  not g50077 (n_23370, n27091);
  and g50078 (n27092, n_23369, n_23370);
  not g50079 (n_23371, n27090);
  and g50080 (n27093, n_23371, n27092);
  not g50081 (n_23372, n27093);
  and g50082 (n27094, n_23369, n_23372);
  and g50083 (n27095, n_23370, n_23372);
  and g50084 (n27096, n_23371, n27095);
  not g50085 (n_23373, n27094);
  not g50086 (n_23374, n27096);
  and g50087 (n27097, n_23373, n_23374);
  and g50088 (n27098, n_23318, n_23321);
  and g50089 (n27099, n27097, n27098);
  not g50090 (n_23375, n27097);
  not g50091 (n_23376, n27098);
  and g50092 (n27100, n_23375, n_23376);
  not g50093 (n_23377, n27099);
  not g50094 (n_23378, n27100);
  and g50095 (n27101, n_23377, n_23378);
  and g50096 (n27102, n_23327, n_23330);
  not g50097 (n_23379, n27102);
  and g50098 (n27103, n27101, n_23379);
  not g50099 (n_23380, n27101);
  and g50100 (n27104, n_23380, n27102);
  not g50101 (n_23381, n27103);
  not g50102 (n_23382, n27104);
  and g50103 (\f[120] , n_23381, n_23382);
  and g50104 (n27106, n_23358, n_23371);
  and g50105 (n27107, \b[57] , n13903);
  and g50106 (n27108, \b[58] , n_11555);
  not g50107 (n_23383, n27107);
  not g50108 (n_23384, n27108);
  and g50109 (n27109, n_23383, n_23384);
  and g50110 (n27110, n_23348, n_23352);
  not g50111 (n_23385, n27109);
  and g50112 (n27111, n_23385, n27110);
  not g50113 (n_23386, n27110);
  and g50114 (n27112, n27109, n_23386);
  not g50115 (n_23387, n27111);
  not g50116 (n_23388, n27112);
  and g50117 (n27113, n_23387, n_23388);
  and g50118 (n27114, \b[61] , n12668);
  and g50119 (n27115, \b[59] , n13047);
  and g50120 (n27116, \b[60] , n12663);
  not g50121 (n_23389, n27115);
  not g50122 (n_23390, n27116);
  and g50123 (n27117, n_23389, n_23390);
  not g50124 (n_23391, n27114);
  and g50125 (n27118, n_23391, n27117);
  and g50126 (n27119, n_12644, n27118);
  and g50127 (n27120, n_13180, n27118);
  not g50128 (n_23392, n27119);
  not g50129 (n_23393, n27120);
  and g50130 (n27121, n_23392, n_23393);
  not g50131 (n_23394, n27121);
  and g50132 (n27122, \a[62] , n_23394);
  and g50133 (n27123, n_10843, n27121);
  not g50134 (n_23395, n27122);
  not g50135 (n_23396, n27123);
  and g50136 (n27124, n_23395, n_23396);
  not g50137 (n_23397, n27124);
  and g50138 (n27125, n27113, n_23397);
  not g50139 (n_23398, n27113);
  and g50140 (n27126, n_23398, n27124);
  not g50141 (n_23399, n27125);
  not g50142 (n_23400, n27126);
  and g50143 (n27127, n_23399, n_23400);
  not g50144 (n_23401, n27106);
  and g50145 (n27128, n_23401, n27127);
  not g50146 (n_23402, n27127);
  and g50147 (n27129, n27106, n_23402);
  not g50148 (n_23403, n27128);
  not g50149 (n_23404, n27129);
  and g50150 (n27130, n_23403, n_23404);
  and g50151 (n27131, \b[62] , n11896);
  and g50152 (n27132, \b[63] , n11526);
  not g50153 (n_23405, n27131);
  not g50154 (n_23406, n27132);
  and g50155 (n27133, n_23405, n_23406);
  and g50156 (n27134, n11534, n_11843);
  not g50157 (n_23407, n27134);
  and g50158 (n27135, n27133, n_23407);
  not g50159 (n_23408, n27135);
  and g50160 (n27136, \a[59] , n_23408);
  not g50161 (n_23409, n27136);
  and g50162 (n27137, \a[59] , n_23409);
  and g50163 (n27138, n_23408, n_23409);
  not g50164 (n_23410, n27137);
  not g50165 (n_23411, n27138);
  and g50166 (n27139, n_23410, n_23411);
  not g50167 (n_23412, n27139);
  and g50168 (n27140, n27130, n_23412);
  not g50169 (n_23413, n27140);
  and g50170 (n27141, n27130, n_23413);
  and g50171 (n27142, n_23412, n_23413);
  not g50172 (n_23414, n27141);
  not g50173 (n_23415, n27142);
  and g50174 (n27143, n_23414, n_23415);
  and g50175 (n27144, n_23342, n_23372);
  and g50176 (n27145, n27143, n27144);
  not g50177 (n_23416, n27143);
  not g50178 (n_23417, n27144);
  and g50179 (n27146, n_23416, n_23417);
  not g50180 (n_23418, n27145);
  not g50181 (n_23419, n27146);
  and g50182 (n27147, n_23418, n_23419);
  and g50183 (n27148, n_23378, n_23381);
  not g50184 (n_23420, n27148);
  and g50185 (n27149, n27147, n_23420);
  not g50186 (n_23421, n27147);
  and g50187 (n27150, n_23421, n27148);
  not g50188 (n_23422, n27149);
  not g50189 (n_23423, n27150);
  and g50190 (\f[121] , n_23422, n_23423);
  and g50191 (n27152, n_23419, n_23422);
  and g50192 (n27153, n_23403, n_23413);
  and g50193 (n27154, n_23388, n_23399);
  and g50194 (n27155, \b[58] , n13903);
  and g50195 (n27156, \b[59] , n_11555);
  not g50196 (n_23424, n27155);
  not g50197 (n_23425, n27156);
  and g50198 (n27157, n_23424, n_23425);
  not g50199 (n_23426, n27157);
  and g50200 (n27158, n27109, n_23426);
  and g50201 (n27159, n_23385, n27157);
  not g50202 (n_23427, n27154);
  not g50203 (n_23428, n27159);
  and g50204 (n27160, n_23427, n_23428);
  not g50205 (n_23429, n27158);
  and g50206 (n27161, n_23429, n27160);
  not g50207 (n_23430, n27161);
  and g50208 (n27162, n_23427, n_23430);
  and g50209 (n27163, n_23428, n_23430);
  and g50210 (n27164, n_23429, n27163);
  not g50211 (n_23431, n27162);
  not g50212 (n_23432, n27164);
  and g50213 (n27165, n_23431, n_23432);
  and g50214 (n27166, \b[62] , n12668);
  and g50215 (n27167, \b[60] , n13047);
  and g50216 (n27168, \b[61] , n12663);
  and g50222 (n27171, n12671, n13370);
  not g50225 (n_23437, n27172);
  and g50226 (n27173, \a[62] , n_23437);
  not g50227 (n_23438, n27173);
  and g50228 (n27174, \a[62] , n_23438);
  and g50229 (n27175, n_23437, n_23438);
  not g50230 (n_23439, n27174);
  not g50231 (n_23440, n27175);
  and g50232 (n27176, n_23439, n_23440);
  and g50233 (n27177, \b[63] , n11896);
  and g50234 (n27178, n11534, n13797);
  not g50235 (n_23441, n27177);
  not g50236 (n_23442, n27178);
  and g50237 (n27179, n_23441, n_23442);
  not g50238 (n_23443, n27179);
  and g50239 (n27180, \a[59] , n_23443);
  not g50240 (n_23444, n27180);
  and g50241 (n27181, \a[59] , n_23444);
  and g50242 (n27182, n_23443, n_23444);
  not g50243 (n_23445, n27181);
  not g50244 (n_23446, n27182);
  and g50245 (n27183, n_23445, n_23446);
  not g50246 (n_23447, n27176);
  not g50247 (n_23448, n27183);
  and g50248 (n27184, n_23447, n_23448);
  not g50249 (n_23449, n27184);
  and g50250 (n27185, n_23447, n_23449);
  and g50251 (n27186, n_23448, n_23449);
  not g50252 (n_23450, n27185);
  not g50253 (n_23451, n27186);
  and g50254 (n27187, n_23450, n_23451);
  not g50255 (n_23452, n27165);
  and g50256 (n27188, n_23452, n27187);
  not g50257 (n_23453, n27187);
  and g50258 (n27189, n27165, n_23453);
  not g50259 (n_23454, n27188);
  not g50260 (n_23455, n27189);
  and g50261 (n27190, n_23454, n_23455);
  not g50262 (n_23456, n27153);
  not g50263 (n_23457, n27190);
  and g50264 (n27191, n_23456, n_23457);
  not g50265 (n_23458, n27191);
  and g50266 (n27192, n_23456, n_23458);
  and g50267 (n27193, n_23457, n_23458);
  not g50268 (n_23459, n27192);
  not g50269 (n_23460, n27193);
  and g50270 (n27194, n_23459, n_23460);
  not g50271 (n_23461, n27152);
  not g50272 (n_23462, n27194);
  and g50273 (n27195, n_23461, n_23462);
  and g50274 (n27196, n27152, n_23460);
  and g50275 (n27197, n_23459, n27196);
  not g50276 (n_23463, n27195);
  not g50277 (n_23464, n27197);
  and g50278 (\f[122] , n_23463, n_23464);
  and g50279 (n27199, n_23458, n_23463);
  and g50280 (n27200, n_23452, n_23453);
  not g50281 (n_23465, n27200);
  and g50282 (n27201, n_23449, n_23465);
  and g50283 (n27202, \a[59] , n_23426);
  and g50284 (n27203, n_9855, n27157);
  not g50285 (n_23466, n27202);
  not g50286 (n_23467, n27203);
  and g50287 (n27204, n_23466, n_23467);
  and g50288 (n27205, \b[59] , n13903);
  and g50289 (n27206, \b[60] , n_11555);
  not g50290 (n_23468, n27205);
  not g50291 (n_23469, n27206);
  and g50292 (n27207, n_23468, n_23469);
  and g50293 (n27208, n27204, n27207);
  not g50294 (n_23470, n27204);
  not g50295 (n_23471, n27207);
  and g50296 (n27209, n_23470, n_23471);
  not g50297 (n_23472, n27208);
  not g50298 (n_23473, n27209);
  and g50299 (n27210, n_23472, n_23473);
  and g50300 (n27211, \b[63] , n12668);
  and g50301 (n27212, \b[61] , n13047);
  and g50302 (n27213, \b[62] , n12663);
  and g50308 (n27216, n12671, n13771);
  not g50311 (n_23478, n27217);
  and g50312 (n27218, \a[62] , n_23478);
  not g50313 (n_23479, n27218);
  and g50314 (n27219, \a[62] , n_23479);
  and g50315 (n27220, n_23478, n_23479);
  not g50316 (n_23480, n27219);
  not g50317 (n_23481, n27220);
  and g50318 (n27221, n_23480, n_23481);
  not g50319 (n_23482, n27221);
  and g50320 (n27222, n27210, n_23482);
  not g50321 (n_23483, n27222);
  and g50322 (n27223, n27210, n_23483);
  and g50323 (n27224, n_23482, n_23483);
  not g50324 (n_23484, n27223);
  not g50325 (n_23485, n27224);
  and g50326 (n27225, n_23484, n_23485);
  not g50327 (n_23486, n27163);
  not g50328 (n_23487, n27225);
  and g50329 (n27226, n_23486, n_23487);
  and g50330 (n27227, n27163, n27225);
  not g50331 (n_23488, n27226);
  not g50332 (n_23489, n27227);
  and g50333 (n27228, n_23488, n_23489);
  not g50334 (n_23490, n27201);
  and g50335 (n27229, n_23490, n27228);
  not g50336 (n_23491, n27229);
  and g50337 (n27230, n_23490, n_23491);
  and g50338 (n27231, n27228, n_23491);
  not g50339 (n_23492, n27230);
  not g50340 (n_23493, n27231);
  and g50341 (n27232, n_23492, n_23493);
  not g50342 (n_23494, n27199);
  not g50343 (n_23495, n27232);
  and g50344 (n27233, n_23494, n_23495);
  and g50345 (n27234, n27199, n_23493);
  and g50346 (n27235, n_23492, n27234);
  not g50347 (n_23496, n27233);
  not g50348 (n_23497, n27235);
  and g50349 (\f[123] , n_23496, n_23497);
  and g50350 (n27237, n_23491, n_23496);
  and g50351 (n27238, n_23483, n_23488);
  and g50352 (n27239, \b[60] , n13903);
  and g50353 (n27240, \b[61] , n_11555);
  not g50354 (n_23498, n27239);
  not g50355 (n_23499, n27240);
  and g50356 (n27241, n_23498, n_23499);
  and g50357 (n27242, n_9855, n_23426);
  not g50358 (n_23500, n27242);
  and g50359 (n27243, n_23473, n_23500);
  not g50360 (n_23501, n27243);
  and g50361 (n27244, n27241, n_23501);
  not g50362 (n_23502, n27241);
  and g50363 (n27245, n_23502, n27243);
  not g50364 (n_23503, n27244);
  not g50365 (n_23504, n27245);
  and g50366 (n27246, n_23503, n_23504);
  and g50367 (n27247, \b[62] , n13047);
  and g50368 (n27248, \b[63] , n12663);
  not g50369 (n_23505, n27247);
  not g50370 (n_23506, n27248);
  and g50371 (n27249, n_23505, n_23506);
  and g50372 (n27250, n_12644, n27249);
  and g50373 (n27251, n13800, n27249);
  not g50374 (n_23507, n27250);
  not g50375 (n_23508, n27251);
  and g50376 (n27252, n_23507, n_23508);
  not g50377 (n_23509, n27252);
  and g50378 (n27253, \a[62] , n_23509);
  and g50379 (n27254, n_10843, n27252);
  not g50380 (n_23510, n27253);
  not g50381 (n_23511, n27254);
  and g50382 (n27255, n_23510, n_23511);
  not g50383 (n_23512, n27255);
  and g50384 (n27256, n27246, n_23512);
  not g50385 (n_23513, n27246);
  and g50386 (n27257, n_23513, n27255);
  not g50387 (n_23514, n27256);
  not g50388 (n_23515, n27257);
  and g50389 (n27258, n_23514, n_23515);
  not g50390 (n_23516, n27238);
  and g50391 (n27259, n_23516, n27258);
  not g50392 (n_23517, n27259);
  and g50393 (n27260, n_23516, n_23517);
  and g50394 (n27261, n27258, n_23517);
  not g50395 (n_23518, n27260);
  not g50396 (n_23519, n27261);
  and g50397 (n27262, n_23518, n_23519);
  not g50398 (n_23520, n27237);
  not g50399 (n_23521, n27262);
  and g50400 (n27263, n_23520, n_23521);
  and g50401 (n27264, n27237, n_23519);
  and g50402 (n27265, n_23518, n27264);
  not g50403 (n_23522, n27263);
  not g50404 (n_23523, n27265);
  and g50405 (\f[124] , n_23522, n_23523);
  and g50406 (n27267, n_23517, n_23522);
  and g50407 (n27268, n_23503, n_23514);
  and g50408 (n27269, \b[61] , n13903);
  and g50409 (n27270, \b[62] , n_11555);
  not g50410 (n_23524, n27269);
  not g50411 (n_23525, n27270);
  and g50412 (n27271, n_23524, n_23525);
  not g50413 (n_23526, n27271);
  and g50414 (n27272, n27241, n_23526);
  and g50415 (n27273, n_23502, n27271);
  not g50416 (n_23527, n27272);
  not g50417 (n_23528, n27273);
  and g50418 (n27274, n_23527, n_23528);
  and g50419 (n27275, \b[63] , n13047);
  not g50420 (n_23529, n27275);
  and g50421 (n27276, n_12644, n_23529);
  and g50422 (n27277, n_11840, n_23529);
  not g50423 (n_23530, n27276);
  not g50424 (n_23531, n27277);
  and g50425 (n27278, n_23530, n_23531);
  not g50426 (n_23532, n27278);
  and g50427 (n27279, \a[62] , n_23532);
  and g50428 (n27280, n_10843, n27278);
  not g50429 (n_23533, n27279);
  not g50430 (n_23534, n27280);
  and g50431 (n27281, n_23533, n_23534);
  not g50432 (n_23535, n27281);
  and g50433 (n27282, n27274, n_23535);
  not g50434 (n_23536, n27274);
  and g50435 (n27283, n_23536, n27281);
  not g50436 (n_23537, n27282);
  not g50437 (n_23538, n27283);
  and g50438 (n27284, n_23537, n_23538);
  not g50439 (n_23539, n27268);
  and g50440 (n27285, n_23539, n27284);
  not g50441 (n_23540, n27285);
  and g50442 (n27286, n_23539, n_23540);
  and g50443 (n27287, n27284, n_23540);
  not g50444 (n_23541, n27286);
  not g50445 (n_23542, n27287);
  and g50446 (n27288, n_23541, n_23542);
  not g50447 (n_23543, n27267);
  not g50448 (n_23544, n27288);
  and g50449 (n27289, n_23543, n_23544);
  and g50450 (n27290, n27267, n_23542);
  and g50451 (n27291, n_23541, n27290);
  not g50452 (n_23545, n27289);
  not g50453 (n_23546, n27291);
  and g50454 (\f[125] , n_23545, n_23546);
  and g50455 (n27293, n_23540, n_23545);
  and g50456 (n27294, n_23527, n_23537);
  and g50457 (n27295, \b[62] , n13903);
  and g50458 (n27296, \b[63] , n_11555);
  not g50459 (n_23547, n27295);
  not g50460 (n_23548, n27296);
  and g50461 (n27297, n_23547, n_23548);
  not g50462 (n_23549, n27297);
  and g50463 (n27298, n_10843, n_23549);
  and g50464 (n27299, \a[62] , n27297);
  not g50465 (n_23550, n27298);
  not g50466 (n_23551, n27299);
  and g50467 (n27300, n_23550, n_23551);
  and g50468 (n27301, n_23502, n27300);
  not g50469 (n_23552, n27300);
  and g50470 (n27302, n27241, n_23552);
  not g50471 (n_23553, n27301);
  not g50472 (n_23554, n27302);
  and g50473 (n27303, n_23553, n_23554);
  not g50474 (n_23555, n27294);
  and g50475 (n27304, n_23555, n27303);
  not g50476 (n_23556, n27303);
  and g50477 (n27305, n27294, n_23556);
  not g50478 (n_23557, n27304);
  not g50479 (n_23558, n27305);
  and g50480 (n27306, n_23557, n_23558);
  not g50481 (n_23559, n27293);
  and g50482 (n27307, n_23559, n27306);
  not g50483 (n_23560, n27306);
  and g50484 (n27308, n27293, n_23560);
  not g50485 (n_23561, n27307);
  not g50486 (n_23562, n27308);
  and g50487 (\f[126] , n_23561, n_23562);
  and g50488 (n27310, n_23550, n_23553);
  and g50489 (n27311, \b[63] , n13903);
  not g50490 (n_23563, n27310);
  and g50491 (n27312, n_23563, n27311);
  not g50492 (n_23564, n27311);
  and g50493 (n27313, n27310, n_23564);
  not g50494 (n_23565, n27312);
  not g50495 (n_23566, n27313);
  and g50496 (n27314, n_23565, n_23566);
  and g50497 (n27315, n_23557, n_23561);
  and g50498 (n27316, n27314, n27315);
  not g50499 (n_23567, n27314);
  not g50500 (n_23568, n27315);
  and g50501 (n27317, n_23567, n_23568);
  not g50502 (n_23569, n27316);
  not g50503 (n_23570, n27317);
  and g50504 (\f[127] , n_23569, n_23570);
  nor g50505 (n298, n282, n285, n286, n297);
  nor g50506 (n320, n306, n307, n308, n319);
  nor g50507 (n348, n335, n336, n337, n347);
  nor g50508 (n396, n383, n384, n385, n395);
  nor g50509 (n461, n448, n449, n450, n460);
  nor g50510 (n440, n434, n435, n436, n439);
  nor g50511 (n486, n473, n474, n475, n485);
  nor g50512 (n497, n491, n492, n493, n496);
  nor g50513 (n587, n574, n575, n576, n586);
  nor g50514 (n561, n555, n556, n557, n560);
  nor g50515 (n547, n539, n542, n543, n546);
  nor g50516 (n653, n640, n641, n642, n652);
  nor g50517 (n606, n600, n601, n602, n605);
  nor g50518 (n624, n618, n619, n620, n623);
  nor g50519 (n740, n727, n728, n729, n739);
  nor g50520 (n673, n667, n668, n669, n672);
  nor g50521 (n686, n680, n681, n682, n685);
  nor g50522 (n820, n807, n808, n809, n819);
  nor g50523 (n759, n753, n754, n755, n758);
  nor g50524 (n787, n781, n782, n783, n786);
  nor g50525 (n773, n765, n768, n769, n772);
  nor g50526 (n844, n831, n832, n833, n843);
  nor g50527 (n895, n889, n890, n891, n894);
  nor g50528 (n855, n849, n850, n851, n854);
  nor g50529 (n873, n867, n868, n869, n872);
  nor g50530 (n1010, n997, n998, n999, n1009);
  nor g50531 (n984, n978, n979, n980, n983);
  nor g50532 (n924, n918, n919, n920, n923);
  nor g50533 (n937, n931, n932, n933, n936);
  nor g50534 (n1036, n1023, n1024, n1025, n1035);
  nor g50535 (n1047, n1041, n1042, n1043, n1046);
  nor g50536 (n1095, n1089, n1090, n1091, n1094);
  nor g50537 (n1076, n1070, n1071, n1072, n1075);
  nor g50538 (n1062, n1054, n1057, n1058, n1061);
  nor g50539 (n1133, n1120, n1121, n1122, n1132);
  nor g50540 (n1145, n1139, n1140, n1141, n1144);
  nor g50541 (n1157, n1151, n1152, n1153, n1156);
  nor g50542 (n1168, n1162, n1163, n1164, n1167);
  nor g50543 (n1186, n1180, n1181, n1182, n1185);
  nor g50544 (n1239, n1226, n1227, n1228, n1238);
  nor g50545 (n1251, n1245, n1246, n1247, n1250);
  nor g50546 (n1263, n1257, n1258, n1259, n1262);
  nor g50547 (n1275, n1269, n1270, n1271, n1274);
  nor g50548 (n1288, n1282, n1283, n1284, n1287);
  nor g50549 (n1358, n1345, n1346, n1347, n1357);
  nor g50550 (n1370, n1364, n1365, n1366, n1369);
  nor g50551 (n1382, n1376, n1377, n1378, n1381);
  nor g50552 (n1430, n1424, n1425, n1426, n1429);
  nor g50553 (n1411, n1405, n1406, n1407, n1410);
  nor g50554 (n1397, n1389, n1392, n1393, n1396);
  nor g50555 (n1568, n1555, n1556, n1557, n1567);
  nor g50556 (n1469, n1463, n1464, n1465, n1468);
  nor g50557 (n1481, n1475, n1476, n1477, n1480);
  nor g50558 (n1532, n1526, n1527, n1528, n1531);
  nor g50559 (n1493, n1487, n1488, n1489, n1492);
  nor g50560 (n1511, n1505, n1506, n1507, n1510);
  nor g50561 (n1710, n1697, n1698, n1699, n1709);
  nor g50562 (n1587, n1581, n1582, n1583, n1586);
  nor g50563 (n1677, n1671, n1672, n1673, n1676);
  nor g50564 (n1658, n1652, n1653, n1654, n1657);
  nor g50565 (n1600, n1594, n1595, n1596, n1599);
  nor g50566 (n1613, n1607, n1608, n1609, n1612);
  nor g50567 (n1848, n1835, n1836, n1837, n1847);
  nor g50568 (n1730, n1724, n1725, n1726, n1729);
  nor g50569 (n1741, n1735, n1736, n1737, n1740);
  nor g50570 (n1753, n1747, n1748, n1749, n1752);
  nor g50571 (n1802, n1796, n1797, n1798, n1801);
  nor g50572 (n1783, n1777, n1778, n1779, n1782);
  nor g50573 (n1769, n1761, n1764, n1765, n1768);
  nor g50574 (n1986, n1973, n1974, n1975, n1985);
  nor g50575 (n1960, n1954, n1955, n1956, n1959);
  nor g50576 (n1868, n1862, n1863, n1864, n1867);
  nor g50577 (n1880, n1874, n1875, n1876, n1879);
  nor g50578 (n1931, n1925, n1926, n1927, n1930);
  nor g50579 (n1892, n1886, n1887, n1888, n1891);
  nor g50580 (n1910, n1904, n1905, n1906, n1909);
  nor g50581 (n2147, n2134, n2135, n2136, n2146);
  nor g50582 (n2121, n2115, n2116, n2117, n2120);
  nor g50583 (n2007, n2001, n2002, n2003, n2006);
  nor g50584 (n2098, n2092, n2093, n2094, n2097);
  nor g50585 (n2079, n2073, n2074, n2075, n2078);
  nor g50586 (n2021, n2015, n2016, n2017, n2020);
  nor g50587 (n2034, n2028, n2029, n2030, n2033);
  nor g50588 (n2302, n2289, n2290, n2291, n2301);
  nor g50589 (n2276, n2270, n2271, n2272, n2275);
  nor g50590 (n2165, n2159, n2160, n2161, n2164);
  nor g50591 (n2176, n2170, n2171, n2172, n2175);
  nor g50592 (n2188, n2182, n2183, n2184, n2187);
  nor g50593 (n2237, n2231, n2232, n2233, n2236);
  nor g50594 (n2218, n2212, n2213, n2214, n2217);
  nor g50595 (n2204, n2196, n2199, n2200, n2203);
  nor g50596 (n2460, n2447, n2448, n2449, n2459);
  nor g50597 (n2322, n2316, n2317, n2318, n2321);
  nor g50598 (n2428, n2422, n2423, n2424, n2427);
  nor g50599 (n2334, n2328, n2329, n2330, n2333);
  nor g50600 (n2346, n2340, n2341, n2342, n2345);
  nor g50601 (n2397, n2391, n2392, n2393, n2396);
  nor g50602 (n2358, n2352, n2353, n2354, n2357);
  nor g50603 (n2376, n2370, n2371, n2372, n2375);
  nor g50604 (n2487, n2474, n2475, n2476, n2486);
  nor g50605 (n2635, n2629, n2630, n2631, n2634);
  nor g50606 (n2615, n2609, n2610, n2611, n2614);
  nor g50607 (n2499, n2493, n2494, n2495, n2498);
  nor g50608 (n2589, n2583, n2584, n2585, n2588);
  nor g50609 (n2570, n2564, n2565, n2566, n2569);
  nor g50610 (n2512, n2506, n2507, n2508, n2511);
  nor g50611 (n2525, n2519, n2520, n2521, n2524);
  nor g50612 (n2815, n2802, n2803, n2804, n2814);
  nor g50613 (n2790, n2784, n2785, n2786, n2789);
  nor g50614 (n2771, n2765, n2766, n2767, n2770);
  nor g50615 (n2754, n2748, n2749, n2750, n2753);
  nor g50616 (n2663, n2657, n2658, n2659, n2662);
  nor g50617 (n2675, n2669, n2670, n2671, n2674);
  nor g50618 (n2724, n2718, n2719, n2720, n2723);
  nor g50619 (n2705, n2699, n2700, n2701, n2704);
  nor g50620 (n2691, n2683, n2686, n2687, n2690);
  nor g50621 (n2992, n2979, n2980, n2981, n2991);
  nor g50622 (n2833, n2827, n2828, n2829, n2832);
  nor g50623 (n2958, n2952, n2953, n2954, n2957);
  nor g50624 (n2939, n2933, n2934, n2935, n2938);
  nor g50625 (n2844, n2838, n2839, n2840, n2843);
  nor g50626 (n2856, n2850, n2851, n2852, n2855);
  nor g50627 (n2907, n2901, n2902, n2903, n2906);
  nor g50628 (n2868, n2862, n2863, n2864, n2867);
  nor g50629 (n2886, n2880, n2881, n2882, n2885);
  nor g50630 (n3191, n3178, n3179, n3180, n3190);
  nor g50631 (n3010, n3004, n3005, n3006, n3009);
  nor g50632 (n3158, n3152, n3153, n3154, n3157);
  nor g50633 (n3139, n3133, n3134, n3135, n3138);
  nor g50634 (n3120, n3114, n3115, n3116, n3119);
  nor g50635 (n3100, n3094, n3095, n3096, n3099);
  nor g50636 (n3081, n3075, n3076, n3077, n3080);
  nor g50637 (n3023, n3017, n3018, n3019, n3022);
  nor g50638 (n3036, n3030, n3031, n3032, n3035);
  nor g50639 (n3385, n3372, n3373, n3374, n3384);
  nor g50640 (n3209, n3203, n3204, n3205, n3208);
  nor g50641 (n3351, n3345, n3346, n3347, n3350);
  nor g50642 (n3332, n3326, n3327, n3328, n3331);
  nor g50643 (n3313, n3307, n3308, n3309, n3312);
  nor g50644 (n3221, n3215, n3216, n3217, n3220);
  nor g50645 (n3233, n3227, n3228, n3229, n3232);
  nor g50646 (n3282, n3276, n3277, n3278, n3281);
  nor g50647 (n3263, n3257, n3258, n3259, n3262);
  nor g50648 (n3249, n3241, n3244, n3245, n3248);
  nor g50649 (n3579, n3566, n3567, n3568, n3578);
  nor g50650 (n3553, n3547, n3548, n3549, n3552);
  nor g50651 (n3536, n3530, n3531, n3532, n3535);
  nor g50652 (n3518, n3512, n3513, n3514, n3517);
  nor g50653 (n3499, n3493, n3494, n3495, n3498);
  nor g50654 (n3405, n3399, n3400, n3401, n3404);
  nor g50655 (n3417, n3411, n3412, n3413, n3416);
  nor g50656 (n3468, n3462, n3463, n3464, n3467);
  nor g50657 (n3429, n3423, n3424, n3425, n3428);
  nor g50658 (n3447, n3441, n3442, n3443, n3446);
  nor g50659 (n3798, n3785, n3786, n3787, n3797);
  nor g50660 (n3772, n3766, n3767, n3768, n3771);
  nor g50661 (n3753, n3747, n3748, n3749, n3752);
  nor g50662 (n3733, n3727, n3728, n3729, n3732);
  nor g50663 (n3714, n3708, n3709, n3710, n3713);
  nor g50664 (n3598, n3592, n3593, n3594, n3597);
  nor g50665 (n3688, n3682, n3683, n3684, n3687);
  nor g50666 (n3669, n3663, n3664, n3665, n3668);
  nor g50667 (n3611, n3605, n3606, n3607, n3610);
  nor g50668 (n3624, n3618, n3619, n3620, n3623);
  nor g50669 (n4015, n4002, n4003, n4004, n4014);
  nor g50670 (n3989, n3983, n3984, n3985, n3988);
  nor g50671 (n3819, n3813, n3814, n3815, n3818);
  nor g50672 (n3964, n3958, n3959, n3960, n3963);
  nor g50673 (n3945, n3939, n3940, n3941, n3944);
  nor g50674 (n3832, n3826, n3827, n3828, n3831);
  nor g50675 (n3920, n3914, n3915, n3916, n3919);
  nor g50676 (n3901, n3895, n3896, n3897, n3900);
  nor g50677 (n3882, n3876, n3877, n3878, n3881);
  nor g50678 (n3863, n3857, n3858, n3859, n3862);
  nor g50679 (n3849, n3841, n3844, n3845, n3848);
  nor g50680 (n4225, n4212, n4213, n4214, n4224);
  nor g50681 (n4200, n4194, n4195, n4196, n4199);
  nor g50682 (n4034, n4028, n4029, n4030, n4033);
  nor g50683 (n4175, n4169, n4170, n4171, n4174);
  nor g50684 (n4157, n4151, n4152, n4153, n4156);
  nor g50685 (n4140, n4134, n4135, n4136, n4139);
  nor g50686 (n4048, n4042, n4043, n4044, n4047);
  nor g50687 (n4116, n4110, n4111, n4112, n4115);
  nor g50688 (n4099, n4093, n4094, n4095, n4098);
  nor g50689 (n4060, n4054, n4055, n4056, n4059);
  nor g50690 (n4078, n4072, n4073, n4074, n4077);
  nor g50691 (n4468, n4455, n4456, n4457, n4467);
  nor g50692 (n4442, n4436, n4437, n4438, n4441);
  nor g50693 (n4423, n4417, n4418, n4419, n4422);
  nor g50694 (n4404, n4398, n4399, n4400, n4403);
  nor g50695 (n4384, n4378, n4379, n4380, n4383);
  nor g50696 (n4365, n4359, n4360, n4361, n4364);
  nor g50697 (n4345, n4339, n4340, n4341, n4344);
  nor g50698 (n4326, n4320, n4321, n4322, n4325);
  nor g50699 (n4247, n4241, n4242, n4243, n4246);
  nor g50700 (n4260, n4254, n4255, n4256, n4259);
  nor g50701 (n4273, n4267, n4268, n4269, n4272);
  nor g50702 (n4698, n4685, n4686, n4687, n4697);
  nor g50703 (n4672, n4666, n4667, n4668, n4671);
  nor g50704 (n4487, n4481, n4482, n4483, n4486);
  nor g50705 (n4498, n4492, n4493, n4494, n4497);
  nor g50706 (n4641, n4635, n4636, n4637, n4640);
  nor g50707 (n4622, n4616, n4617, n4618, n4621);
  nor g50708 (n4511, n4505, n4506, n4507, n4510);
  nor g50709 (n4597, n4591, n4592, n4593, n4596);
  nor g50710 (n4523, n4517, n4518, n4519, n4522);
  nor g50711 (n4571, n4565, n4566, n4567, n4570);
  nor g50712 (n4552, n4546, n4547, n4548, n4551);
  nor g50713 (n4538, n4530, n4533, n4534, n4537);
  nor g50714 (n4924, n4911, n4912, n4913, n4923);
  nor g50715 (n4715, n4709, n4710, n4711, n4714);
  nor g50716 (n4894, n4888, n4889, n4890, n4893);
  nor g50717 (n4728, n4722, n4723, n4724, n4727);
  nor g50718 (n4870, n4864, n4865, n4866, n4869);
  nor g50719 (n4852, n4846, n4847, n4848, n4851);
  nor g50720 (n4835, n4829, n4830, n4831, n4834);
  nor g50721 (n4742, n4736, n4737, n4738, n4741);
  nor g50722 (n4810, n4804, n4805, n4806, n4809);
  nor g50723 (n4793, n4787, n4788, n4789, n4792);
  nor g50724 (n4754, n4748, n4749, n4750, n4753);
  nor g50725 (n4772, n4766, n4767, n4768, n4771);
  nor g50726 (n5183, n5170, n5171, n5172, n5182);
  nor g50727 (n4945, n4939, n4940, n4941, n4944);
  nor g50728 (n4957, n4951, n4952, n4953, n4956);
  nor g50729 (n5145, n5139, n5140, n5141, n5144);
  nor g50730 (n5126, n5120, n5121, n5122, n5125);
  nor g50731 (n5106, n5100, n5101, n5102, n5105);
  nor g50732 (n5087, n5081, n5082, n5083, n5086);
  nor g50733 (n4971, n4965, n4966, n4967, n4970);
  nor g50734 (n4983, n4977, n4978, n4979, n4982);
  nor g50735 (n4995, n4989, n4990, n4991, n4994);
  nor g50736 (n5008, n5002, n5003, n5004, n5007);
  nor g50737 (n5021, n5015, n5016, n5017, n5020);
  nor g50738 (n5207, n5194, n5195, n5196, n5206);
  nor g50739 (n5219, n5213, n5214, n5215, n5218);
  nor g50740 (n5231, n5225, n5226, n5227, n5230);
  nor g50741 (n5243, n5237, n5238, n5239, n5242);
  nor g50742 (n5403, n5397, n5398, n5399, n5402);
  nor g50743 (n5384, n5378, n5379, n5380, n5383);
  nor g50744 (n5365, n5359, n5360, n5361, n5364);
  nor g50745 (n5255, n5249, n5250, n5251, n5254);
  nor g50746 (n5340, n5334, n5335, n5336, n5339);
  nor g50747 (n5268, n5262, n5263, n5264, n5267);
  nor g50748 (n5315, n5309, n5310, n5311, n5314);
  nor g50749 (n5297, n5291, n5292, n5293, n5296);
  nor g50750 (n5283, n5275, n5278, n5279, n5282);
  nor g50751 (n5453, n5440, n5441, n5442, n5452);
  nor g50752 (n5672, n5666, n5667, n5668, n5671);
  nor g50753 (n5466, n5460, n5461, n5462, n5465);
  nor g50754 (n5648, n5642, n5643, n5644, n5647);
  nor g50755 (n5479, n5473, n5474, n5475, n5478);
  nor g50756 (n5624, n5618, n5619, n5620, n5623);
  nor g50757 (n5605, n5599, n5600, n5601, n5604);
  nor g50758 (n5588, n5582, n5583, n5584, n5587);
  nor g50759 (n5492, n5486, n5487, n5488, n5491);
  nor g50760 (n5563, n5557, n5558, n5559, n5562);
  nor g50761 (n5544, n5538, n5539, n5540, n5543);
  nor g50762 (n5503, n5497, n5498, n5499, n5502);
  nor g50763 (n5521, n5515, n5516, n5517, n5520);
  nor g50764 (n5957, n5944, n5945, n5946, n5956);
  nor g50765 (n5699, n5693, n5694, n5695, n5698);
  nor g50766 (n5712, n5706, n5707, n5708, n5711);
  nor g50767 (n5920, n5914, n5915, n5916, n5919);
  nor g50768 (n5726, n5720, n5721, n5722, n5725);
  nor g50769 (n5893, n5887, n5888, n5889, n5892);
  nor g50770 (n5874, n5868, n5869, n5870, n5873);
  nor g50771 (n5855, n5849, n5850, n5851, n5854);
  nor g50772 (n5737, n5731, n5732, n5733, n5736);
  nor g50773 (n5829, n5823, n5824, n5825, n5828);
  nor g50774 (n5810, n5804, n5805, n5806, n5809);
  nor g50775 (n5750, n5744, n5745, n5746, n5749);
  nor g50776 (n5763, n5757, n5758, n5759, n5762);
  nor g50777 (n6221, n6208, n6209, n6210, n6220);
  nor g50778 (n6197, n6191, n6192, n6193, n6196);
  nor g50779 (n5978, n5972, n5973, n5974, n5977);
  nor g50780 (n5990, n5984, n5985, n5986, n5989);
  nor g50781 (n6002, n5996, n5997, n5998, n6001);
  nor g50782 (n6161, n6155, n6156, n6157, n6160);
  nor g50783 (n6142, n6136, n6137, n6138, n6141);
  nor g50784 (n6015, n6009, n6010, n6011, n6014);
  nor g50785 (n6027, n6021, n6022, n6023, n6026);
  nor g50786 (n6039, n6033, n6034, n6035, n6038);
  nor g50787 (n6105, n6099, n6100, n6101, n6104);
  nor g50788 (n6051, n6045, n6046, n6047, n6050);
  nor g50789 (n6079, n6073, n6074, n6075, n6078);
  nor g50790 (n6065, n6057, n6060, n6061, n6064);
  nor g50791 (n6491, n6478, n6479, n6480, n6490);
  nor g50792 (n6239, n6233, n6234, n6235, n6238);
  nor g50793 (n6459, n6453, n6454, n6455, n6458);
  nor g50794 (n6253, n6247, n6248, n6249, n6252);
  nor g50795 (n6435, n6429, n6430, n6431, n6434);
  nor g50796 (n6266, n6260, n6261, n6262, n6265);
  nor g50797 (n6411, n6405, n6406, n6407, n6410);
  nor g50798 (n6277, n6271, n6272, n6273, n6276);
  nor g50799 (n6386, n6380, n6381, n6382, n6385);
  nor g50800 (n6368, n6362, n6363, n6364, n6367);
  nor g50801 (n6291, n6285, n6286, n6287, n6290);
  nor g50802 (n6343, n6337, n6338, n6339, n6342);
  nor g50803 (n6303, n6297, n6298, n6299, n6302);
  nor g50804 (n6321, n6315, n6316, n6317, n6320);
  nor g50805 (n6517, n6504, n6505, n6506, n6516);
  nor g50806 (n6783, n6777, n6778, n6779, n6782);
  nor g50807 (n6764, n6758, n6759, n6760, n6763);
  nor g50808 (n6530, n6524, n6525, n6526, n6529);
  nor g50809 (n6738, n6732, n6733, n6734, n6737);
  nor g50810 (n6544, n6538, n6539, n6540, n6543);
  nor g50811 (n6711, n6705, n6706, n6707, n6710);
  nor g50812 (n6692, n6686, n6687, n6688, n6691);
  nor g50813 (n6673, n6667, n6668, n6669, n6672);
  nor g50814 (n6555, n6549, n6550, n6551, n6554);
  nor g50815 (n6647, n6641, n6642, n6643, n6646);
  nor g50816 (n6628, n6622, n6623, n6624, n6627);
  nor g50817 (n6568, n6562, n6563, n6564, n6567);
  nor g50818 (n6581, n6575, n6576, n6577, n6580);
  nor g50819 (n7074, n7061, n7062, n7063, n7073);
  nor g50820 (n6810, n6804, n6805, n6806, n6809);
  nor g50821 (n7041, n7035, n7036, n7037, n7040);
  nor g50822 (n6821, n6815, n6816, n6817, n6820);
  nor g50823 (n6833, n6827, n6828, n6829, n6832);
  nor g50824 (n6845, n6839, n6840, n6841, n6844);
  nor g50825 (n7004, n6998, n6999, n7000, n7003);
  nor g50826 (n6985, n6979, n6980, n6981, n6984);
  nor g50827 (n6858, n6852, n6853, n6854, n6857);
  nor g50828 (n6870, n6864, n6865, n6866, n6869);
  nor g50829 (n6882, n6876, n6877, n6878, n6881);
  nor g50830 (n6948, n6942, n6943, n6944, n6947);
  nor g50831 (n6894, n6888, n6889, n6890, n6893);
  nor g50832 (n6922, n6916, n6917, n6918, n6921);
  nor g50833 (n6908, n6900, n6903, n6904, n6907);
  nor g50834 (n7363, n7350, n7351, n7352, n7362);
  nor g50835 (n7337, n7331, n7332, n7333, n7336);
  nor g50836 (n7318, n7312, n7313, n7314, n7317);
  nor g50837 (n7301, n7295, n7296, n7297, n7300);
  nor g50838 (n7095, n7089, n7090, n7091, n7094);
  nor g50839 (n7277, n7271, n7272, n7273, n7276);
  nor g50840 (n7108, n7102, n7103, n7104, n7107);
  nor g50841 (n7253, n7247, n7248, n7249, n7252);
  nor g50842 (n7119, n7113, n7114, n7115, n7118);
  nor g50843 (n7228, n7222, n7223, n7224, n7227);
  nor g50844 (n7210, n7204, n7205, n7206, n7209);
  nor g50845 (n7133, n7127, n7128, n7129, n7132);
  nor g50846 (n7185, n7179, n7180, n7181, n7184);
  nor g50847 (n7145, n7139, n7140, n7141, n7144);
  nor g50848 (n7163, n7157, n7158, n7159, n7162);
  nor g50849 (n7679, n7666, n7667, n7668, n7678);
  nor g50850 (n7653, n7647, n7648, n7649, n7652);
  nor g50851 (n7634, n7628, n7629, n7630, n7633);
  nor g50852 (n7615, n7609, n7610, n7611, n7614);
  nor g50853 (n7381, n7375, n7376, n7377, n7380);
  nor g50854 (n7589, n7583, n7584, n7585, n7588);
  nor g50855 (n7395, n7389, n7390, n7391, n7394);
  nor g50856 (n7562, n7556, n7557, n7558, n7561);
  nor g50857 (n7543, n7537, n7538, n7539, n7542);
  nor g50858 (n7524, n7518, n7519, n7520, n7523);
  nor g50859 (n7406, n7400, n7401, n7402, n7405);
  nor g50860 (n7498, n7492, n7493, n7494, n7497);
  nor g50861 (n7479, n7473, n7474, n7475, n7478);
  nor g50862 (n7419, n7413, n7414, n7415, n7418);
  nor g50863 (n7432, n7426, n7427, n7428, n7431);
  nor g50864 (n7705, n7692, n7693, n7694, n7704);
  nor g50865 (n7978, n7972, n7973, n7974, n7977);
  nor g50866 (n7959, n7953, n7954, n7955, n7958);
  nor g50867 (n7940, n7934, n7935, n7936, n7939);
  nor g50868 (n7717, n7711, n7712, n7713, n7716);
  nor g50869 (n7729, n7723, n7724, n7725, n7728);
  nor g50870 (n7741, n7735, n7736, n7737, n7740);
  nor g50871 (n7903, n7897, n7898, n7899, n7902);
  nor g50872 (n7884, n7878, n7879, n7880, n7883);
  nor g50873 (n7865, n7859, n7860, n7861, n7864);
  nor g50874 (n7755, n7749, n7750, n7751, n7754);
  nor g50875 (n7767, n7761, n7762, n7763, n7766);
  nor g50876 (n7833, n7827, n7828, n7829, n7832);
  nor g50877 (n7779, n7773, n7774, n7775, n7778);
  nor g50878 (n7807, n7801, n7802, n7803, n7806);
  nor g50879 (n7793, n7785, n7788, n7789, n7792);
  nor g50880 (n8011, n7998, n7999, n8000, n8010);
  nor g50881 (n8285, n8279, n8280, n8281, n8284);
  nor g50882 (n8267, n8261, n8262, n8263, n8266);
  nor g50883 (n8248, n8242, n8243, n8244, n8247);
  nor g50884 (n8231, n8225, n8226, n8227, n8230);
  nor g50885 (n8025, n8019, n8020, n8021, n8024);
  nor g50886 (n8207, n8201, n8202, n8203, n8206);
  nor g50887 (n8038, n8032, n8033, n8034, n8037);
  nor g50888 (n8183, n8177, n8178, n8179, n8182);
  nor g50889 (n8164, n8158, n8159, n8160, n8163);
  nor g50890 (n8145, n8139, n8140, n8141, n8144);
  nor g50891 (n8050, n8044, n8045, n8046, n8049);
  nor g50892 (n8062, n8056, n8057, n8058, n8061);
  nor g50893 (n8114, n8108, n8109, n8110, n8113);
  nor g50894 (n8074, n8068, n8069, n8070, n8073);
  nor g50895 (n8092, n8086, n8087, n8088, n8091);
  nor g50896 (n8627, n8614, n8615, n8616, n8626);
  nor g50897 (n8601, n8595, n8596, n8597, n8600);
  nor g50898 (n8581, n8575, n8576, n8577, n8580);
  nor g50899 (n8562, n8556, n8557, n8558, n8561);
  nor g50900 (n8543, n8537, n8538, n8539, n8542);
  nor g50901 (n8523, n8517, n8518, n8519, n8522);
  nor g50902 (n8504, n8498, n8499, n8500, n8503);
  nor g50903 (n8311, n8305, n8306, n8307, n8310);
  nor g50904 (n8477, n8471, n8472, n8473, n8476);
  nor g50905 (n8458, n8452, n8453, n8454, n8457);
  nor g50906 (n8439, n8433, n8434, n8435, n8438);
  nor g50907 (n8322, n8316, n8317, n8318, n8321);
  nor g50908 (n8414, n8408, n8409, n8410, n8413);
  nor g50909 (n8395, n8389, n8390, n8391, n8394);
  nor g50910 (n8335, n8329, n8330, n8331, n8334);
  nor g50911 (n8348, n8342, n8343, n8344, n8347);
  nor g50912 (n8951, n8938, n8939, n8940, n8950);
  nor g50913 (n8925, n8919, n8920, n8921, n8924);
  nor g50914 (n8906, n8900, n8901, n8902, n8905);
  nor g50915 (n8887, n8881, n8882, n8883, n8886);
  nor g50916 (n8868, n8862, n8863, n8864, n8867);
  nor g50917 (n8645, n8639, n8640, n8641, n8644);
  nor g50918 (n8657, n8651, n8652, n8653, n8656);
  nor g50919 (n8669, n8663, n8664, n8665, n8668);
  nor g50920 (n8831, n8825, n8826, n8827, n8830);
  nor g50921 (n8812, n8806, n8807, n8808, n8811);
  nor g50922 (n8793, n8787, n8788, n8789, n8792);
  nor g50923 (n8683, n8677, n8678, n8679, n8682);
  nor g50924 (n8695, n8689, n8690, n8691, n8694);
  nor g50925 (n8761, n8755, n8756, n8757, n8760);
  nor g50926 (n8707, n8701, n8702, n8703, n8706);
  nor g50927 (n8735, n8729, n8730, n8731, n8734);
  nor g50928 (n8721, n8713, n8716, n8717, n8720);
  nor g50929 (n8978, n8965, n8966, n8967, n8977);
  nor g50930 (n9269, n9263, n9264, n9265, n9268);
  nor g50931 (n8990, n8984, n8985, n8986, n8989);
  nor g50932 (n9244, n9238, n9239, n9240, n9243);
  nor g50933 (n9225, n9219, n9220, n9221, n9224);
  nor g50934 (n9208, n9202, n9203, n9204, n9207);
  nor g50935 (n9003, n8997, n8998, n8999, n9002);
  nor g50936 (n9184, n9178, n9179, n9180, n9183);
  nor g50937 (n9016, n9010, n9011, n9012, n9015);
  nor g50938 (n9160, n9154, n9155, n9156, n9159);
  nor g50939 (n9141, n9135, n9136, n9137, n9140);
  nor g50940 (n9028, n9022, n9023, n9024, n9027);
  nor g50941 (n9040, n9034, n9035, n9036, n9039);
  nor g50942 (n9052, n9046, n9047, n9048, n9051);
  nor g50943 (n9104, n9098, n9099, n9100, n9103);
  nor g50944 (n9064, n9058, n9059, n9060, n9063);
  nor g50945 (n9082, n9076, n9077, n9078, n9081);
  nor g50946 (n9630, n9617, n9618, n9619, n9629);
  nor g50947 (n9605, n9599, n9600, n9601, n9604);
  nor g50948 (n9585, n9579, n9580, n9581, n9584);
  nor g50949 (n9566, n9560, n9561, n9562, n9565);
  nor g50950 (n9547, n9541, n9542, n9543, n9546);
  nor g50951 (n9528, n9522, n9523, n9524, n9527);
  nor g50952 (n9508, n9502, n9503, n9504, n9507);
  nor g50953 (n9489, n9483, n9484, n9485, n9488);
  nor g50954 (n9472, n9466, n9467, n9468, n9471);
  nor g50955 (n9454, n9448, n9449, n9450, n9453);
  nor g50956 (n9435, n9429, n9430, n9431, n9434);
  nor g50957 (n9416, n9410, n9411, n9412, n9415);
  nor g50958 (n9299, n9293, n9294, n9295, n9298);
  nor g50959 (n9391, n9385, n9386, n9387, n9390);
  nor g50960 (n9372, n9366, n9367, n9368, n9371);
  nor g50961 (n9312, n9306, n9307, n9308, n9311);
  nor g50962 (n9325, n9319, n9320, n9321, n9324);
  nor g50963 (n9974, n9961, n9962, n9963, n9973);
  nor g50964 (n9948, n9942, n9943, n9944, n9947);
  nor g50965 (n9929, n9923, n9924, n9925, n9928);
  nor g50966 (n9910, n9904, n9905, n9906, n9909);
  nor g50967 (n9891, n9885, n9886, n9887, n9890);
  nor g50968 (n9872, n9866, n9867, n9868, n9871);
  nor g50969 (n9650, n9644, n9645, n9646, n9649);
  nor g50970 (n9662, n9656, n9657, n9658, n9661);
  nor g50971 (n9674, n9668, n9669, n9670, n9673);
  nor g50972 (n9835, n9829, n9830, n9831, n9834);
  nor g50973 (n9688, n9682, n9683, n9684, n9687);
  nor g50974 (n9809, n9803, n9804, n9805, n9808);
  nor g50975 (n9700, n9694, n9695, n9696, n9699);
  nor g50976 (n9712, n9706, n9707, n9708, n9711);
  nor g50977 (n9723, n9717, n9718, n9719, n9722);
  nor g50978 (n9771, n9765, n9766, n9767, n9770);
  nor g50979 (n9752, n9746, n9747, n9748, n9751);
  nor g50980 (n9738, n9730, n9733, n9734, n9737);
  nor g50981 (n10000, n9987, n9988, n9989, n9999);
  nor g50982 (n10312, n10306, n10307, n10308, n10311);
  nor g50983 (n10293, n10287, n10288, n10289, n10292);
  nor g50984 (n10011, n10005, n10006, n10007, n10010);
  nor g50985 (n10268, n10262, n10263, n10264, n10267);
  nor g50986 (n10249, n10243, n10244, n10245, n10248);
  nor g50987 (n10232, n10226, n10227, n10228, n10231);
  nor g50988 (n10214, n10208, n10209, n10210, n10213);
  nor g50989 (n10026, n10020, n10021, n10022, n10025);
  nor g50990 (n10038, n10032, n10033, n10034, n10037);
  nor g50991 (n10050, n10044, n10045, n10046, n10049);
  nor g50992 (n10062, n10056, n10057, n10058, n10061);
  nor g50993 (n10074, n10068, n10069, n10070, n10073);
  nor g50994 (n10086, n10080, n10081, n10082, n10085);
  nor g50995 (n10098, n10092, n10093, n10094, n10097);
  nor g50996 (n10110, n10104, n10105, n10106, n10109);
  nor g50997 (n10121, n10115, n10116, n10117, n10120);
  nor g50998 (n10139, n10133, n10134, n10135, n10138);
  nor g50999 (n10686, n10673, n10674, n10675, n10685);
  nor g51000 (n10337, n10331, n10332, n10333, n10336);
  nor g51001 (n10349, n10343, n10344, n10345, n10348);
  nor g51002 (n10649, n10643, n10644, n10645, n10648);
  nor g51003 (n10630, n10624, n10625, n10626, n10629);
  nor g51004 (n10611, n10605, n10606, n10607, n10610);
  nor g51005 (n10592, n10586, n10587, n10588, n10591);
  nor g51006 (n10572, n10566, n10567, n10568, n10571);
  nor g51007 (n10553, n10547, n10548, n10549, n10552);
  nor g51008 (n10534, n10528, n10529, n10530, n10533);
  nor g51009 (n10515, n10509, n10510, n10511, n10514);
  nor g51010 (n10496, n10490, n10491, n10492, n10495);
  nor g51011 (n10477, n10471, n10472, n10473, n10476);
  nor g51012 (n10363, n10357, n10358, n10359, n10362);
  nor g51013 (n10375, n10369, n10370, n10371, n10374);
  nor g51014 (n10387, n10381, n10382, n10383, n10386);
  nor g51015 (n10399, n10393, n10394, n10395, n10398);
  nor g51016 (n10412, n10406, n10407, n10408, n10411);
  nor g51017 (n10710, n10697, n10698, n10699, n10709);
  nor g51018 (n11041, n11035, n11036, n11037, n11040);
  nor g51019 (n10724, n10718, n10719, n10720, n10723);
  nor g51020 (n11015, n11009, n11010, n11011, n11014);
  nor g51021 (n10996, n10990, n10991, n10992, n10995);
  nor g51022 (n10977, n10971, n10972, n10973, n10976);
  nor g51023 (n10958, n10952, n10953, n10954, n10957);
  nor g51024 (n10736, n10730, n10731, n10732, n10735);
  nor g51025 (n10748, n10742, n10743, n10744, n10747);
  nor g51026 (n10927, n10921, n10922, n10923, n10926);
  nor g51027 (n10908, n10902, n10903, n10904, n10907);
  nor g51028 (n10891, n10885, n10886, n10887, n10890);
  nor g51029 (n10873, n10867, n10868, n10869, n10872);
  nor g51030 (n10763, n10757, n10758, n10759, n10762);
  nor g51031 (n10775, n10769, n10770, n10771, n10774);
  nor g51032 (n10787, n10781, n10782, n10783, n10786);
  nor g51033 (n10835, n10829, n10830, n10831, n10834);
  nor g51034 (n10816, n10810, n10811, n10812, n10815);
  nor g51035 (n10802, n10794, n10797, n10798, n10801);
  nor g51036 (n11412, n11399, n11400, n11401, n11411);
  nor g51037 (n11067, n11061, n11062, n11063, n11066);
  nor g51038 (n11079, n11073, n11074, n11075, n11078);
  nor g51039 (n11091, n11085, n11086, n11087, n11090);
  nor g51040 (n11102, n11096, n11097, n11098, n11101);
  nor g51041 (n11356, n11350, n11351, n11352, n11355);
  nor g51042 (n11337, n11331, n11332, n11333, n11336);
  nor g51043 (n11320, n11314, n11315, n11316, n11319);
  nor g51044 (n11302, n11296, n11297, n11298, n11301);
  nor g51045 (n11117, n11111, n11112, n11113, n11116);
  nor g51046 (n11279, n11273, n11274, n11275, n11278);
  nor g51047 (n11260, n11254, n11255, n11256, n11259);
  nor g51048 (n11130, n11124, n11125, n11126, n11129);
  nor g51049 (n11142, n11136, n11137, n11138, n11141);
  nor g51050 (n11154, n11148, n11149, n11150, n11153);
  nor g51051 (n11166, n11160, n11161, n11162, n11165);
  nor g51052 (n11217, n11211, n11212, n11213, n11216);
  nor g51053 (n11178, n11172, n11173, n11174, n11177);
  nor g51054 (n11196, n11190, n11191, n11192, n11195);
  nor g51055 (n11438, n11425, n11426, n11427, n11437);
  nor g51056 (n11450, n11444, n11445, n11446, n11449);
  nor g51057 (n11462, n11456, n11457, n11458, n11461);
  nor g51058 (n11474, n11468, n11469, n11470, n11473);
  nor g51059 (n11777, n11771, n11772, n11773, n11776);
  nor g51060 (n11758, n11752, n11753, n11754, n11757);
  nor g51061 (n11739, n11733, n11734, n11735, n11738);
  nor g51062 (n11720, n11714, n11715, n11716, n11719);
  nor g51063 (n11700, n11694, n11695, n11696, n11699);
  nor g51064 (n11683, n11677, n11678, n11679, n11682);
  nor g51065 (n11665, n11659, n11660, n11661, n11664);
  nor g51066 (n11646, n11640, n11641, n11642, n11645);
  nor g51067 (n11627, n11621, n11622, n11623, n11626);
  nor g51068 (n11608, n11602, n11603, n11604, n11607);
  nor g51069 (n11589, n11583, n11584, n11585, n11588);
  nor g51070 (n11570, n11564, n11565, n11566, n11569);
  nor g51071 (n11491, n11485, n11486, n11487, n11490);
  nor g51072 (n11504, n11498, n11499, n11500, n11503);
  nor g51073 (n11517, n11511, n11512, n11513, n11516);
  nor g51074 (n12181, n12168, n12169, n12170, n12180);
  nor g51075 (n12159, n12153, n12154, n12155, n12158);
  nor g51076 (n11823, n11817, n11818, n11819, n11822);
  nor g51077 (n11835, n11829, n11830, n11831, n11834);
  nor g51078 (n12127, n12121, n12122, n12123, n12126);
  nor g51079 (n12109, n12103, n12104, n12105, n12108);
  nor g51080 (n12090, n12084, n12085, n12086, n12089);
  nor g51081 (n12071, n12065, n12066, n12067, n12070);
  nor g51082 (n11848, n11842, n11843, n11844, n11847);
  nor g51083 (n12046, n12040, n12041, n12042, n12045);
  nor g51084 (n12027, n12021, n12022, n12023, n12026);
  nor g51085 (n12008, n12002, n12003, n12004, n12007);
  nor g51086 (n11991, n11985, n11986, n11987, n11990);
  nor g51087 (n11973, n11967, n11968, n11969, n11972);
  nor g51088 (n11864, n11858, n11859, n11860, n11863);
  nor g51089 (n11875, n11869, n11870, n11871, n11874);
  nor g51090 (n11887, n11881, n11882, n11883, n11886);
  nor g51091 (n11935, n11929, n11930, n11931, n11934);
  nor g51092 (n11916, n11910, n11911, n11912, n11915);
  nor g51093 (n11902, n11894, n11897, n11898, n11901);
  nor g51094 (n12213, n12200, n12201, n12202, n12212);
  nor g51095 (n12224, n12218, n12219, n12220, n12223);
  nor g51096 (n12236, n12230, n12231, n12232, n12235);
  nor g51097 (n12248, n12242, n12243, n12244, n12247);
  nor g51098 (n12260, n12254, n12255, n12256, n12259);
  nor g51099 (n12273, n12267, n12268, n12269, n12272);
  nor g51100 (n12527, n12521, n12522, n12523, n12526);
  nor g51101 (n12508, n12502, n12503, n12504, n12507);
  nor g51102 (n12491, n12485, n12486, n12487, n12490);
  nor g51103 (n12286, n12280, n12281, n12282, n12285);
  nor g51104 (n12467, n12461, n12462, n12463, n12466);
  nor g51105 (n12448, n12442, n12443, n12444, n12447);
  nor g51106 (n12429, n12423, n12424, n12425, n12428);
  nor g51107 (n12299, n12293, n12294, n12295, n12298);
  nor g51108 (n12311, n12305, n12306, n12307, n12310);
  nor g51109 (n12323, n12317, n12318, n12319, n12322);
  nor g51110 (n12335, n12329, n12330, n12331, n12334);
  nor g51111 (n12386, n12380, n12381, n12382, n12385);
  nor g51112 (n12347, n12341, n12342, n12343, n12346);
  nor g51113 (n12365, n12359, n12360, n12361, n12364);
  nor g51114 (n12971, n12958, n12959, n12960, n12970);
  nor g51115 (n12950, n12944, n12945, n12946, n12949);
  nor g51116 (n12586, n12580, n12581, n12582, n12585);
  nor g51117 (n12598, n12592, n12593, n12594, n12597);
  nor g51118 (n12610, n12604, n12605, n12606, n12609);
  nor g51119 (n12913, n12907, n12908, n12909, n12912);
  nor g51120 (n12894, n12888, n12889, n12890, n12893);
  nor g51121 (n12875, n12869, n12870, n12871, n12874);
  nor g51122 (n12856, n12850, n12851, n12852, n12855);
  nor g51123 (n12839, n12833, n12834, n12835, n12838);
  nor g51124 (n12821, n12815, n12816, n12817, n12820);
  nor g51125 (n12802, n12796, n12797, n12798, n12801);
  nor g51126 (n12783, n12777, n12778, n12779, n12782);
  nor g51127 (n12764, n12758, n12759, n12760, n12763);
  nor g51128 (n12745, n12739, n12740, n12741, n12744);
  nor g51129 (n12726, n12720, n12721, n12722, n12725);
  nor g51130 (n12707, n12701, n12702, n12703, n12706);
  nor g51131 (n12628, n12622, n12623, n12624, n12627);
  nor g51132 (n12641, n12635, n12636, n12637, n12640);
  nor g51133 (n12654, n12648, n12649, n12650, n12653);
  nor g51134 (n13372, n13359, n13360, n13361, n13371);
  nor g51135 (n13346, n13340, n13341, n13342, n13345);
  nor g51136 (n13332, n13326, n13327, n13328, n13331);
  nor g51137 (n13315, n13309, n13310, n13311, n13314);
  nor g51138 (n12998, n12992, n12993, n12994, n12997);
  nor g51139 (n13291, n13285, n13286, n13287, n13290);
  nor g51140 (n13273, n13267, n13268, n13269, n13272);
  nor g51141 (n13254, n13248, n13249, n13250, n13253);
  nor g51142 (n13235, n13229, n13230, n13231, n13234);
  nor g51143 (n13216, n13210, n13211, n13212, n13215);
  nor g51144 (n13197, n13191, n13192, n13193, n13196);
  nor g51145 (n13178, n13172, n13173, n13174, n13177);
  nor g51146 (n13159, n13153, n13154, n13155, n13158);
  nor g51147 (n13142, n13136, n13137, n13138, n13141);
  nor g51148 (n13124, n13118, n13119, n13120, n13123);
  nor g51149 (n13015, n13009, n13010, n13011, n13014);
  nor g51150 (n13026, n13020, n13021, n13022, n13025);
  nor g51151 (n13038, n13032, n13033, n13034, n13037);
  nor g51152 (n13086, n13080, n13081, n13082, n13085);
  nor g51153 (n13067, n13061, n13062, n13063, n13066);
  nor g51154 (n13053, n13045, n13048, n13049, n13052);
  nor g51155 (n13773, n13760, n13761, n13762, n13772);
  nor g51156 (n13748, n13742, n13743, n13744, n13747);
  nor g51157 (n13733, n13727, n13728, n13729, n13732);
  nor g51158 (n13714, n13708, n13709, n13710, n13713);
  nor g51159 (n13394, n13388, n13389, n13390, n13393);
  nor g51160 (n13406, n13400, n13401, n13402, n13405);
  nor g51161 (n13419, n13413, n13414, n13415, n13418);
  nor g51162 (n13430, n13424, n13425, n13426, n13429);
  nor g51163 (n13667, n13661, n13662, n13663, n13666);
  nor g51164 (n13650, n13644, n13645, n13646, n13649);
  nor g51165 (n13443, n13437, n13438, n13439, n13442);
  nor g51166 (n13625, n13619, n13620, n13621, n13624);
  nor g51167 (n13606, n13600, n13601, n13602, n13605);
  nor g51168 (n13587, n13581, n13582, n13583, n13586);
  nor g51169 (n13456, n13450, n13451, n13452, n13455);
  nor g51170 (n13564, n13558, n13559, n13560, n13563);
  nor g51171 (n13468, n13462, n13463, n13464, n13467);
  nor g51172 (n13539, n13533, n13534, n13535, n13538);
  nor g51173 (n13481, n13475, n13476, n13477, n13480);
  nor g51174 (n13515, n13509, n13510, n13511, n13514);
  nor g51175 (n13500, n13494, n13495, n13496, n13499);
  nor g51176 (n14174, n14168, n14169, n14170, n14173);
  nor g51177 (n14159, n14153, n14154, n14155, n14158);
  nor g51178 (n13816, n13810, n13811, n13812, n13815);
  nor g51179 (n13828, n13822, n13823, n13824, n13827);
  nor g51180 (n13840, n13834, n13835, n13836, n13839);
  nor g51181 (n13852, n13846, n13847, n13848, n13851);
  nor g51182 (n14114, n14108, n14109, n14110, n14113);
  nor g51183 (n14094, n14088, n14089, n14090, n14093);
  nor g51184 (n14075, n14069, n14070, n14071, n14074);
  nor g51185 (n13864, n13858, n13859, n13860, n13863);
  nor g51186 (n14048, n14042, n14043, n14044, n14047);
  nor g51187 (n14029, n14023, n14024, n14025, n14028);
  nor g51188 (n14010, n14004, n14005, n14006, n14009);
  nor g51189 (n13875, n13869, n13870, n13871, n13874);
  nor g51190 (n13984, n13978, n13979, n13980, n13983);
  nor g51191 (n13886, n13880, n13881, n13882, n13885);
  nor g51192 (n13958, n13952, n13953, n13954, n13957);
  nor g51193 (n13897, n13891, n13892, n13893, n13896);
  nor g51194 (n13932, n13926, n13927, n13928, n13931);
  nor g51195 (n13913, n13907, n13908, n13909, n13912);
  nor g51196 (n14560, n14554, n14555, n14556, n14559);
  nor g51197 (n14541, n14535, n14536, n14537, n14540);
  nor g51198 (n14527, n14521, n14522, n14523, n14526);
  nor g51199 (n14200, n14194, n14195, n14196, n14199);
  nor g51200 (n14502, n14496, n14497, n14498, n14501);
  nor g51201 (n14213, n14207, n14208, n14209, n14212);
  nor g51202 (n14474, n14468, n14469, n14470, n14473);
  nor g51203 (n14455, n14449, n14450, n14451, n14454);
  nor g51204 (n14436, n14430, n14431, n14432, n14435);
  nor g51205 (n14417, n14411, n14412, n14413, n14416);
  nor g51206 (n14398, n14392, n14393, n14394, n14397);
  nor g51207 (n14379, n14373, n14374, n14375, n14378);
  nor g51208 (n14360, n14354, n14355, n14356, n14359);
  nor g51209 (n14343, n14337, n14338, n14339, n14342);
  nor g51210 (n14325, n14319, n14320, n14321, n14324);
  nor g51211 (n14308, n14302, n14303, n14304, n14307);
  nor g51212 (n14230, n14224, n14225, n14226, n14229);
  nor g51213 (n14284, n14278, n14279, n14280, n14283);
  nor g51214 (n14265, n14259, n14260, n14261, n14264);
  nor g51215 (n14246, n14240, n14241, n14242, n14245);
  nor g51216 (n14599, n14593, n14594, n14595, n14598);
  nor g51217 (n14955, n14949, n14950, n14951, n14954);
  nor g51218 (n14614, n14608, n14609, n14610, n14613);
  nor g51219 (n14629, n14623, n14624, n14625, n14628);
  nor g51220 (n14644, n14638, n14639, n14640, n14643);
  nor g51221 (n14659, n14653, n14654, n14655, n14658);
  nor g51222 (n14673, n14667, n14668, n14669, n14672);
  nor g51223 (n14703, n14697, n14698, n14699, n14702);
  nor g51224 (n14870, n14864, n14865, n14866, n14869);
  nor g51225 (n14851, n14845, n14846, n14847, n14850);
  nor g51226 (n14714, n14708, n14709, n14710, n14713);
  nor g51227 (n14824, n14818, n14819, n14820, n14823);
  nor g51228 (n14805, n14799, n14800, n14801, n14804);
  nor g51229 (n14725, n14719, n14720, n14721, n14724);
  nor g51230 (n14779, n14773, n14774, n14775, n14778);
  nor g51231 (n14761, n14755, n14756, n14757, n14760);
  nor g51232 (n14989, n14983, n14984, n14985, n14988);
  nor g51233 (n15294, n15288, n15289, n15290, n15293);
  nor g51234 (n15004, n14998, n14999, n15000, n15003);
  nor g51235 (n15271, n15265, n15266, n15267, n15270);
  nor g51236 (n15020, n15014, n15015, n15016, n15019);
  nor g51237 (n15050, n15044, n15045, n15046, n15049);
  nor g51238 (n15222, n15216, n15217, n15218, n15221);
  nor g51239 (n15203, n15197, n15198, n15199, n15202);
  nor g51240 (n15184, n15178, n15179, n15180, n15183);
  nor g51241 (n15164, n15158, n15159, n15160, n15163);
  nor g51242 (n15145, n15139, n15140, n15141, n15144);
  nor g51243 (n15062, n15056, n15057, n15058, n15061);
  nor g51244 (n15118, n15112, n15113, n15114, n15117);
  nor g51245 (n15099, n15093, n15094, n15095, n15098);
  nor g51246 (n15073, n15067, n15068, n15069, n15072);
  nor g51247 (n15397, n15391, n15392, n15393, n15396);
  nor g51248 (n15412, n15406, n15407, n15408, n15411);
  nor g51249 (n15444, n15438, n15439, n15440, n15443);
  nor g51250 (n15461, n15455, n15456, n15457, n15460);
  nor g51251 (n15476, n15470, n15471, n15472, n15475);
  nor g51252 (n15491, n15485, n15486, n15487, n15490);
  nor g51253 (n15660, n15654, n15655, n15656, n15659);
  nor g51254 (n15641, n15635, n15636, n15637, n15640);
  nor g51255 (n15622, n15616, n15617, n15618, n15621);
  nor g51256 (n15502, n15496, n15497, n15498, n15501);
  nor g51257 (n15596, n15590, n15591, n15592, n15595);
  nor g51258 (n15577, n15571, n15572, n15573, n15576);
  nor g51259 (n15513, n15507, n15508, n15509, n15512);
  nor g51260 (n15550, n15544, n15545, n15546, n15549);
  nor g51261 (n15524, n15518, n15519, n15520, n15523);
  nor g51262 (n15777, n15771, n15772, n15773, n15776);
  nor g51263 (n15792, n15786, n15787, n15788, n15791);
  nor g51264 (n16119, n16113, n16114, n16115, n16118);
  nor g51265 (n15808, n15802, n15803, n15804, n15807);
  nor g51266 (n16095, n16089, n16090, n16091, n16094);
  nor g51267 (n15823, n15817, n15818, n15819, n15822);
  nor g51268 (n15839, n15833, n15834, n15835, n15838);
  nor g51269 (n15854, n15848, n15849, n15850, n15853);
  nor g51270 (n16067, n16061, n16062, n16063, n16066);
  nor g51271 (n16050, n16044, n16045, n16046, n16049);
  nor g51272 (n16032, n16026, n16027, n16028, n16031);
  nor g51273 (n16013, n16007, n16008, n16009, n16012);
  nor g51274 (n15994, n15988, n15989, n15990, n15993);
  nor g51275 (n15977, n15971, n15972, n15973, n15976);
  nor g51276 (n15959, n15953, n15954, n15955, n15958);
  nor g51277 (n15940, n15934, n15935, n15936, n15939);
  nor g51278 (n15921, n15915, n15916, n15917, n15920);
  nor g51279 (n15875, n15869, n15870, n15871, n15874);
  nor g51280 (n15899, n15893, n15894, n15895, n15898);
  nor g51281 (n16165, n16159, n16160, n16161, n16164);
  nor g51282 (n16195, n16189, n16190, n16191, n16194);
  nor g51283 (n16210, n16204, n16205, n16206, n16209);
  nor g51284 (n16225, n16219, n16220, n16221, n16224);
  nor g51285 (n16257, n16251, n16252, n16253, n16256);
  nor g51286 (n16273, n16267, n16268, n16269, n16272);
  nor g51287 (n16288, n16282, n16283, n16284, n16287);
  nor g51288 (n16301, n16295, n16296, n16297, n16300);
  nor g51289 (n16453, n16447, n16448, n16449, n16452);
  nor g51290 (n16434, n16428, n16429, n16430, n16433);
  nor g51291 (n16415, n16409, n16410, n16411, n16414);
  nor g51292 (n16395, n16389, n16390, n16391, n16394);
  nor g51293 (n16376, n16370, n16371, n16372, n16375);
  nor g51294 (n16357, n16351, n16352, n16353, n16356);
  nor g51295 (n16338, n16332, n16333, n16334, n16337);
  nor g51296 (n16847, n16841, n16842, n16843, n16846);
  nor g51297 (n16538, n16532, n16533, n16534, n16537);
  nor g51298 (n16553, n16547, n16548, n16549, n16552);
  nor g51299 (n16568, n16562, n16563, n16564, n16567);
  nor g51300 (n16585, n16579, n16580, n16581, n16584);
  nor g51301 (n16776, n16770, n16771, n16772, n16775);
  nor g51302 (n16600, n16594, n16595, n16596, n16599);
  nor g51303 (n16750, n16744, n16745, n16746, n16749);
  nor g51304 (n16731, n16725, n16726, n16727, n16730);
  nor g51305 (n16611, n16605, n16606, n16607, n16610);
  nor g51306 (n16623, n16617, n16618, n16619, n16622);
  nor g51307 (n16698, n16692, n16693, n16694, n16697);
  nor g51308 (n16679, n16673, n16674, n16675, n16678);
  nor g51309 (n16662, n16656, n16657, n16658, n16661);
  nor g51310 (n16648, n16642, n16643, n16644, n16647);
  nor g51311 (n16900, n16894, n16895, n16896, n16899);
  nor g51312 (n16917, n16911, n16912, n16913, n16916);
  nor g51313 (n16931, n16925, n16926, n16927, n16930);
  nor g51314 (n16947, n16941, n16942, n16943, n16946);
  nor g51315 (n17219, n17213, n17214, n17215, n17218);
  nor g51316 (n16962, n16956, n16957, n16958, n16961);
  nor g51317 (n16978, n16972, n16973, n16974, n16977);
  nor g51318 (n16994, n16988, n16989, n16990, n16993);
  nor g51319 (n17188, n17182, n17183, n17184, n17187);
  nor g51320 (n17171, n17165, n17166, n17167, n17170);
  nor g51321 (n17153, n17147, n17148, n17149, n17152);
  nor g51322 (n17134, n17128, n17129, n17130, n17133);
  nor g51323 (n17115, n17109, n17110, n17111, n17114);
  nor g51324 (n17013, n17007, n17008, n17009, n17012);
  nor g51325 (n17088, n17082, n17083, n17084, n17087);
  nor g51326 (n17024, n17018, n17019, n17020, n17023);
  nor g51327 (n17063, n17057, n17058, n17059, n17062);
  nor g51328 (n17037, n17031, n17032, n17033, n17036);
  nor g51329 (n17264, n17258, n17259, n17260, n17263);
  nor g51330 (n17280, n17274, n17275, n17276, n17279);
  nor g51331 (n17295, n17289, n17290, n17291, n17294);
  nor g51332 (n17310, n17304, n17305, n17306, n17309);
  nor g51333 (n17327, n17321, n17322, n17323, n17326);
  nor g51334 (n17342, n17336, n17337, n17338, n17341);
  nor g51335 (n17354, n17348, n17349, n17350, n17353);
  nor g51336 (n17367, n17361, n17362, n17363, n17366);
  nor g51337 (n17503, n17497, n17498, n17499, n17502);
  nor g51338 (n17484, n17478, n17479, n17480, n17483);
  nor g51339 (n17465, n17459, n17460, n17461, n17464);
  nor g51340 (n17446, n17440, n17441, n17442, n17445);
  nor g51341 (n17427, n17421, n17422, n17423, n17426);
  nor g51342 (n17408, n17402, n17403, n17404, n17407);
  nor g51343 (n17378, n17372, n17373, n17374, n17377);
  nor g51344 (n17655, n17649, n17650, n17651, n17654);
  nor g51345 (n17670, n17664, n17665, n17666, n17669);
  nor g51346 (n17701, n17695, n17696, n17697, n17700);
  nor g51347 (n17731, n17725, n17726, n17727, n17730);
  nor g51348 (n17901, n17895, n17896, n17897, n17900);
  nor g51349 (n17743, n17737, n17738, n17739, n17742);
  nor g51350 (n17875, n17869, n17870, n17871, n17874);
  nor g51351 (n17856, n17850, n17851, n17852, n17855);
  nor g51352 (n17755, n17749, n17750, n17751, n17754);
  nor g51353 (n17767, n17761, n17762, n17763, n17766);
  nor g51354 (n17825, n17819, n17820, n17821, n17824);
  nor g51355 (n17806, n17800, n17801, n17802, n17805);
  nor g51356 (n17791, n17785, n17786, n17787, n17790);
  nor g51357 (n17981, n17975, n17976, n17977, n17980);
  nor g51358 (n17997, n17991, n17992, n17993, n17996);
  nor g51359 (n18011, n18005, n18006, n18007, n18010);
  nor g51360 (n18027, n18021, n18022, n18023, n18026);
  nor g51361 (n18042, n18036, n18037, n18038, n18041);
  nor g51362 (n18058, n18052, n18053, n18054, n18057);
  nor g51363 (n18273, n18267, n18268, n18269, n18272);
  nor g51364 (n18255, n18249, n18250, n18251, n18254);
  nor g51365 (n18237, n18231, n18232, n18233, n18236);
  nor g51366 (n18220, n18214, n18215, n18216, n18219);
  nor g51367 (n18202, n18196, n18197, n18198, n18201);
  nor g51368 (n18183, n18177, n18178, n18179, n18182);
  nor g51369 (n18164, n18158, n18159, n18160, n18163);
  nor g51370 (n18078, n18072, n18073, n18074, n18077);
  nor g51371 (n18137, n18131, n18132, n18133, n18136);
  nor g51372 (n18118, n18112, n18113, n18114, n18117);
  nor g51373 (n18090, n18084, n18085, n18086, n18089);
  nor g51374 (n18326, n18320, n18321, n18322, n18325);
  nor g51375 (n18342, n18336, n18337, n18338, n18341);
  nor g51376 (n18358, n18352, n18353, n18354, n18357);
  nor g51377 (n18374, n18368, n18369, n18370, n18373);
  nor g51378 (n18387, n18381, n18382, n18383, n18386);
  nor g51379 (n18399, n18393, n18394, n18395, n18398);
  nor g51380 (n18412, n18406, n18407, n18408, n18411);
  nor g51381 (n18423, n18417, n18418, n18419, n18422);
  nor g51382 (n18519, n18513, n18514, n18515, n18518);
  nor g51383 (n18500, n18494, n18495, n18496, n18499);
  nor g51384 (n18481, n18475, n18476, n18477, n18480);
  nor g51385 (n18462, n18456, n18457, n18458, n18461);
  nor g51386 (n18444, n18438, n18439, n18440, n18443);
  nor g51387 (n18683, n18677, n18678, n18679, n18682);
  nor g51388 (n18698, n18692, n18693, n18694, n18697);
  nor g51389 (n18713, n18707, n18708, n18709, n18712);
  nor g51390 (n18743, n18737, n18738, n18739, n18742);
  nor g51391 (n18755, n18749, n18750, n18751, n18754);
  nor g51392 (n18904, n18898, n18899, n18900, n18903);
  nor g51393 (n18885, n18879, n18880, n18881, n18884);
  nor g51394 (n18868, n18862, n18863, n18864, n18867);
  nor g51395 (n18848, n18842, n18843, n18844, n18847);
  nor g51396 (n18769, n18763, n18764, n18765, n18768);
  nor g51397 (n18825, n18819, n18820, n18821, n18824);
  nor g51398 (n18806, n18800, n18801, n18802, n18805);
  nor g51399 (n18996, n18990, n18991, n18992, n18995);
  nor g51400 (n19011, n19005, n19006, n19007, n19010);
  nor g51401 (n19027, n19021, n19022, n19023, n19026);
  nor g51402 (n19041, n19035, n19036, n19037, n19040);
  nor g51403 (n19056, n19050, n19051, n19052, n19055);
  nor g51404 (n19273, n19267, n19268, n19269, n19272);
  nor g51405 (n19253, n19247, n19248, n19249, n19252);
  nor g51406 (n19236, n19230, n19231, n19232, n19235);
  nor g51407 (n19218, n19212, n19213, n19214, n19217);
  nor g51408 (n19201, n19195, n19196, n19197, n19200);
  nor g51409 (n19183, n19177, n19178, n19179, n19182);
  nor g51410 (n19164, n19158, n19159, n19160, n19163);
  nor g51411 (n19145, n19139, n19140, n19141, n19144);
  nor g51412 (n19126, n19120, n19121, n19122, n19125);
  nor g51413 (n19107, n19101, n19102, n19103, n19106);
  nor g51414 (n19088, n19082, n19083, n19084, n19087);
  nor g51415 (n19333, n19327, n19328, n19329, n19332);
  nor g51416 (n19364, n19358, n19359, n19360, n19363);
  nor g51417 (n19379, n19373, n19374, n19375, n19378);
  nor g51418 (n19395, n19389, n19390, n19391, n19394);
  nor g51419 (n19588, n19582, n19583, n19584, n19587);
  nor g51420 (n19410, n19404, n19405, n19406, n19409);
  nor g51421 (n19423, n19417, n19418, n19419, n19422);
  nor g51422 (n19435, n19429, n19430, n19431, n19434);
  nor g51423 (n19547, n19541, n19542, n19543, n19546);
  nor g51424 (n19448, n19442, n19443, n19444, n19447);
  nor g51425 (n19521, n19515, n19516, n19517, n19520);
  nor g51426 (n19503, n19497, n19498, n19499, n19502);
  nor g51427 (n19484, n19478, n19479, n19480, n19483);
  nor g51428 (n19649, n19643, n19644, n19645, n19648);
  nor g51429 (n19664, n19658, n19659, n19660, n19663);
  nor g51430 (n19680, n19674, n19675, n19676, n19679);
  nor g51431 (n19695, n19689, n19690, n19691, n19694);
  nor g51432 (n19711, n19705, n19706, n19707, n19710);
  nor g51433 (n19901, n19895, n19896, n19897, n19900);
  nor g51434 (n19727, n19721, n19722, n19723, n19726);
  nor g51435 (n19739, n19733, n19734, n19735, n19738);
  nor g51436 (n19872, n19866, n19867, n19868, n19871);
  nor g51437 (n19852, n19846, n19847, n19848, n19851);
  nor g51438 (n19834, n19828, n19829, n19830, n19833);
  nor g51439 (n19813, n19807, n19808, n19809, n19812);
  nor g51440 (n19752, n19746, n19747, n19748, n19751);
  nor g51441 (n19790, n19784, n19785, n19786, n19789);
  nor g51442 (n19764, n19758, n19759, n19760, n19763);
  nor g51443 (n19949, n19943, n19944, n19945, n19948);
  nor g51444 (n19964, n19958, n19959, n19960, n19963);
  nor g51445 (n20214, n20208, n20209, n20210, n20213);
  nor g51446 (n19979, n19973, n19974, n19975, n19978);
  nor g51447 (n20191, n20185, n20186, n20187, n20190);
  nor g51448 (n20172, n20166, n20167, n20168, n20171);
  nor g51449 (n20153, n20147, n20148, n20149, n20152);
  nor g51450 (n20136, n20130, n20131, n20132, n20135);
  nor g51451 (n20118, n20112, n20113, n20114, n20117);
  nor g51452 (n20101, n20095, n20096, n20097, n20100);
  nor g51453 (n20082, n20076, n20077, n20078, n20081);
  nor g51454 (n20063, n20057, n20058, n20059, n20062);
  nor g51455 (n19998, n19992, n19993, n19994, n19997);
  nor g51456 (n20038, n20032, n20033, n20034, n20037);
  nor g51457 (n20010, n20004, n20005, n20006, n20009);
  nor g51458 (n20251, n20245, n20246, n20247, n20250);
  nor g51459 (n20266, n20260, n20261, n20262, n20265);
  nor g51460 (n20281, n20275, n20276, n20277, n20280);
  nor g51461 (n20296, n20290, n20291, n20292, n20295);
  nor g51462 (n20489, n20483, n20484, n20485, n20488);
  nor g51463 (n20470, n20464, n20465, n20466, n20469);
  nor g51464 (n20311, n20305, n20306, n20307, n20310);
  nor g51465 (n20324, n20318, n20319, n20320, n20323);
  nor g51466 (n20437, n20431, n20432, n20433, n20436);
  nor g51467 (n20417, n20411, n20412, n20413, n20416);
  nor g51468 (n20336, n20330, n20331, n20332, n20335);
  nor g51469 (n20391, n20385, n20386, n20387, n20390);
  nor g51470 (n20348, n20342, n20343, n20344, n20347);
  nor g51471 (n20366, n20360, n20361, n20362, n20365);
  nor g51472 (n20560, n20554, n20555, n20556, n20559);
  nor g51473 (n20576, n20570, n20571, n20572, n20575);
  nor g51474 (n20591, n20585, n20586, n20587, n20590);
  nor g51475 (n20607, n20601, n20602, n20603, n20606);
  nor g51476 (n20794, n20788, n20789, n20790, n20793);
  nor g51477 (n20775, n20769, n20770, n20771, n20774);
  nor g51478 (n20623, n20617, n20618, n20619, n20622);
  nor g51479 (n20635, n20629, n20630, n20631, n20634);
  nor g51480 (n20647, n20641, n20642, n20643, n20646);
  nor g51481 (n20659, n20653, n20654, n20655, n20658);
  nor g51482 (n20734, n20728, n20729, n20730, n20733);
  nor g51483 (n20713, n20707, n20708, n20709, n20712);
  nor g51484 (n20672, n20666, n20667, n20668, n20671);
  nor g51485 (n20834, n20828, n20829, n20830, n20833);
  nor g51486 (n20849, n20843, n20844, n20845, n20848);
  nor g51487 (n20866, n20860, n20861, n20862, n20865);
  nor g51488 (n20880, n20874, n20875, n20876, n20879);
  nor g51489 (n21076, n21070, n21071, n21072, n21075);
  nor g51490 (n21057, n21051, n21052, n21053, n21056);
  nor g51491 (n21038, n21032, n21033, n21034, n21037);
  nor g51492 (n21019, n21013, n21014, n21015, n21018);
  nor g51493 (n21000, n20994, n20995, n20996, n20999);
  nor g51494 (n20983, n20977, n20978, n20979, n20982);
  nor g51495 (n20964, n20958, n20959, n20960, n20963);
  nor g51496 (n20945, n20939, n20940, n20941, n20944);
  nor g51497 (n20926, n20920, n20921, n20922, n20925);
  nor g51498 (n20906, n20900, n20901, n20902, n20905);
  nor g51499 (n21132, n21126, n21127, n21128, n21131);
  nor g51500 (n21163, n21157, n21158, n21159, n21162);
  nor g51501 (n21354, n21348, n21349, n21350, n21353);
  nor g51502 (n21335, n21329, n21330, n21331, n21334);
  nor g51503 (n21316, n21310, n21311, n21312, n21315);
  nor g51504 (n21177, n21171, n21172, n21173, n21176);
  nor g51505 (n21189, n21183, n21184, n21185, n21188);
  nor g51506 (n21283, n21277, n21278, n21279, n21282);
  nor g51507 (n21263, n21257, n21258, n21259, n21262);
  nor g51508 (n21244, n21238, n21239, n21240, n21243);
  nor g51509 (n21202, n21196, n21197, n21198, n21201);
  nor g51510 (n21407, n21401, n21402, n21403, n21406);
  nor g51511 (n21422, n21416, n21417, n21418, n21421);
  nor g51512 (n21439, n21433, n21434, n21435, n21438);
  nor g51513 (n21454, n21448, n21449, n21450, n21453);
  nor g51514 (n21620, n21614, n21615, n21616, n21619);
  nor g51515 (n21601, n21595, n21596, n21597, n21600);
  nor g51516 (n21467, n21461, n21462, n21463, n21466);
  nor g51517 (n21578, n21572, n21573, n21574, n21577);
  nor g51518 (n21558, n21552, n21553, n21554, n21557);
  nor g51519 (n21480, n21474, n21475, n21476, n21479);
  nor g51520 (n21535, n21529, n21530, n21531, n21534);
  nor g51521 (n21516, n21510, n21511, n21512, n21515);
  nor g51522 (n21668, n21662, n21663, n21664, n21667);
  nor g51523 (n21685, n21679, n21680, n21681, n21684);
  nor g51524 (n21699, n21693, n21694, n21695, n21698);
  nor g51525 (n21894, n21888, n21889, n21890, n21893);
  nor g51526 (n21875, n21869, n21870, n21871, n21874);
  nor g51527 (n21856, n21850, n21851, n21852, n21855);
  nor g51528 (n21839, n21833, n21834, n21835, n21838);
  nor g51529 (n21821, n21815, n21816, n21817, n21820);
  nor g51530 (n21802, n21796, n21797, n21798, n21801);
  nor g51531 (n21719, n21713, n21714, n21715, n21718);
  nor g51532 (n21776, n21770, n21771, n21772, n21775);
  nor g51533 (n21759, n21753, n21754, n21755, n21758);
  nor g51534 (n21741, n21735, n21736, n21737, n21740);
  nor g51535 (n21933, n21927, n21928, n21929, n21932);
  nor g51536 (n22142, n22136, n22137, n22138, n22141);
  nor g51537 (n22124, n22118, n22119, n22120, n22123);
  nor g51538 (n22105, n22099, n22100, n22101, n22104);
  nor g51539 (n22086, n22080, n22081, n22082, n22085);
  nor g51540 (n21964, n21958, n21959, n21960, n21963);
  nor g51541 (n21976, n21970, n21971, n21972, n21975);
  nor g51542 (n22052, n22046, n22047, n22048, n22051);
  nor g51543 (n22033, n22027, n22028, n22029, n22032);
  nor g51544 (n22014, n22008, n22009, n22010, n22013);
  nor g51545 (n22204, n22198, n22199, n22200, n22203);
  nor g51546 (n22219, n22213, n22214, n22215, n22218);
  nor g51547 (n22235, n22229, n22230, n22231, n22234);
  nor g51548 (n22247, n22241, n22242, n22243, n22246);
  nor g51549 (n22394, n22388, n22389, n22390, n22393);
  nor g51550 (n22375, n22369, n22370, n22371, n22374);
  nor g51551 (n22260, n22254, n22255, n22256, n22259);
  nor g51552 (n22352, n22346, n22347, n22348, n22351);
  nor g51553 (n22332, n22326, n22327, n22328, n22331);
  nor g51554 (n22273, n22267, n22268, n22269, n22272);
  nor g51555 (n22285, n22279, n22280, n22281, n22284);
  nor g51556 (n22441, n22435, n22436, n22437, n22440);
  nor g51557 (n22654, n22648, n22649, n22650, n22653);
  nor g51558 (n22456, n22450, n22451, n22452, n22455);
  nor g51559 (n22629, n22623, n22624, n22625, n22628);
  nor g51560 (n22610, n22604, n22605, n22606, n22609);
  nor g51561 (n22591, n22585, n22586, n22587, n22590);
  nor g51562 (n22574, n22568, n22569, n22570, n22573);
  nor g51563 (n22556, n22550, n22551, n22552, n22555);
  nor g51564 (n22537, n22531, n22532, n22533, n22536);
  nor g51565 (n22518, n22512, n22513, n22514, n22517);
  nor g51566 (n22472, n22466, n22467, n22468, n22471);
  nor g51567 (n22500, n22494, n22495, n22496, n22499);
  nor g51568 (n22696, n22690, n22691, n22692, n22695);
  nor g51569 (n22711, n22705, n22706, n22707, n22710);
  nor g51570 (n22882, n22876, n22877, n22878, n22881);
  nor g51571 (n22864, n22858, n22859, n22860, n22863);
  nor g51572 (n22845, n22839, n22840, n22841, n22844);
  nor g51573 (n22826, n22820, n22821, n22822, n22825);
  nor g51574 (n22723, n22717, n22718, n22719, n22722);
  nor g51575 (n22735, n22729, n22730, n22731, n22734);
  nor g51576 (n22792, n22786, n22787, n22788, n22791);
  nor g51577 (n22747, n22741, n22742, n22743, n22746);
  nor g51578 (n22765, n22759, n22760, n22761, n22764);
  nor g51579 (n22933, n22927, n22928, n22929, n22932);
  nor g51580 (n23125, n23119, n23120, n23121, n23124);
  nor g51581 (n22950, n22944, n22945, n22946, n22949);
  nor g51582 (n22962, n22956, n22957, n22958, n22961);
  nor g51583 (n23094, n23088, n23089, n23090, n23093);
  nor g51584 (n23075, n23069, n23070, n23071, n23074);
  nor g51585 (n22975, n22969, n22970, n22971, n22974);
  nor g51586 (n23052, n23046, n23047, n23048, n23051);
  nor g51587 (n23031, n23025, n23026, n23027, n23030);
  nor g51588 (n22988, n22982, n22983, n22984, n22987);
  nor g51589 (n23011, n23005, n23006, n23007, n23010);
  nor g51590 (n23356, n23350, n23351, n23352, n23355);
  nor g51591 (n23336, n23330, n23331, n23332, n23335);
  nor g51592 (n23156, n23150, n23151, n23152, n23155);
  nor g51593 (n23311, n23305, n23306, n23307, n23310);
  nor g51594 (n23292, n23286, n23287, n23288, n23291);
  nor g51595 (n23273, n23267, n23268, n23269, n23272);
  nor g51596 (n23256, n23250, n23251, n23252, n23255);
  nor g51597 (n23238, n23232, n23233, n23234, n23237);
  nor g51598 (n23172, n23166, n23167, n23168, n23171);
  nor g51599 (n23213, n23207, n23208, n23209, n23212);
  nor g51600 (n23199, n23193, n23194, n23195, n23198);
  nor g51601 (n23572, n23566, n23567, n23568, n23571);
  nor g51602 (n23393, n23387, n23388, n23389, n23392);
  nor g51603 (n23547, n23541, n23542, n23543, n23546);
  nor g51604 (n23529, n23523, n23524, n23525, n23528);
  nor g51605 (n23510, n23504, n23505, n23506, n23509);
  nor g51606 (n23491, n23485, n23486, n23487, n23490);
  nor g51607 (n23405, n23399, n23400, n23401, n23404);
  nor g51608 (n23417, n23411, n23412, n23413, n23416);
  nor g51609 (n23429, n23423, n23424, n23425, n23428);
  nor g51610 (n23449, n23443, n23444, n23445, n23448);
  nor g51611 (n23790, n23784, n23785, n23786, n23789);
  nor g51612 (n23771, n23765, n23766, n23767, n23770);
  nor g51613 (n23616, n23610, n23611, n23612, n23615);
  nor g51614 (n23628, n23622, n23623, n23624, n23627);
  nor g51615 (n23740, n23734, n23735, n23736, n23739);
  nor g51616 (n23721, n23715, n23716, n23717, n23720);
  nor g51617 (n23641, n23635, n23636, n23637, n23640);
  nor g51618 (n23653, n23647, n23648, n23649, n23652);
  nor g51619 (n23692, n23686, n23687, n23688, n23691);
  nor g51620 (n23677, n23671, n23672, n23673, n23676);
  nor g51621 (n24000, n23994, n23995, n23996, n23999);
  nor g51622 (n23980, n23974, n23975, n23976, n23979);
  nor g51623 (n23819, n23813, n23814, n23815, n23818);
  nor g51624 (n23955, n23949, n23950, n23951, n23954);
  nor g51625 (n23936, n23930, n23931, n23932, n23935);
  nor g51626 (n23917, n23911, n23912, n23913, n23916);
  nor g51627 (n23898, n23892, n23893, n23894, n23897);
  nor g51628 (n23832, n23826, n23827, n23828, n23831);
  nor g51629 (n23873, n23867, n23868, n23869, n23872);
  nor g51630 (n23859, n23853, n23854, n23855, n23858);
  nor g51631 (n24195, n24189, n24190, n24191, n24194);
  nor g51632 (n24037, n24031, n24032, n24033, n24036);
  nor g51633 (n24170, n24164, n24165, n24166, n24169);
  nor g51634 (n24152, n24146, n24147, n24148, n24151);
  nor g51635 (n24133, n24127, n24128, n24129, n24132);
  nor g51636 (n24114, n24108, n24109, n24110, n24113);
  nor g51637 (n24049, n24043, n24044, n24045, n24048);
  nor g51638 (n24061, n24055, n24056, n24057, n24060);
  nor g51639 (n24081, n24075, n24076, n24077, n24080);
  nor g51640 (n24395, n24389, n24390, n24391, n24394);
  nor g51641 (n24376, n24370, n24371, n24372, n24375);
  nor g51642 (n24239, n24233, n24234, n24235, n24238);
  nor g51643 (n24251, n24245, n24246, n24247, n24250);
  nor g51644 (n24345, n24339, n24340, n24341, n24344);
  nor g51645 (n24326, n24320, n24321, n24322, n24325);
  nor g51646 (n24264, n24258, n24259, n24260, n24263);
  nor g51647 (n24303, n24297, n24298, n24299, n24302);
  nor g51648 (n24288, n24282, n24283, n24284, n24287);
  nor g51649 (n24579, n24573, n24574, n24575, n24578);
  nor g51650 (n24560, n24554, n24555, n24556, n24559);
  nor g51651 (n24541, n24535, n24536, n24537, n24540);
  nor g51652 (n24421, n24415, n24416, n24417, n24420);
  nor g51653 (n24518, n24512, n24513, n24514, n24517);
  nor g51654 (n24499, n24493, n24494, n24495, n24498);
  nor g51655 (n24480, n24474, n24475, n24476, n24479);
  nor g51656 (n24459, n24453, n24454, n24455, n24458);
  nor g51657 (n24445, n24439, n24440, n24441, n24444);
  nor g51658 (n24762, n24756, n24757, n24758, n24761);
  nor g51659 (n24743, n24737, n24738, n24739, n24742);
  nor g51660 (n24724, n24718, n24719, n24720, n24723);
  nor g51661 (n24704, n24698, n24699, n24700, n24703);
  nor g51662 (n24685, n24679, n24680, n24681, n24684);
  nor g51663 (n24666, n24660, n24661, n24662, n24665);
  nor g51664 (n24647, n24641, n24642, n24643, n24646);
  nor g51665 (n24619, n24613, n24614, n24615, n24618);
  nor g51666 (n24942, n24936, n24937, n24938, n24941);
  nor g51667 (n24923, n24917, n24918, n24919, n24922);
  nor g51668 (n24804, n24798, n24799, n24800, n24803);
  nor g51669 (n24816, n24810, n24811, n24812, n24815);
  nor g51670 (n24892, n24886, n24887, n24888, n24891);
  nor g51671 (n24873, n24867, n24868, n24869, n24872);
  nor g51672 (n24855, n24849, n24850, n24851, n24854);
  nor g51673 (n24840, n24834, n24835, n24836, n24839);
  nor g51674 (n25109, n25103, n25104, n25105, n25108);
  nor g51675 (n25090, n25084, n25085, n25086, n25089);
  nor g51676 (n25071, n25065, n25066, n25067, n25070);
  nor g51677 (n24968, n24962, n24963, n24964, n24967);
  nor g51678 (n25048, n25042, n25043, n25044, n25047);
  nor g51679 (n25029, n25023, n25024, n25025, n25028);
  nor g51680 (n25008, n25002, n25003, n25004, n25007);
  nor g51681 (n24993, n24987, n24988, n24989, n24992);
  nor g51682 (n25271, n25265, n25266, n25267, n25270);
  nor g51683 (n25252, n25246, n25247, n25248, n25251);
  nor g51684 (n25233, n25227, n25228, n25229, n25232);
  nor g51685 (n25213, n25207, n25208, n25209, n25212);
  nor g51686 (n25194, n25188, n25189, n25190, n25193);
  nor g51687 (n25175, n25169, n25170, n25171, n25174);
  nor g51688 (n25433, n25427, n25428, n25429, n25432);
  nor g51689 (n25312, n25306, n25307, n25308, n25311);
  nor g51690 (n25324, n25318, n25319, n25320, n25323);
  nor g51691 (n25336, n25330, n25331, n25332, n25335);
  nor g51692 (n25392, n25386, n25387, n25388, n25391);
  nor g51693 (n25375, n25369, n25370, n25371, n25374);
  nor g51694 (n25361, n25355, n25356, n25357, n25360);
  nor g51695 (n25581, n25575, n25576, n25577, n25580);
  nor g51696 (n25458, n25452, n25453, n25454, n25457);
  nor g51697 (n25470, n25464, n25465, n25466, n25469);
  nor g51698 (n25550, n25544, n25545, n25546, n25549);
  nor g51699 (n25483, n25477, n25478, n25479, n25482);
  nor g51700 (n25522, n25516, n25517, n25518, n25521);
  nor g51701 (n25503, n25497, n25498, n25499, n25502);
  nor g51702 (n25621, n25615, n25616, n25617, n25620);
  nor g51703 (n25717, n25711, n25712, n25713, n25716);
  nor g51704 (n25699, n25693, n25694, n25695, n25698);
  nor g51705 (n25680, n25674, n25675, n25676, n25679);
  nor g51706 (n25661, n25655, n25656, n25657, n25660);
  nor g51707 (n25870, n25864, n25865, n25866, n25869);
  nor g51708 (n25765, n25759, n25760, n25761, n25764);
  nor g51709 (n25777, n25771, n25772, n25773, n25776);
  nor g51710 (n25789, n25783, n25784, n25785, n25788);
  nor g51711 (n25801, n25795, n25796, n25797, n25800);
  nor g51712 (n25895, n25889, n25890, n25891, n25894);
  nor g51713 (n25907, n25901, n25902, n25903, n25906);
  nor g51714 (n25919, n25913, n25914, n25915, n25918);
  nor g51715 (n25931, n25925, n25926, n25927, n25930);
  nor g51716 (n25973, n25967, n25968, n25969, n25972);
  nor g51717 (n25958, n25952, n25953, n25954, n25957);
  nor g51718 (n26037, n26031, n26032, n26033, n26036);
  nor g51719 (n26113, n26107, n26108, n26109, n26112);
  nor g51720 (n26050, n26044, n26045, n26046, n26049);
  nor g51721 (n26062, n26056, n26057, n26058, n26061);
  nor g51722 (n26081, n26075, n26076, n26077, n26080);
  nor g51723 (n26232, n26226, n26227, n26228, n26231);
  nor g51724 (n26147, n26141, n26142, n26143, n26146);
  nor g51725 (n26159, n26153, n26154, n26155, n26158);
  nor g51726 (n26171, n26165, n26166, n26167, n26170);
  nor g51727 (n26194, n26188, n26189, n26190, n26193);
  nor g51728 (n26270, n26264, n26265, n26266, n26269);
  nor g51729 (n26282, n26276, n26277, n26278, n26281);
  nor g51730 (n26294, n26288, n26289, n26290, n26293);
  nor g51731 (n26335, n26329, n26330, n26331, n26334);
  nor g51732 (n26307, n26301, n26302, n26303, n26306);
  nor g51733 (n26390, n26384, n26385, n26386, n26389);
  nor g51734 (n26402, n26396, n26397, n26398, n26401);
  nor g51735 (n26414, n26408, n26409, n26410, n26413);
  nor g51736 (n26548, n26542, n26543, n26544, n26547);
  nor g51737 (n26485, n26479, n26480, n26481, n26484);
  nor g51738 (n26523, n26517, n26518, n26519, n26522);
  nor g51739 (n26497, n26491, n26492, n26493, n26496);
  nor g51740 (n26653, n26647, n26648, n26649, n26652);
  nor g51741 (n26587, n26581, n26582, n26583, n26586);
  nor g51742 (n26599, n26593, n26594, n26595, n26598);
  nor g51743 (n26610, n26604, n26605, n26606, n26609);
  nor g51744 (n26690, n26684, n26685, n26686, n26689);
  nor g51745 (n26702, n26696, n26697, n26698, n26701);
  nor g51746 (n26721, n26715, n26716, n26717, n26720);
  nor g51747 (n26808, n26802, n26803, n26804, n26807);
  nor g51748 (n26791, n26785, n26786, n26787, n26790);
  nor g51749 (n26777, n26771, n26772, n26773, n26776);
  nor g51750 (n26849, n26843, n26844, n26845, n26848);
  nor g51751 (n26866, n26860, n26861, n26862, n26865);
  nor g51752 (n26886, n26880, n26881, n26882, n26885);
  nor g51753 (n26931, n26925, n26926, n26927, n26930);
  nor g51754 (n27016, n27010, n27011, n27012, n27015);
  nor g51755 (n26990, n26984, n26985, n26986, n26989);
  nor g51756 (n27085, n27079, n27080, n27081, n27084);
  nor g51757 (n27055, n27049, n27050, n27051, n27054);
  nor g51758 (n27172, n27166, n27167, n27168, n27171);
  nor g51759 (n27217, n27211, n27212, n27213, n27216);
endmodule
