VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO oaTaper STRING ;
END PROPERTYDEFINITIONS

MACRO AND2X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AND2X1 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.125 1.07 0.545 1.17 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.48 0.83 0.9 0.93 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.9 1.85 1 1.95 ;
        RECT 0.9 1.65 1 1.75 ;
        RECT 0.9 0.4 1 0.5 ;
        RECT 0.9 0.2 1 0.3 ;
      LAYER ME1 ;
        RECT 0.89 0.17 1.01 0.53 ;
        RECT 0.89 1.62 1.01 1.98 ;
      LAYER ME2 ;
        RECT 0.9 0.17 1 1.98 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.125 1.62 0.215 2.52 ;
        RECT 0.645 1.62 0.735 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.645 -0.22 0.735 0.53 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.18 0.17 0.3 0.53 ;
      RECT 0.37 1.62 0.49 1.98 ;
      RECT 0.125 1.07 0.545 1.17 ;
      RECT 0.35 1.27 0.88 1.37 ;
      RECT 0.48 0.83 0.9 0.93 ;
      RECT 0.89 1.62 1.01 1.98 ;
      RECT 0.89 0.17 1.01 0.53 ;
      RECT 0.125 1.62 0.215 2.52 ;
      RECT 0.645 1.62 0.735 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.645 -0.22 0.735 0.53 ;
    LAYER VI1 ;
      RECT 0.19 0.4 0.29 0.5 ;
      RECT 0.19 0.2 0.29 0.3 ;
      RECT 0.38 1.85 0.48 1.95 ;
      RECT 0.38 1.65 0.48 1.75 ;
      RECT 0.38 1.27 0.48 1.37 ;
      RECT 0.9 1.85 1 1.95 ;
      RECT 0.9 1.65 1 1.75 ;
      RECT 0.9 0.4 1 0.5 ;
      RECT 0.9 0.2 1 0.3 ;
    LAYER ME2 ;
      RECT 0.19 0.17 0.29 0.53 ;
      RECT 0.19 0.43 0.48 0.53 ;
      RECT 0.35 1.27 0.51 1.37 ;
      RECT 0.38 0.43 0.48 1.98 ;
      RECT 0.9 0.17 1 1.98 ;
  END
END AND2X1

MACRO AND2X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AND2X2 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.13 1.07 0.41 1.22 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.5 0.96 0.92 1.06 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.9 1.79 1 1.89 ;
        RECT 0.9 1.59 1 1.69 ;
        RECT 0.9 1.39 1 1.49 ;
        RECT 0.9 0.55 1 0.65 ;
        RECT 0.9 0.35 1 0.45 ;
      LAYER ME1 ;
        RECT 0.89 0.32 1.01 0.68 ;
        RECT 0.9 1.36 1 1.92 ;
        RECT 0.905 1.32 0.995 1.92 ;
      LAYER ME2 ;
        RECT 0.9 0.32 1 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.125 1.32 0.215 2.52 ;
        RECT 0.645 1.32 0.735 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.645 -0.22 0.735 0.68 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.18 0.32 0.3 0.68 ;
      RECT 0.13 1.07 0.41 1.22 ;
      RECT 0.385 1.32 0.475 1.92 ;
      RECT 0.38 1.36 0.48 1.92 ;
      RECT 0.35 0.77 0.88 0.87 ;
      RECT 0.5 0.96 0.92 1.06 ;
      RECT 0.905 1.32 0.995 1.92 ;
      RECT 0.9 1.36 1 1.92 ;
      RECT 0.89 0.32 1.01 0.68 ;
      RECT 0.125 1.32 0.215 2.52 ;
      RECT 0.645 1.32 0.735 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.645 -0.22 0.735 0.68 ;
    LAYER VI1 ;
      RECT 0.19 0.55 0.29 0.65 ;
      RECT 0.19 0.35 0.29 0.45 ;
      RECT 0.38 1.79 0.48 1.89 ;
      RECT 0.38 1.59 0.48 1.69 ;
      RECT 0.38 1.39 0.48 1.49 ;
      RECT 0.38 0.77 0.48 0.87 ;
      RECT 0.9 1.79 1 1.89 ;
      RECT 0.9 1.59 1 1.69 ;
      RECT 0.9 1.39 1 1.49 ;
      RECT 0.9 0.55 1 0.65 ;
      RECT 0.9 0.35 1 0.45 ;
    LAYER ME2 ;
      RECT 0.19 0.32 0.29 0.68 ;
      RECT 0.19 0.58 0.48 0.68 ;
      RECT 0.38 0.58 0.48 1.92 ;
      RECT 0.9 0.32 1 1.92 ;
  END
END AND2X2

MACRO AND2X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AND2X4 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.005 0.42 1.155 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.51 1.08 0.93 1.18 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.91 1.79 1.01 1.89 ;
        RECT 0.91 1.59 1.01 1.69 ;
        RECT 0.91 1.39 1.01 1.49 ;
        RECT 0.91 0.55 1.01 0.65 ;
        RECT 0.91 0.35 1.01 0.45 ;
      LAYER ME1 ;
        RECT 0.9 0.32 1.02 0.68 ;
        RECT 0.91 1.36 1.01 1.92 ;
        RECT 0.915 1.32 1.005 1.92 ;
      LAYER ME2 ;
        RECT 0.91 0.32 1.01 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 1.32 0.225 2.52 ;
        RECT 0.655 1.32 0.745 2.52 ;
        RECT 1.175 1.32 1.265 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.655 -0.22 0.745 0.68 ;
        RECT 1.175 -0.22 1.265 0.68 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.19 0.32 0.31 0.68 ;
      RECT 0.14 1.005 0.42 1.155 ;
      RECT 0.395 1.32 0.485 1.92 ;
      RECT 0.39 1.36 0.49 1.92 ;
      RECT 0.51 1.08 0.93 1.18 ;
      RECT 0.915 1.32 1.005 1.92 ;
      RECT 0.91 1.36 1.01 1.92 ;
      RECT 0.9 0.32 1.02 0.68 ;
      RECT 0.36 0.8 1.12 0.89 ;
      RECT 0.36 0.795 0.52 0.895 ;
      RECT 0.135 1.32 0.225 2.52 ;
      RECT 0.655 1.32 0.745 2.52 ;
      RECT 1.175 1.32 1.265 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.655 -0.22 0.745 0.68 ;
      RECT 1.175 -0.22 1.265 0.68 ;
    LAYER VI1 ;
      RECT 0.2 0.55 0.3 0.65 ;
      RECT 0.2 0.35 0.3 0.45 ;
      RECT 0.39 1.79 0.49 1.89 ;
      RECT 0.39 1.59 0.49 1.69 ;
      RECT 0.39 1.39 0.49 1.49 ;
      RECT 0.39 0.795 0.49 0.895 ;
      RECT 0.91 1.79 1.01 1.89 ;
      RECT 0.91 1.59 1.01 1.69 ;
      RECT 0.91 1.39 1.01 1.49 ;
      RECT 0.91 0.55 1.01 0.65 ;
      RECT 0.91 0.35 1.01 0.45 ;
    LAYER ME2 ;
      RECT 0.2 0.32 0.3 0.68 ;
      RECT 0.2 0.58 0.49 0.68 ;
      RECT 0.39 0.58 0.49 1.92 ;
      RECT 0.91 0.32 1.01 1.92 ;
  END
END AND2X4

MACRO AOI211X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI211X1 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.3 1.165 0.72 1.265 ;
    END
  END A2
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.43 1.62 0.52 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.17 -0.22 0.26 0.53 ;
        RECT 0.88 -0.22 0.97 0.53 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.17 0.865 0.59 0.965 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.815 1.145 1.235 1.245 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.135 1.85 1.235 1.95 ;
        RECT 1.135 1.65 1.235 1.75 ;
        RECT 1.135 0.61 1.235 0.71 ;
        RECT 1.135 0.41 1.235 0.51 ;
      LAYER ME1 ;
        RECT 0.62 0.65 1.245 0.74 ;
        RECT 1.125 0.38 1.245 0.74 ;
        RECT 0.62 0.38 0.71 0.74 ;
        RECT 1.125 1.62 1.245 1.98 ;
      LAYER ME2 ;
        RECT 1.135 0.38 1.235 1.98 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.685 0.885 1.105 0.985 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.17 0.865 0.59 0.965 ;
      RECT 0.3 1.165 0.72 1.265 ;
      RECT 0.17 1.44 0.78 1.53 ;
      RECT 0.17 1.44 0.26 1.92 ;
      RECT 0.69 1.44 0.78 1.92 ;
      RECT 0.685 0.885 1.105 0.985 ;
      RECT 0.815 1.145 1.235 1.245 ;
      RECT 1.125 1.62 1.245 1.98 ;
      RECT 0.62 0.38 0.71 0.74 ;
      RECT 1.125 0.38 1.245 0.74 ;
      RECT 0.62 0.65 1.245 0.74 ;
      RECT 0.43 1.62 0.52 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.17 -0.22 0.26 0.53 ;
      RECT 0.88 -0.22 0.97 0.53 ;
    LAYER VI1 ;
      RECT 1.135 1.85 1.235 1.95 ;
      RECT 1.135 1.65 1.235 1.75 ;
      RECT 1.135 0.61 1.235 0.71 ;
      RECT 1.135 0.41 1.235 0.51 ;
    LAYER ME2 ;
      RECT 1.135 0.38 1.235 1.98 ;
  END
END AOI211X1

MACRO AOI211X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI211X2 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.31 1.105 0.73 1.205 ;
    END
  END A2
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.43 1.32 0.52 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.17 -0.22 0.26 0.68 ;
        RECT 0.88 -0.22 0.97 0.68 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.17 0.835 0.59 0.935 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.845 1.075 1.265 1.175 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.61 0.21 0.71 0.31 ;
        RECT 1.135 1.79 1.235 1.89 ;
        RECT 1.135 1.59 1.235 1.69 ;
        RECT 1.135 1.39 1.235 1.49 ;
        RECT 1.135 0.55 1.235 0.65 ;
        RECT 1.135 0.35 1.235 0.45 ;
      LAYER ME1 ;
        RECT 1.125 0.32 1.245 0.68 ;
        RECT 1.135 1.36 1.235 1.92 ;
        RECT 1.14 1.32 1.23 1.92 ;
        RECT 0.58 0.21 0.74 0.31 ;
        RECT 0.62 0.21 0.71 0.68 ;
      LAYER ME2 ;
        RECT 1.135 0.21 1.235 1.92 ;
        RECT 0.58 0.21 1.235 0.31 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.715 0.835 1.135 0.935 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.17 1.32 0.26 2.11 ;
      RECT 0.17 2.01 0.33 2.11 ;
      RECT 0.17 0.835 0.59 0.935 ;
      RECT 0.31 1.105 0.73 1.205 ;
      RECT 0.58 0.21 0.74 0.31 ;
      RECT 0.62 0.21 0.71 0.68 ;
      RECT 0.69 1.32 0.78 2.11 ;
      RECT 0.66 2.01 0.82 2.11 ;
      RECT 0.715 0.835 1.135 0.935 ;
      RECT 1.14 1.32 1.23 1.92 ;
      RECT 1.135 1.36 1.235 1.92 ;
      RECT 1.125 0.32 1.245 0.68 ;
      RECT 0.845 1.075 1.265 1.175 ;
      RECT 0.43 1.32 0.52 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.17 -0.22 0.26 0.68 ;
      RECT 0.88 -0.22 0.97 0.68 ;
    LAYER VI1 ;
      RECT 0.2 2.01 0.3 2.11 ;
      RECT 0.61 0.21 0.71 0.31 ;
      RECT 0.69 2.01 0.79 2.11 ;
      RECT 1.135 1.79 1.235 1.89 ;
      RECT 1.135 1.59 1.235 1.69 ;
      RECT 1.135 1.39 1.235 1.49 ;
      RECT 1.135 0.55 1.235 0.65 ;
      RECT 1.135 0.35 1.235 0.45 ;
    LAYER ME2 ;
      RECT 0.17 2.01 0.82 2.11 ;
      RECT 0.58 0.21 1.235 0.31 ;
      RECT 1.135 0.21 1.235 1.92 ;
  END
END AOI211X2

MACRO AOI211X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI211X4 0 -0.11 ;
  SIZE 2.24 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.105 1.105 0.525 1.205 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.55 0.55 0.65 0.65 ;
        RECT 0.55 0.35 0.65 0.45 ;
        RECT 1.26 0.55 1.36 0.65 ;
        RECT 1.26 0.35 1.36 0.45 ;
        RECT 1.33 1.79 1.43 1.89 ;
        RECT 1.33 1.59 1.43 1.69 ;
        RECT 1.33 1.39 1.43 1.49 ;
        RECT 1.78 0.55 1.88 0.65 ;
        RECT 1.78 0.35 1.88 0.45 ;
      LAYER ME1 ;
        RECT 1.77 0.32 1.89 0.68 ;
        RECT 1.33 1.36 1.43 1.92 ;
        RECT 1.335 1.32 1.425 1.92 ;
        RECT 1.25 0.32 1.37 0.68 ;
        RECT 0.54 0.32 0.66 0.68 ;
      LAYER ME2 ;
        RECT 1.78 0.32 1.88 0.68 ;
        RECT 0.55 0.55 1.88 0.65 ;
        RECT 1.33 1.36 1.445 1.92 ;
        RECT 1.345 0.38 1.445 1.92 ;
        RECT 1.26 0.32 1.36 0.68 ;
        RECT 0.55 0.32 0.65 0.68 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 1.32 0.195 2.52 ;
        RECT 0.625 1.32 0.715 2.52 ;
        RECT 2.045 1.32 2.135 2.52 ;
        RECT 0 2.3 2.24 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 -0.22 0.195 0.68 ;
        RECT 1.005 -0.22 1.095 0.68 ;
        RECT 1.525 -0.22 1.615 0.68 ;
        RECT 2.045 -0.22 2.135 0.68 ;
        RECT 0 -0.22 2.24 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.7 1.105 2.05 1.205 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.89 0.8 1.31 0.9 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.59 0.775 2.01 0.875 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.365 1.32 0.455 1.92 ;
      RECT 0.36 1.36 0.46 1.92 ;
      RECT 0.105 1.105 0.525 1.205 ;
      RECT 0.54 0.32 0.66 0.68 ;
      RECT 0.89 0.8 1.31 0.9 ;
      RECT 1.25 0.32 1.37 0.68 ;
      RECT 1.335 1.32 1.425 1.92 ;
      RECT 1.33 1.36 1.43 1.92 ;
      RECT 0.88 1.36 0.98 1.92 ;
      RECT 0.885 1.32 0.975 2.12 ;
      RECT 1.785 1.32 1.875 2.12 ;
      RECT 0.885 2.03 1.875 2.12 ;
      RECT 1.77 0.32 1.89 0.68 ;
      RECT 1.59 0.775 2.01 0.875 ;
      RECT 0.7 1.105 2.05 1.205 ;
      RECT 0.105 1.32 0.195 2.52 ;
      RECT 0.625 1.32 0.715 2.52 ;
      RECT 2.045 1.32 2.135 2.52 ;
      RECT 0 2.3 2.24 2.52 ;
      RECT 0 -0.22 2.24 0 ;
      RECT 0.105 -0.22 0.195 0.68 ;
      RECT 1.005 -0.22 1.095 0.68 ;
      RECT 1.525 -0.22 1.615 0.68 ;
      RECT 2.045 -0.22 2.135 0.68 ;
    LAYER VI1 ;
      RECT 0.36 1.79 0.46 1.89 ;
      RECT 0.36 1.59 0.46 1.69 ;
      RECT 0.36 1.39 0.46 1.49 ;
      RECT 0.55 0.55 0.65 0.65 ;
      RECT 0.55 0.35 0.65 0.45 ;
      RECT 0.88 1.79 0.98 1.89 ;
      RECT 0.88 1.59 0.98 1.69 ;
      RECT 0.88 1.39 0.98 1.49 ;
      RECT 1.26 0.55 1.36 0.65 ;
      RECT 1.26 0.35 1.36 0.45 ;
      RECT 1.33 1.79 1.43 1.89 ;
      RECT 1.33 1.59 1.43 1.69 ;
      RECT 1.33 1.39 1.43 1.49 ;
      RECT 1.78 0.55 1.88 0.65 ;
      RECT 1.78 0.35 1.88 0.45 ;
    LAYER ME2 ;
      RECT 0.36 1.59 0.98 1.69 ;
      RECT 0.36 1.36 0.46 1.92 ;
      RECT 0.88 1.36 0.98 1.92 ;
      RECT 0.55 0.55 1.88 0.65 ;
      RECT 0.55 0.32 0.65 0.68 ;
      RECT 1.26 0.32 1.36 0.68 ;
      RECT 1.78 0.32 1.88 0.68 ;
      RECT 1.345 0.38 1.445 1.92 ;
      RECT 1.33 1.36 1.445 1.92 ;
  END
END AOI211X4

MACRO AOI21X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI21X1 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.355 1.24 0.775 1.34 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.83 0.58 0.93 0.68 ;
        RECT 0.83 0.38 0.93 0.48 ;
        RECT 0.9 1.85 1 1.95 ;
        RECT 0.9 1.65 1 1.75 ;
      LAYER ME1 ;
        RECT 0.89 1.62 1.01 1.98 ;
        RECT 0.125 0.62 0.93 0.71 ;
        RECT 0.83 0.35 0.93 0.71 ;
        RECT 0.125 0.38 0.215 0.71 ;
      LAYER ME2 ;
        RECT 0.83 1.62 1 1.98 ;
        RECT 0.83 0.35 0.93 1.98 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.385 1.62 0.475 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.575 -0.22 0.665 0.53 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.125 0.82 0.545 0.92 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.51 1.025 0.93 1.125 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.125 0.82 0.545 0.92 ;
      RECT 0.125 1.44 0.735 1.53 ;
      RECT 0.125 1.44 0.215 1.92 ;
      RECT 0.645 1.44 0.735 1.92 ;
      RECT 0.355 1.24 0.775 1.34 ;
      RECT 0.51 1.025 0.93 1.125 ;
      RECT 0.125 0.38 0.215 0.71 ;
      RECT 0.83 0.35 0.93 0.71 ;
      RECT 0.125 0.62 0.93 0.71 ;
      RECT 0.89 1.62 1.01 1.98 ;
      RECT 0.385 1.62 0.475 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.575 -0.22 0.665 0.53 ;
    LAYER VI1 ;
      RECT 0.83 0.58 0.93 0.68 ;
      RECT 0.83 0.38 0.93 0.48 ;
      RECT 0.9 1.85 1 1.95 ;
      RECT 0.9 1.65 1 1.75 ;
    LAYER ME2 ;
      RECT 0.83 0.35 0.93 1.98 ;
      RECT 0.83 1.62 1 1.98 ;
  END
END AOI21X1

MACRO AOI21X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI21X2 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.305 1.095 0.725 1.195 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.12 0.55 0.22 0.65 ;
        RECT 0.12 0.35 0.22 0.45 ;
        RECT 0.83 0.55 0.93 0.65 ;
        RECT 0.83 0.35 0.93 0.45 ;
        RECT 0.9 1.79 1 1.89 ;
        RECT 0.9 1.59 1 1.69 ;
        RECT 0.9 1.39 1 1.49 ;
      LAYER ME1 ;
        RECT 0.9 1.36 1 1.92 ;
        RECT 0.905 1.32 0.995 1.92 ;
        RECT 0.82 0.32 0.94 0.68 ;
        RECT 0.11 0.32 0.23 0.68 ;
      LAYER ME2 ;
        RECT 0.9 0.32 1 1.92 ;
        RECT 0.83 0.32 1 0.68 ;
        RECT 0.12 0.45 1 0.55 ;
        RECT 0.12 0.32 0.22 0.68 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.385 1.32 0.475 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.575 -0.22 0.665 0.68 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.09 0.87 0.51 0.97 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.6 0.87 1.02 0.97 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.125 1.32 0.215 1.92 ;
      RECT 0.12 1.36 0.22 1.92 ;
      RECT 0.11 0.32 0.23 0.68 ;
      RECT 0.09 0.87 0.51 0.97 ;
      RECT 0.305 1.095 0.725 1.195 ;
      RECT 0.645 1.32 0.735 1.92 ;
      RECT 0.64 1.36 0.74 1.92 ;
      RECT 0.82 0.32 0.94 0.68 ;
      RECT 0.905 1.32 0.995 1.92 ;
      RECT 0.9 1.36 1 1.92 ;
      RECT 0.6 0.87 1.02 0.97 ;
      RECT 0.385 1.32 0.475 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.575 -0.22 0.665 0.68 ;
    LAYER VI1 ;
      RECT 0.12 1.79 0.22 1.89 ;
      RECT 0.12 1.59 0.22 1.69 ;
      RECT 0.12 1.39 0.22 1.49 ;
      RECT 0.12 0.55 0.22 0.65 ;
      RECT 0.12 0.35 0.22 0.45 ;
      RECT 0.64 1.79 0.74 1.89 ;
      RECT 0.64 1.59 0.74 1.69 ;
      RECT 0.64 1.39 0.74 1.49 ;
      RECT 0.83 0.55 0.93 0.65 ;
      RECT 0.83 0.35 0.93 0.45 ;
      RECT 0.9 1.79 1 1.89 ;
      RECT 0.9 1.59 1 1.69 ;
      RECT 0.9 1.39 1 1.49 ;
    LAYER ME2 ;
      RECT 0.12 1.59 0.74 1.69 ;
      RECT 0.12 1.36 0.22 1.92 ;
      RECT 0.64 1.36 0.74 1.92 ;
      RECT 0.12 0.45 1 0.55 ;
      RECT 0.12 0.32 0.22 0.68 ;
      RECT 0.83 0.32 1 0.68 ;
      RECT 0.9 0.32 1 1.92 ;
  END
END AOI21X2

MACRO AOI21X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI21X4 0 -0.11 ;
  SIZE 1.96 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.22 0.865 0.64 0.965 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.665 0.55 0.765 0.65 ;
        RECT 0.665 0.35 0.765 0.45 ;
        RECT 1.185 1.79 1.285 1.89 ;
        RECT 1.185 1.59 1.285 1.69 ;
        RECT 1.185 1.39 1.285 1.49 ;
        RECT 1.375 0.55 1.475 0.65 ;
        RECT 1.375 0.35 1.475 0.45 ;
      LAYER ME1 ;
        RECT 1.365 0.32 1.485 0.68 ;
        RECT 1.185 1.36 1.285 1.92 ;
        RECT 1.19 1.32 1.28 1.92 ;
        RECT 0.655 0.32 0.775 0.68 ;
      LAYER ME2 ;
        RECT 1.185 1.26 1.475 1.36 ;
        RECT 1.375 0.32 1.475 1.36 ;
        RECT 0.665 0.45 1.475 0.55 ;
        RECT 1.185 1.26 1.285 1.92 ;
        RECT 0.665 0.32 0.765 0.68 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.15 1.32 0.24 2.52 ;
        RECT 0.67 1.32 0.76 2.52 ;
        RECT 1.725 1.32 1.815 2.52 ;
        RECT 0 2.3 1.96 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.22 -0.22 0.31 0.68 ;
        RECT 1.12 -0.22 1.21 0.68 ;
        RECT 1.64 -0.22 1.73 0.68 ;
        RECT 0 -0.22 1.96 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.67 1.095 1.09 1.195 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.32 0.865 1.74 0.965 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.41 1.32 0.5 1.92 ;
      RECT 0.405 1.36 0.505 1.92 ;
      RECT 0.22 0.865 0.64 0.965 ;
      RECT 0.655 0.32 0.775 0.68 ;
      RECT 0.67 1.095 1.09 1.195 ;
      RECT 1.19 1.32 1.28 1.92 ;
      RECT 1.185 1.36 1.285 1.92 ;
      RECT 1.365 0.32 1.485 0.68 ;
      RECT 0.925 1.36 1.025 1.92 ;
      RECT 0.93 1.32 1.02 2.12 ;
      RECT 1.465 1.32 1.555 2.12 ;
      RECT 0.93 2.03 1.555 2.12 ;
      RECT 1.32 0.865 1.74 0.965 ;
      RECT 0.15 1.32 0.24 2.52 ;
      RECT 0.67 1.32 0.76 2.52 ;
      RECT 1.725 1.32 1.815 2.52 ;
      RECT 0 2.3 1.96 2.52 ;
      RECT 0 -0.22 1.96 0 ;
      RECT 0.22 -0.22 0.31 0.68 ;
      RECT 1.12 -0.22 1.21 0.68 ;
      RECT 1.64 -0.22 1.73 0.68 ;
    LAYER VI1 ;
      RECT 0.405 1.79 0.505 1.89 ;
      RECT 0.405 1.59 0.505 1.69 ;
      RECT 0.405 1.39 0.505 1.49 ;
      RECT 0.665 0.55 0.765 0.65 ;
      RECT 0.665 0.35 0.765 0.45 ;
      RECT 0.925 1.79 1.025 1.89 ;
      RECT 0.925 1.59 1.025 1.69 ;
      RECT 0.925 1.39 1.025 1.49 ;
      RECT 1.185 1.79 1.285 1.89 ;
      RECT 1.185 1.59 1.285 1.69 ;
      RECT 1.185 1.39 1.285 1.49 ;
      RECT 1.375 0.55 1.475 0.65 ;
      RECT 1.375 0.35 1.475 0.45 ;
    LAYER ME2 ;
      RECT 0.405 1.59 1.025 1.69 ;
      RECT 0.405 1.36 0.505 1.92 ;
      RECT 0.925 1.36 1.025 1.92 ;
      RECT 0.665 0.45 1.475 0.55 ;
      RECT 0.665 0.32 0.765 0.68 ;
      RECT 1.375 0.32 1.475 1.36 ;
      RECT 1.185 1.26 1.475 1.36 ;
      RECT 1.185 1.26 1.285 1.92 ;
  END
END AOI21X4

MACRO AOI22X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI22X1 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.26 1.165 0.68 1.265 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.8 1.145 1.22 1.245 ;
    END
  END B2
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.395 1.62 0.485 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 -0.22 0.225 0.53 ;
        RECT 1.035 -0.22 1.125 0.53 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.135 0.865 0.555 0.965 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.67 0.885 1.09 0.985 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.58 0.4 0.68 0.5 ;
        RECT 0.58 0.2 0.68 0.3 ;
        RECT 0.91 1.855 1.01 1.955 ;
        RECT 0.91 1.655 1.01 1.755 ;
      LAYER ME1 ;
        RECT 0.9 1.62 1.02 1.98 ;
        RECT 0.91 1.62 1.01 1.985 ;
        RECT 0.57 0.17 0.69 0.53 ;
      LAYER ME2 ;
        RECT 0.91 1.625 1.01 1.985 ;
        RECT 0.58 1.625 1.01 1.725 ;
        RECT 0.58 0.17 0.68 1.725 ;
    END
  END Y
  OBS
    LAYER ME1 ;
      RECT 0.135 0.865 0.555 0.965 ;
      RECT 0.26 1.165 0.68 1.265 ;
      RECT 0.57 0.17 0.69 0.53 ;
      RECT 0.9 1.62 1.02 1.98 ;
      RECT 0.91 1.62 1.01 1.985 ;
      RECT 0.67 0.885 1.09 0.985 ;
      RECT 0.8 1.145 1.22 1.245 ;
      RECT 0.135 1.44 0.745 1.53 ;
      RECT 0.135 1.44 0.225 1.92 ;
      RECT 0.655 1.44 0.745 2.165 ;
      RECT 1.175 1.62 1.265 2.165 ;
      RECT 0.655 2.075 1.265 2.165 ;
      RECT 0.395 1.62 0.485 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.135 -0.22 0.225 0.53 ;
      RECT 1.035 -0.22 1.125 0.53 ;
    LAYER VI1 ;
      RECT 0.58 0.4 0.68 0.5 ;
      RECT 0.58 0.2 0.68 0.3 ;
      RECT 0.91 1.855 1.01 1.955 ;
      RECT 0.91 1.655 1.01 1.755 ;
    LAYER ME2 ;
      RECT 0.58 0.17 0.68 1.725 ;
      RECT 0.58 1.625 1.01 1.725 ;
      RECT 0.91 1.625 1.01 1.985 ;
  END
END AOI22X1

MACRO AOI22X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI22X2 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.21 1.115 0.63 1.215 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.845 0.835 1.265 0.935 ;
    END
  END B2
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.395 1.32 0.485 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 -0.22 0.225 0.68 ;
        RECT 1.035 -0.22 1.125 0.68 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.135 0.835 0.555 0.935 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.77 1.095 1.19 1.195 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.58 0.55 0.68 0.65 ;
        RECT 0.58 0.35 0.68 0.45 ;
        RECT 0.91 1.79 1.01 1.89 ;
        RECT 0.91 1.59 1.01 1.69 ;
        RECT 0.91 1.39 1.01 1.49 ;
      LAYER ME1 ;
        RECT 0.91 1.36 1.01 1.92 ;
        RECT 0.915 1.32 1.005 1.92 ;
        RECT 0.57 0.32 0.69 0.68 ;
      LAYER ME2 ;
        RECT 0.91 1.36 1.01 1.92 ;
        RECT 0.58 1.36 1.01 1.46 ;
        RECT 0.58 0.32 0.68 1.46 ;
    END
  END Y
  OBS
    LAYER ME1 ;
      RECT 0.135 1.32 0.225 2.11 ;
      RECT 0.135 2.01 0.295 2.11 ;
      RECT 0.135 0.835 0.555 0.935 ;
      RECT 0.21 1.115 0.63 1.215 ;
      RECT 0.57 0.32 0.69 0.68 ;
      RECT 0.915 1.32 1.005 1.92 ;
      RECT 0.91 1.36 1.01 1.92 ;
      RECT 0.77 1.095 1.19 1.195 ;
      RECT 0.655 1.32 0.745 2.11 ;
      RECT 1.175 1.32 1.265 2.11 ;
      RECT 0.625 2.01 1.265 2.11 ;
      RECT 0.845 0.835 1.265 0.935 ;
      RECT 0.395 1.32 0.485 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.135 -0.22 0.225 0.68 ;
      RECT 1.035 -0.22 1.125 0.68 ;
    LAYER VI1 ;
      RECT 0.165 2.01 0.265 2.11 ;
      RECT 0.58 0.55 0.68 0.65 ;
      RECT 0.58 0.35 0.68 0.45 ;
      RECT 0.655 2.01 0.755 2.11 ;
      RECT 0.91 1.79 1.01 1.89 ;
      RECT 0.91 1.59 1.01 1.69 ;
      RECT 0.91 1.39 1.01 1.49 ;
    LAYER ME2 ;
      RECT 0.135 2.01 0.785 2.11 ;
      RECT 0.58 0.32 0.68 1.46 ;
      RECT 0.58 1.36 1.01 1.46 ;
      RECT 0.91 1.36 1.01 1.92 ;
  END
END AOI22X2

MACRO AOI22X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN AOI22X4 0 -0.11 ;
  SIZE 2.52 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.62 0.55 0.72 0.65 ;
        RECT 0.62 0.35 0.72 0.45 ;
        RECT 1.47 1.22 1.57 1.32 ;
        RECT 1.52 0.55 1.62 0.65 ;
        RECT 1.52 0.35 1.62 0.45 ;
      LAYER ME2 ;
        RECT 1.52 0.32 1.62 0.68 ;
        RECT 1.47 0.38 1.57 1.35 ;
        RECT 0.62 0.445 1.62 0.555 ;
        RECT 0.62 0.32 0.72 0.68 ;
      LAYER ME1 ;
        RECT 1.475 2.01 2.085 2.1 ;
        RECT 1.995 1.32 2.085 2.1 ;
        RECT 1.47 1.19 1.57 1.35 ;
        RECT 1.475 1.19 1.565 2.1 ;
        RECT 1.51 0.32 1.63 0.68 ;
        RECT 0.61 0.32 0.73 0.68 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.61 0.855 2.03 0.955 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.545 1.065 0.965 1.165 ;
    END
  END A1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.435 1.32 0.525 2.52 ;
        RECT 0.955 1.32 1.045 2.52 ;
        RECT 0 2.3 2.52 2.52 ;
    END
  END vdd!
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.07 0.945 1.49 1.045 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.175 0.845 0.595 0.945 ;
    END
  END A2
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.175 -0.22 0.265 0.68 ;
        RECT 1.075 -0.22 1.165 0.68 ;
        RECT 1.975 -0.22 2.065 0.68 ;
        RECT 0 -0.22 2.52 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.175 1.32 0.265 1.92 ;
      RECT 0.17 1.36 0.27 1.92 ;
      RECT 0.175 0.845 0.595 0.945 ;
      RECT 0.61 0.32 0.73 0.68 ;
      RECT 0.695 1.32 0.785 1.92 ;
      RECT 0.69 1.36 0.79 1.92 ;
      RECT 0.545 1.065 0.965 1.165 ;
      RECT 1.215 1.32 1.305 1.92 ;
      RECT 1.21 1.36 1.31 1.92 ;
      RECT 1.07 0.945 1.49 1.045 ;
      RECT 1.51 0.32 1.63 0.68 ;
      RECT 1.735 1.32 1.825 1.92 ;
      RECT 1.73 1.36 1.83 1.92 ;
      RECT 1.61 0.855 2.03 0.955 ;
      RECT 1.47 1.19 1.57 1.35 ;
      RECT 1.475 1.19 1.565 2.1 ;
      RECT 1.995 1.32 2.085 2.1 ;
      RECT 1.475 2.01 2.085 2.1 ;
      RECT 2.255 1.32 2.345 1.92 ;
      RECT 2.25 1.36 2.35 1.92 ;
      RECT 0.435 1.32 0.525 2.52 ;
      RECT 0.955 1.32 1.045 2.52 ;
      RECT 0 2.3 2.52 2.52 ;
      RECT 0 -0.22 2.52 0 ;
      RECT 0.175 -0.22 0.265 0.68 ;
      RECT 1.075 -0.22 1.165 0.68 ;
      RECT 1.975 -0.22 2.065 0.68 ;
    LAYER VI1 ;
      RECT 0.17 1.79 0.27 1.89 ;
      RECT 0.17 1.59 0.27 1.69 ;
      RECT 0.17 1.39 0.27 1.49 ;
      RECT 0.62 0.55 0.72 0.65 ;
      RECT 0.62 0.35 0.72 0.45 ;
      RECT 0.69 1.79 0.79 1.89 ;
      RECT 0.69 1.59 0.79 1.69 ;
      RECT 0.69 1.39 0.79 1.49 ;
      RECT 1.21 1.79 1.31 1.89 ;
      RECT 1.21 1.59 1.31 1.69 ;
      RECT 1.21 1.39 1.31 1.49 ;
      RECT 1.47 1.22 1.57 1.32 ;
      RECT 1.52 0.55 1.62 0.65 ;
      RECT 1.52 0.35 1.62 0.45 ;
      RECT 1.73 1.79 1.83 1.89 ;
      RECT 1.73 1.59 1.83 1.69 ;
      RECT 1.73 1.39 1.83 1.49 ;
      RECT 2.25 1.79 2.35 1.89 ;
      RECT 2.25 1.59 2.35 1.69 ;
      RECT 2.25 1.39 2.35 1.49 ;
    LAYER ME2 ;
      RECT 0.62 0.445 1.62 0.555 ;
      RECT 0.62 0.32 0.72 0.68 ;
      RECT 1.52 0.32 1.62 0.68 ;
      RECT 1.47 0.38 1.57 1.35 ;
      RECT 0.17 1.585 2.35 1.695 ;
      RECT 0.17 1.36 0.27 1.92 ;
      RECT 0.69 1.36 0.79 1.92 ;
      RECT 1.21 1.36 1.31 1.92 ;
      RECT 1.73 1.36 1.83 1.92 ;
      RECT 2.25 1.36 2.35 1.92 ;
  END
END AOI22X4

MACRO BUFENX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN BUFENX1 0 -0.11 ;
  SIZE 1.68 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.175 0.845 0.595 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.41 1.85 1.51 1.95 ;
        RECT 1.41 1.65 1.51 1.75 ;
        RECT 1.41 0.4 1.51 0.5 ;
        RECT 1.41 0.2 1.51 0.3 ;
      LAYER ME1 ;
        RECT 1.4 0.17 1.52 0.53 ;
        RECT 1.4 1.62 1.52 1.98 ;
      LAYER ME2 ;
        RECT 1.41 0.17 1.51 1.98 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.175 1.62 0.265 2.52 ;
        RECT 0.965 1.62 1.055 2.52 ;
        RECT 0 2.3 1.68 2.52 ;
    END
  END vdd!
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.76 0.845 1.18 0.945 ;
    END
  END EN
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.175 -0.22 0.265 0.53 ;
        RECT 0.965 -0.22 1.055 0.53 ;
        RECT 0 -0.22 1.68 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.42 1.62 0.54 1.98 ;
      RECT 0.42 0.17 0.54 0.53 ;
      RECT 0.175 0.845 0.595 0.945 ;
      RECT 0.69 1.62 0.81 1.98 ;
      RECT 0.69 0.17 0.81 0.53 ;
      RECT 0.76 0.845 1.18 0.945 ;
      RECT 0.4 1.06 1.23 1.16 ;
      RECT 0.67 1.365 1.46 1.465 ;
      RECT 1.4 1.62 1.52 1.98 ;
      RECT 1.4 0.17 1.52 0.53 ;
      RECT 0.175 1.62 0.265 2.52 ;
      RECT 0.965 1.62 1.055 2.52 ;
      RECT 0 2.3 1.68 2.52 ;
      RECT 0 -0.22 1.68 0 ;
      RECT 0.175 -0.22 0.265 0.53 ;
      RECT 0.965 -0.22 1.055 0.53 ;
    LAYER VI1 ;
      RECT 0.43 1.85 0.53 1.95 ;
      RECT 0.43 1.65 0.53 1.75 ;
      RECT 0.43 1.06 0.53 1.16 ;
      RECT 0.43 0.4 0.53 0.5 ;
      RECT 0.43 0.2 0.53 0.3 ;
      RECT 0.7 1.85 0.8 1.95 ;
      RECT 0.7 1.65 0.8 1.75 ;
      RECT 0.7 1.365 0.8 1.465 ;
      RECT 0.7 0.4 0.8 0.5 ;
      RECT 0.7 0.2 0.8 0.3 ;
      RECT 1.41 1.85 1.51 1.95 ;
      RECT 1.41 1.65 1.51 1.75 ;
      RECT 1.41 0.4 1.51 0.5 ;
      RECT 1.41 0.2 1.51 0.3 ;
    LAYER ME2 ;
      RECT 0.43 0.17 0.53 1.98 ;
      RECT 0.7 0.17 0.8 1.98 ;
      RECT 1.41 0.17 1.51 1.98 ;
  END
END BUFENX1

MACRO BUFENX2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN BUFENX2 0 -0.11 ;
  SIZE 1.68 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.175 1.245 0.595 1.345 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.41 1.79 1.51 1.89 ;
        RECT 1.41 1.59 1.51 1.69 ;
        RECT 1.41 1.39 1.51 1.49 ;
        RECT 1.41 0.55 1.51 0.65 ;
        RECT 1.41 0.35 1.51 0.45 ;
      LAYER ME1 ;
        RECT 1.4 0.32 1.52 0.68 ;
        RECT 1.41 1.36 1.51 1.92 ;
        RECT 1.415 1.32 1.505 1.92 ;
      LAYER ME2 ;
        RECT 1.41 0.32 1.51 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.175 1.62 0.265 2.52 ;
        RECT 0.965 1.32 1.055 2.52 ;
        RECT 0 2.3 1.68 2.52 ;
    END
  END vdd!
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.52 0.99 0.94 1.09 ;
    END
  END EN
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.175 -0.22 0.265 0.53 ;
        RECT 0.965 -0.22 1.055 0.68 ;
        RECT 0 -0.22 1.68 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.42 1.56 0.54 1.92 ;
      RECT 0.42 0.32 0.54 0.68 ;
      RECT 0.175 1.245 0.595 1.345 ;
      RECT 0.705 1.32 0.795 1.92 ;
      RECT 0.7 1.36 0.8 1.92 ;
      RECT 0.69 0.32 0.81 0.68 ;
      RECT 0.52 0.99 0.94 1.09 ;
      RECT 0.4 0.78 1.2 0.88 ;
      RECT 1.03 1.04 1.45 1.14 ;
      RECT 1.415 1.32 1.505 1.92 ;
      RECT 1.41 1.36 1.51 1.92 ;
      RECT 1.4 0.32 1.52 0.68 ;
      RECT 0.175 1.62 0.265 2.52 ;
      RECT 0.965 1.32 1.055 2.52 ;
      RECT 0 2.3 1.68 2.52 ;
      RECT 0 -0.22 1.68 0 ;
      RECT 0.175 -0.22 0.265 0.53 ;
      RECT 0.965 -0.22 1.055 0.68 ;
    LAYER VI1 ;
      RECT 0.43 1.79 0.53 1.89 ;
      RECT 0.43 1.59 0.53 1.69 ;
      RECT 0.43 0.78 0.53 0.88 ;
      RECT 0.43 0.55 0.53 0.65 ;
      RECT 0.43 0.35 0.53 0.45 ;
      RECT 0.7 1.79 0.8 1.89 ;
      RECT 0.7 1.59 0.8 1.69 ;
      RECT 0.7 1.39 0.8 1.49 ;
      RECT 0.7 0.55 0.8 0.65 ;
      RECT 0.7 0.35 0.8 0.45 ;
      RECT 1.06 1.04 1.16 1.14 ;
      RECT 1.41 1.79 1.51 1.89 ;
      RECT 1.41 1.59 1.51 1.69 ;
      RECT 1.41 1.39 1.51 1.49 ;
      RECT 1.41 0.55 1.51 0.65 ;
      RECT 1.41 0.35 1.51 0.45 ;
    LAYER ME2 ;
      RECT 0.43 0.32 0.53 1.92 ;
      RECT 0.7 1.04 1.19 1.14 ;
      RECT 0.7 0.32 0.8 1.92 ;
      RECT 1.41 0.32 1.51 1.92 ;
  END
END BUFENX2

MACRO BUFENX4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN BUFENX4 0 -0.11 ;
  SIZE 2.24 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.23 1.245 0.65 1.345 ;
    END
  END A
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.23 1.62 0.32 2.52 ;
        RECT 1.02 1.32 1.11 2.52 ;
        RECT 1.92 1.32 2.01 2.52 ;
        RECT 0 2.3 2.24 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.23 -0.22 0.32 0.53 ;
        RECT 1.02 -0.22 1.11 0.68 ;
        RECT 1.92 -0.22 2.01 0.68 ;
        RECT 0 -0.22 2.24 0 ;
    END
  END gnd!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.465 1.79 1.565 1.89 ;
        RECT 1.465 1.59 1.565 1.69 ;
        RECT 1.465 1.39 1.565 1.49 ;
        RECT 1.465 0.55 1.565 0.65 ;
        RECT 1.465 0.35 1.565 0.45 ;
      LAYER ME1 ;
        RECT 1.455 0.32 1.575 0.68 ;
        RECT 1.465 1.36 1.565 1.92 ;
        RECT 1.47 1.32 1.56 1.92 ;
      LAYER ME2 ;
        RECT 1.465 0.32 1.565 1.92 ;
    END
  END Y
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.575 0.985 0.995 1.085 ;
    END
  END EN
  OBS
    LAYER ME1 ;
      RECT 0.475 1.56 0.595 1.92 ;
      RECT 0.475 0.32 0.595 0.68 ;
      RECT 0.23 1.245 0.65 1.345 ;
      RECT 0.76 1.32 0.85 1.92 ;
      RECT 0.755 1.36 0.855 1.92 ;
      RECT 0.745 0.32 0.865 0.68 ;
      RECT 0.575 0.985 0.995 1.085 ;
      RECT 0.455 0.78 1.255 0.88 ;
      RECT 1.47 1.32 1.56 1.92 ;
      RECT 1.465 1.36 1.565 1.92 ;
      RECT 1.455 0.32 1.575 0.68 ;
      RECT 1.115 1.115 1.675 1.215 ;
      RECT 0.23 1.62 0.32 2.52 ;
      RECT 1.02 1.32 1.11 2.52 ;
      RECT 1.92 1.32 2.01 2.52 ;
      RECT 0 2.3 2.24 2.52 ;
      RECT 0 -0.22 2.24 0 ;
      RECT 0.23 -0.22 0.32 0.53 ;
      RECT 1.02 -0.22 1.11 0.68 ;
      RECT 1.92 -0.22 2.01 0.68 ;
    LAYER VI1 ;
      RECT 0.485 1.79 0.585 1.89 ;
      RECT 0.485 1.59 0.585 1.69 ;
      RECT 0.485 0.78 0.585 0.88 ;
      RECT 0.485 0.55 0.585 0.65 ;
      RECT 0.485 0.35 0.585 0.45 ;
      RECT 0.755 1.79 0.855 1.89 ;
      RECT 0.755 1.59 0.855 1.69 ;
      RECT 0.755 1.39 0.855 1.49 ;
      RECT 0.755 0.55 0.855 0.65 ;
      RECT 0.755 0.35 0.855 0.45 ;
      RECT 1.145 1.115 1.245 1.215 ;
      RECT 1.465 1.79 1.565 1.89 ;
      RECT 1.465 1.59 1.565 1.69 ;
      RECT 1.465 1.39 1.565 1.49 ;
      RECT 1.465 0.55 1.565 0.65 ;
      RECT 1.465 0.35 1.565 0.45 ;
    LAYER ME2 ;
      RECT 0.485 0.32 0.585 1.92 ;
      RECT 0.755 1.115 1.275 1.215 ;
      RECT 0.755 0.32 0.855 1.92 ;
      RECT 1.465 0.32 1.565 1.92 ;
  END
END BUFENX4

MACRO BUFX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN BUFX1 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.17 1.095 0.59 1.195 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.63 1.85 0.73 1.95 ;
        RECT 0.63 1.65 0.73 1.75 ;
        RECT 0.63 0.4 0.73 0.5 ;
        RECT 0.63 0.2 0.73 0.3 ;
      LAYER ME1 ;
        RECT 0.62 0.17 0.74 0.53 ;
        RECT 0.62 1.62 0.74 1.98 ;
      LAYER ME2 ;
        RECT 0.63 0.17 0.73 1.98 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.375 -0.22 0.465 0.53 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.375 1.62 0.465 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.1 1.62 0.22 1.98 ;
      RECT 0.1 0.17 0.22 0.53 ;
      RECT 0.17 1.095 0.59 1.195 ;
      RECT 0.08 1.35 0.64 1.45 ;
      RECT 0.62 1.62 0.74 1.98 ;
      RECT 0.62 0.17 0.74 0.53 ;
      RECT 0.375 1.62 0.465 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.375 -0.22 0.465 0.53 ;
    LAYER VI1 ;
      RECT 0.11 1.85 0.21 1.95 ;
      RECT 0.11 1.65 0.21 1.75 ;
      RECT 0.11 1.35 0.21 1.45 ;
      RECT 0.11 0.4 0.21 0.5 ;
      RECT 0.11 0.2 0.21 0.3 ;
      RECT 0.63 1.85 0.73 1.95 ;
      RECT 0.63 1.65 0.73 1.75 ;
      RECT 0.63 0.4 0.73 0.5 ;
      RECT 0.63 0.2 0.73 0.3 ;
    LAYER ME2 ;
      RECT 0.08 1.35 0.24 1.45 ;
      RECT 0.11 0.17 0.21 1.98 ;
      RECT 0.63 0.17 0.73 1.98 ;
  END
END BUFX1

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN BUFX2 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.13 0.875 0.55 0.975 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.63 1.79 0.73 1.89 ;
        RECT 0.63 1.59 0.73 1.69 ;
        RECT 0.63 1.39 0.73 1.49 ;
        RECT 0.63 0.55 0.73 0.65 ;
        RECT 0.63 0.35 0.73 0.45 ;
      LAYER ME1 ;
        RECT 0.62 0.32 0.74 0.68 ;
        RECT 0.63 1.36 0.73 1.92 ;
        RECT 0.635 1.32 0.725 1.92 ;
      LAYER ME2 ;
        RECT 0.63 0.32 0.73 1.92 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.375 -0.22 0.465 0.68 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.375 1.32 0.465 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.115 1.32 0.205 1.92 ;
      RECT 0.11 1.36 0.21 1.92 ;
      RECT 0.1 0.32 0.22 0.68 ;
      RECT 0.13 0.875 0.55 0.975 ;
      RECT 0.08 1.11 0.64 1.21 ;
      RECT 0.635 1.32 0.725 1.92 ;
      RECT 0.63 1.36 0.73 1.92 ;
      RECT 0.62 0.32 0.74 0.68 ;
      RECT 0.375 1.32 0.465 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.375 -0.22 0.465 0.68 ;
    LAYER VI1 ;
      RECT 0.11 1.79 0.21 1.89 ;
      RECT 0.11 1.59 0.21 1.69 ;
      RECT 0.11 1.39 0.21 1.49 ;
      RECT 0.11 1.11 0.21 1.21 ;
      RECT 0.11 0.55 0.21 0.65 ;
      RECT 0.11 0.35 0.21 0.45 ;
      RECT 0.63 1.79 0.73 1.89 ;
      RECT 0.63 1.59 0.73 1.69 ;
      RECT 0.63 1.39 0.73 1.49 ;
      RECT 0.63 0.55 0.73 0.65 ;
      RECT 0.63 0.35 0.73 0.45 ;
    LAYER ME2 ;
      RECT 0.11 0.32 0.21 1.92 ;
      RECT 0.63 0.32 0.73 1.92 ;
  END
END BUFX2

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN BUFX4 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.145 1.055 0.565 1.155 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.64 1.79 0.74 1.89 ;
        RECT 0.64 1.59 0.74 1.69 ;
        RECT 0.64 1.39 0.74 1.49 ;
        RECT 0.64 0.55 0.74 0.65 ;
        RECT 0.64 0.35 0.74 0.45 ;
      LAYER ME1 ;
        RECT 0.63 0.32 0.75 0.68 ;
        RECT 0.64 1.36 0.74 1.92 ;
        RECT 0.645 1.32 0.735 1.92 ;
      LAYER ME2 ;
        RECT 0.64 0.32 0.74 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.385 1.32 0.475 2.52 ;
        RECT 0.905 1.32 0.995 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.385 -0.22 0.475 0.68 ;
        RECT 0.905 -0.22 0.995 0.68 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.125 1.32 0.215 1.92 ;
      RECT 0.12 1.36 0.22 1.92 ;
      RECT 0.11 0.32 0.23 0.68 ;
      RECT 0.145 1.055 0.565 1.155 ;
      RECT 0.645 1.32 0.735 1.92 ;
      RECT 0.64 1.36 0.74 1.92 ;
      RECT 0.63 0.32 0.75 0.68 ;
      RECT 0.09 0.81 0.88 0.91 ;
      RECT 0.385 1.32 0.475 2.52 ;
      RECT 0.905 1.32 0.995 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.385 -0.22 0.475 0.68 ;
      RECT 0.905 -0.22 0.995 0.68 ;
    LAYER VI1 ;
      RECT 0.12 1.79 0.22 1.89 ;
      RECT 0.12 1.59 0.22 1.69 ;
      RECT 0.12 1.39 0.22 1.49 ;
      RECT 0.12 0.81 0.22 0.91 ;
      RECT 0.12 0.55 0.22 0.65 ;
      RECT 0.12 0.35 0.22 0.45 ;
      RECT 0.64 1.79 0.74 1.89 ;
      RECT 0.64 1.59 0.74 1.69 ;
      RECT 0.64 1.39 0.74 1.49 ;
      RECT 0.64 0.55 0.74 0.65 ;
      RECT 0.64 0.35 0.74 0.45 ;
    LAYER ME2 ;
      RECT 0.12 0.32 0.22 1.92 ;
      RECT 0.64 0.32 0.74 1.92 ;
  END
END BUFX4

MACRO FA1X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN FA1X1 0 -0.11 ;
  SIZE 5.6 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.47 -0.22 0.56 0.53 ;
        RECT 1.37 -0.22 1.46 0.53 ;
        RECT 2.38 -0.22 2.47 0.53 ;
        RECT 3.13 -0.22 3.22 0.53 ;
        RECT 4.14 -0.22 4.23 0.53 ;
        RECT 5.04 -0.22 5.13 0.53 ;
        RECT 0 -0.22 5.6 0 ;
    END
  END gnd!
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 2.705 1.1 4.375 1.2 ;
    END
  END CIN
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.47 1.62 0.56 2.52 ;
        RECT 1.37 1.62 1.46 2.52 ;
        RECT 1.86 1.62 1.95 2.52 ;
        RECT 2.38 1.62 2.47 2.52 ;
        RECT 2.9 1.62 2.99 2.52 ;
        RECT 3.13 1.62 3.22 2.52 ;
        RECT 3.65 1.62 3.74 2.52 ;
        RECT 4.14 1.62 4.23 2.52 ;
        RECT 5.04 1.62 5.13 2.52 ;
        RECT 0 2.3 5.6 2.52 ;
    END
  END vdd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.225 1.1 2.145 1.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.4 0.88 0.49 1.05 ;
        RECT 0.4 0.915 1.135 1.015 ;
        RECT 0.805 0.9 1.135 1.03 ;
        RECT 0.805 0.9 2.355 1 ;
        RECT 2.265 0.865 2.355 1.035 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 4.585 1.72 4.685 1.82 ;
        RECT 4.585 0.4 4.685 0.5 ;
      LAYER ME1 ;
        RECT 4.555 0.23 4.715 0.53 ;
        RECT 4.555 1.62 4.715 1.92 ;
      LAYER ME2 ;
        RECT 4.585 0.37 4.685 1.92 ;
    END
  END S
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 3.385 1.72 3.485 1.82 ;
        RECT 3.575 0.405 3.675 0.505 ;
      LAYER ME1 ;
        RECT 3.545 0.23 3.705 0.53 ;
        RECT 3.575 0.23 3.675 0.535 ;
        RECT 3.355 1.62 3.515 1.92 ;
      LAYER ME2 ;
        RECT 3.385 1.62 3.675 1.72 ;
        RECT 3.575 0.375 3.675 1.72 ;
        RECT 3.385 1.62 3.485 1.92 ;
    END
  END COUT
  OBS
    LAYER ME1 ;
      RECT 0.885 1.62 1.045 1.92 ;
      RECT 0.885 0.23 1.045 0.53 ;
      RECT 0.21 0.65 0.935 0.74 ;
      RECT 0.21 1.19 1.125 1.28 ;
      RECT 1.035 1.15 1.125 1.32 ;
      RECT 0.21 0.38 0.3 1.92 ;
      RECT 1.595 1.62 1.755 1.92 ;
      RECT 0.555 1.41 1.755 1.51 ;
      RECT 1.595 0.23 1.755 0.53 ;
      RECT 1.895 0.23 2.055 0.53 ;
      RECT 1.225 1.1 2.145 1.2 ;
      RECT 2.085 1.62 2.245 1.92 ;
      RECT 0.805 0.9 2.355 1 ;
      RECT 0.4 0.915 1.135 1.015 ;
      RECT 0.805 0.9 1.135 1.03 ;
      RECT 2.265 0.865 2.355 1.035 ;
      RECT 0.4 0.88 0.49 1.05 ;
      RECT 2.605 1.62 2.765 1.92 ;
      RECT 2.795 0.23 2.955 0.53 ;
      RECT 2.825 0.23 2.925 0.535 ;
      RECT 2.795 0.7 3.365 0.8 ;
      RECT 3.355 1.62 3.515 1.92 ;
      RECT 1.895 1.3 3.605 1.4 ;
      RECT 3.545 0.23 3.705 0.53 ;
      RECT 3.575 0.23 3.675 0.535 ;
      RECT 3.845 1.62 4.005 1.92 ;
      RECT 3.845 0.23 4.005 0.53 ;
      RECT 2.705 1.1 4.375 1.2 ;
      RECT 4.555 1.62 4.715 1.92 ;
      RECT 4.555 0.23 4.715 0.53 ;
      RECT 3.845 1.41 5.045 1.51 ;
      RECT 1.335 0.65 2.555 0.74 ;
      RECT 1.335 0.645 1.495 0.745 ;
      RECT 2.465 0.65 2.555 1 ;
      RECT 2.465 0.9 4.795 1 ;
      RECT 4.465 0.915 5.2 1.015 ;
      RECT 4.465 0.9 4.795 1.03 ;
      RECT 5.11 0.88 5.2 1.05 ;
      RECT 4.665 0.65 5.39 0.74 ;
      RECT 4.475 1.19 5.39 1.28 ;
      RECT 4.475 1.15 4.565 1.32 ;
      RECT 5.3 0.38 5.39 1.92 ;
      RECT 0.47 1.62 0.56 2.52 ;
      RECT 1.37 1.62 1.46 2.52 ;
      RECT 1.86 1.62 1.95 2.52 ;
      RECT 2.38 1.62 2.47 2.52 ;
      RECT 2.9 1.62 2.99 2.52 ;
      RECT 3.13 1.62 3.22 2.52 ;
      RECT 3.65 1.62 3.74 2.52 ;
      RECT 4.14 1.62 4.23 2.52 ;
      RECT 5.04 1.62 5.13 2.52 ;
      RECT 0 2.3 5.6 2.52 ;
      RECT 0 -0.22 5.6 0 ;
      RECT 0.47 -0.22 0.56 0.53 ;
      RECT 1.37 -0.22 1.46 0.53 ;
      RECT 2.38 -0.22 2.47 0.53 ;
      RECT 3.13 -0.22 3.22 0.53 ;
      RECT 4.14 -0.22 4.23 0.53 ;
      RECT 5.04 -0.22 5.13 0.53 ;
    LAYER VI1 ;
      RECT 0.915 1.72 1.015 1.82 ;
      RECT 0.915 0.4 1.015 0.5 ;
      RECT 1.365 0.645 1.465 0.745 ;
      RECT 1.625 1.72 1.725 1.82 ;
      RECT 1.625 1.41 1.725 1.51 ;
      RECT 1.625 0.4 1.725 0.5 ;
      RECT 1.925 1.3 2.025 1.4 ;
      RECT 1.925 0.4 2.025 0.5 ;
      RECT 2.115 1.72 2.215 1.82 ;
      RECT 2.635 1.72 2.735 1.82 ;
      RECT 2.825 0.7 2.925 0.8 ;
      RECT 2.825 0.405 2.925 0.505 ;
      RECT 3.385 1.72 3.485 1.82 ;
      RECT 3.575 0.405 3.675 0.505 ;
      RECT 3.875 1.72 3.975 1.82 ;
      RECT 3.875 1.41 3.975 1.51 ;
      RECT 3.875 0.4 3.975 0.5 ;
      RECT 4.585 1.72 4.685 1.82 ;
      RECT 4.585 0.4 4.685 0.5 ;
    LAYER ME2 ;
      RECT 0.915 0.645 1.495 0.745 ;
      RECT 0.915 0.37 1.015 1.92 ;
      RECT 1.625 0.37 1.725 1.92 ;
      RECT 1.925 0.37 2.025 1.72 ;
      RECT 1.925 1.62 2.215 1.72 ;
      RECT 2.115 1.62 2.215 1.92 ;
      RECT 2.825 0.23 2.925 1.72 ;
      RECT 2.635 1.62 2.925 1.72 ;
      RECT 2.635 1.62 2.735 1.92 ;
      RECT 3.575 0.375 3.675 1.72 ;
      RECT 3.385 1.62 3.675 1.72 ;
      RECT 3.385 1.62 3.485 1.92 ;
      RECT 3.875 0.37 3.975 1.92 ;
      RECT 4.585 0.37 4.685 1.92 ;
  END
END FA1X1

MACRO FILL1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN FILL1 0 -0.11 ;
  SIZE 0.28 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.22 0.28 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 2.3 0.28 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0 2.3 0.28 2.52 ;
      RECT 0 -0.22 0.28 0 ;
  END
END FILL1

MACRO FILL2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN FILL2 0 -0.11 ;
  SIZE 0.56 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.22 0.56 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 2.3 0.56 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0 2.3 0.56 2.52 ;
      RECT 0 -0.22 0.56 0 ;
  END
END FILL2

MACRO FILL3
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN FILL3 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
  END
END FILL3

MACRO FILL4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN FILL4 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
  END
END FILL4

MACRO HA1X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN HA1X1 0 -0.11 ;
  SIZE 2.8 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.44 0.9 2.065 1 ;
        RECT 1.735 0.9 2.065 1.03 ;
        RECT 1.735 0.915 2.47 1.015 ;
        RECT 2.38 0.88 2.47 1.05 ;
    END
  END B
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.4 -0.22 0.49 0.53 ;
        RECT 1.41 -0.22 1.5 0.53 ;
        RECT 2.31 -0.22 2.4 0.53 ;
        RECT 0 -0.22 2.8 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.4 1.62 0.49 2.52 ;
        RECT 0.92 1.62 1.01 2.52 ;
        RECT 1.41 1.62 1.5 2.52 ;
        RECT 2.31 1.62 2.4 2.52 ;
        RECT 0 2.3 2.8 2.52 ;
    END
  END vdd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.49 1.1 1.645 1.2 ;
    END
  END A
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.855 1.72 1.955 1.82 ;
        RECT 1.855 0.4 1.955 0.5 ;
      LAYER ME1 ;
        RECT 1.825 0.23 1.985 0.53 ;
        RECT 1.825 1.62 1.985 1.92 ;
      LAYER ME2 ;
        RECT 1.855 0.37 1.955 1.92 ;
    END
  END S
  PIN C
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.135 1.85 0.235 1.95 ;
        RECT 0.135 1.65 0.235 1.75 ;
        RECT 0.135 0.4 0.235 0.5 ;
        RECT 0.135 0.2 0.235 0.3 ;
      LAYER ME1 ;
        RECT 0.125 0.17 0.245 0.53 ;
        RECT 0.125 1.62 0.245 1.98 ;
      LAYER ME2 ;
        RECT 0.135 0.17 0.235 1.98 ;
    END
  END C
  OBS
    LAYER ME1 ;
      RECT 0.125 1.62 0.245 1.98 ;
      RECT 0.125 0.17 0.245 0.53 ;
      RECT 0.645 1.62 0.765 1.98 ;
      RECT 0.835 0.17 0.955 0.53 ;
      RECT 0.255 1.39 0.975 1.49 ;
      RECT 1.115 1.62 1.275 1.92 ;
      RECT 1.115 0.23 1.275 0.53 ;
      RECT 0.49 1.1 1.645 1.2 ;
      RECT 1.825 1.62 1.985 1.92 ;
      RECT 1.825 0.23 1.985 0.53 ;
      RECT 1.115 1.41 2.315 1.51 ;
      RECT 0.44 0.9 2.065 1 ;
      RECT 1.735 0.915 2.47 1.015 ;
      RECT 1.735 0.9 2.065 1.03 ;
      RECT 2.38 0.88 2.47 1.05 ;
      RECT 1.935 0.65 2.66 0.74 ;
      RECT 1.745 1.19 2.66 1.28 ;
      RECT 1.745 1.15 1.835 1.32 ;
      RECT 2.57 0.38 2.66 1.92 ;
      RECT 0.4 1.62 0.49 2.52 ;
      RECT 0.92 1.62 1.01 2.52 ;
      RECT 1.41 1.62 1.5 2.52 ;
      RECT 2.31 1.62 2.4 2.52 ;
      RECT 0 2.3 2.8 2.52 ;
      RECT 0 -0.22 2.8 0 ;
      RECT 0.4 -0.22 0.49 0.53 ;
      RECT 1.41 -0.22 1.5 0.53 ;
      RECT 2.31 -0.22 2.4 0.53 ;
    LAYER VI1 ;
      RECT 0.135 1.85 0.235 1.95 ;
      RECT 0.135 1.65 0.235 1.75 ;
      RECT 0.135 0.4 0.235 0.5 ;
      RECT 0.135 0.2 0.235 0.3 ;
      RECT 0.655 1.85 0.755 1.95 ;
      RECT 0.655 1.65 0.755 1.75 ;
      RECT 0.845 1.39 0.945 1.49 ;
      RECT 0.845 0.4 0.945 0.5 ;
      RECT 0.845 0.2 0.945 0.3 ;
      RECT 1.145 1.72 1.245 1.82 ;
      RECT 1.145 1.41 1.245 1.51 ;
      RECT 1.145 0.4 1.245 0.5 ;
      RECT 1.855 1.72 1.955 1.82 ;
      RECT 1.855 0.4 1.955 0.5 ;
    LAYER ME2 ;
      RECT 0.135 0.17 0.235 1.98 ;
      RECT 0.815 1.39 0.975 1.49 ;
      RECT 0.845 0.17 0.945 1.72 ;
      RECT 0.655 1.62 0.945 1.72 ;
      RECT 0.655 1.62 0.755 1.98 ;
      RECT 1.145 0.37 1.245 1.92 ;
      RECT 1.855 0.37 1.955 1.92 ;
  END
END HA1X1

MACRO HACB1X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN HACB1X1 0 -0.11 ;
  SIZE 2.52 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.205 0.9 1.785 1 ;
        RECT 1.455 0.9 1.785 1.03 ;
        RECT 1.455 0.915 2.19 1.015 ;
        RECT 2.1 0.88 2.19 1.05 ;
    END
  END B
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.12 -0.22 0.21 0.53 ;
        RECT 1.13 -0.22 1.22 0.53 ;
        RECT 2.03 -0.22 2.12 0.53 ;
        RECT 0 -0.22 2.52 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.12 1.62 0.21 2.52 ;
        RECT 0.64 1.62 0.73 2.52 ;
        RECT 1.13 1.62 1.22 2.52 ;
        RECT 2.03 1.62 2.12 2.52 ;
        RECT 0 2.3 2.52 2.52 ;
    END
  END vdd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.205 1.1 1.365 1.2 ;
    END
  END A
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.575 1.72 1.675 1.82 ;
        RECT 1.575 0.4 1.675 0.5 ;
      LAYER ME1 ;
        RECT 1.545 0.23 1.705 0.53 ;
        RECT 1.545 1.62 1.705 1.92 ;
      LAYER ME2 ;
        RECT 1.575 0.37 1.675 1.92 ;
    END
  END S
  PIN CB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.375 1.85 0.475 1.95 ;
        RECT 0.375 1.65 0.475 1.75 ;
        RECT 0.565 0.4 0.665 0.5 ;
        RECT 0.565 0.2 0.665 0.3 ;
      LAYER ME1 ;
        RECT 0.555 0.17 0.675 0.53 ;
        RECT 0.365 1.62 0.485 1.98 ;
      LAYER ME2 ;
        RECT 0.375 1.62 0.665 1.72 ;
        RECT 0.565 0.17 0.665 1.72 ;
        RECT 0.375 1.62 0.475 1.98 ;
    END
  END CB
  OBS
    LAYER ME1 ;
      RECT 0.365 1.62 0.485 1.98 ;
      RECT 0.555 0.17 0.675 0.53 ;
      RECT 0.835 1.62 0.995 1.92 ;
      RECT 0.835 0.23 0.995 0.53 ;
      RECT 0.205 1.1 1.365 1.2 ;
      RECT 1.545 1.62 1.705 1.92 ;
      RECT 1.545 0.23 1.705 0.53 ;
      RECT 0.835 1.41 2.035 1.51 ;
      RECT 0.205 0.9 1.785 1 ;
      RECT 1.455 0.915 2.19 1.015 ;
      RECT 1.455 0.9 1.785 1.03 ;
      RECT 2.1 0.88 2.19 1.05 ;
      RECT 1.655 0.65 2.38 0.74 ;
      RECT 1.465 1.19 2.38 1.28 ;
      RECT 1.465 1.15 1.555 1.32 ;
      RECT 2.29 0.38 2.38 1.92 ;
      RECT 0.12 1.62 0.21 2.52 ;
      RECT 0.64 1.62 0.73 2.52 ;
      RECT 1.13 1.62 1.22 2.52 ;
      RECT 2.03 1.62 2.12 2.52 ;
      RECT 0 2.3 2.52 2.52 ;
      RECT 0 -0.22 2.52 0 ;
      RECT 0.12 -0.22 0.21 0.53 ;
      RECT 1.13 -0.22 1.22 0.53 ;
      RECT 2.03 -0.22 2.12 0.53 ;
    LAYER VI1 ;
      RECT 0.375 1.85 0.475 1.95 ;
      RECT 0.375 1.65 0.475 1.75 ;
      RECT 0.565 0.4 0.665 0.5 ;
      RECT 0.565 0.2 0.665 0.3 ;
      RECT 0.865 1.72 0.965 1.82 ;
      RECT 0.865 1.41 0.965 1.51 ;
      RECT 0.865 0.4 0.965 0.5 ;
      RECT 1.575 1.72 1.675 1.82 ;
      RECT 1.575 0.4 1.675 0.5 ;
    LAYER ME2 ;
      RECT 0.565 0.17 0.665 1.72 ;
      RECT 0.375 1.62 0.665 1.72 ;
      RECT 0.375 1.62 0.475 1.98 ;
      RECT 0.865 0.37 0.965 1.92 ;
      RECT 1.575 0.37 1.675 1.92 ;
  END
END HACB1X1

MACRO INVENX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN INVENX1 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.265 1.145 0.685 1.245 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.865 1.85 0.965 1.95 ;
        RECT 0.865 1.65 0.965 1.75 ;
        RECT 0.865 0.4 0.965 0.5 ;
        RECT 0.865 0.2 0.965 0.3 ;
      LAYER ME1 ;
        RECT 0.855 0.17 0.975 0.53 ;
        RECT 0.855 1.62 0.975 1.98 ;
      LAYER ME2 ;
        RECT 0.865 0.17 0.965 1.98 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.42 1.62 0.51 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.145 0.945 0.565 1.045 ;
    END
  END EN
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.42 -0.22 0.51 0.53 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.145 1.62 0.265 1.98 ;
      RECT 0.145 0.17 0.265 0.53 ;
      RECT 0.145 0.945 0.565 1.045 ;
      RECT 0.265 1.145 0.685 1.245 ;
      RECT 0.125 1.41 0.875 1.52 ;
      RECT 0.855 1.62 0.975 1.98 ;
      RECT 0.855 0.17 0.975 0.53 ;
      RECT 0.42 1.62 0.51 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.42 -0.22 0.51 0.53 ;
    LAYER VI1 ;
      RECT 0.155 1.85 0.255 1.95 ;
      RECT 0.155 1.65 0.255 1.75 ;
      RECT 0.155 1.415 0.255 1.515 ;
      RECT 0.155 0.4 0.255 0.5 ;
      RECT 0.155 0.2 0.255 0.3 ;
      RECT 0.865 1.85 0.965 1.95 ;
      RECT 0.865 1.65 0.965 1.75 ;
      RECT 0.865 0.4 0.965 0.5 ;
      RECT 0.865 0.2 0.965 0.3 ;
    LAYER ME2 ;
      RECT 0.155 0.17 0.255 1.98 ;
      RECT 0.865 0.17 0.965 1.98 ;
  END
END INVENX1

MACRO INVENX2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN INVENX2 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.855 1.79 0.955 1.89 ;
        RECT 0.855 1.59 0.955 1.69 ;
        RECT 0.855 1.39 0.955 1.49 ;
        RECT 0.855 0.55 0.955 0.65 ;
        RECT 0.855 0.35 0.955 0.45 ;
      LAYER ME2 ;
        RECT 0.855 0.32 0.955 1.92 ;
      LAYER ME1 ;
        RECT 0.845 0.32 0.965 0.68 ;
        RECT 0.855 1.36 0.955 1.92 ;
        RECT 0.86 1.32 0.95 1.92 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.495 0.925 0.915 1.025 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.115 0.83 0.395 0.98 ;
    END
  END EN
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.41 -0.22 0.5 0.68 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.41 1.32 0.5 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.15 1.32 0.24 1.92 ;
      RECT 0.145 1.36 0.245 1.92 ;
      RECT 0.135 0.32 0.255 0.68 ;
      RECT 0.115 0.83 0.395 0.98 ;
      RECT 0.115 1.125 0.915 1.225 ;
      RECT 0.495 0.925 0.915 1.025 ;
      RECT 0.86 1.32 0.95 1.92 ;
      RECT 0.855 1.36 0.955 1.92 ;
      RECT 0.845 0.32 0.965 0.68 ;
      RECT 0.41 1.32 0.5 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.41 -0.22 0.5 0.68 ;
    LAYER VI1 ;
      RECT 0.145 1.79 0.245 1.89 ;
      RECT 0.145 1.59 0.245 1.69 ;
      RECT 0.145 1.39 0.245 1.49 ;
      RECT 0.145 1.125 0.245 1.225 ;
      RECT 0.145 0.55 0.245 0.65 ;
      RECT 0.145 0.35 0.245 0.45 ;
      RECT 0.855 1.79 0.955 1.89 ;
      RECT 0.855 1.59 0.955 1.69 ;
      RECT 0.855 1.39 0.955 1.49 ;
      RECT 0.855 0.55 0.955 0.65 ;
      RECT 0.855 0.35 0.955 0.45 ;
    LAYER ME2 ;
      RECT 0.145 0.32 0.245 1.92 ;
      RECT 0.855 0.32 0.955 1.92 ;
  END
END INVENX2

MACRO INVENX4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN INVENX4 0 -0.11 ;
  SIZE 1.68 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.475 1.32 0.565 2.52 ;
        RECT 1.375 1.32 1.465 2.52 ;
        RECT 0 2.3 1.68 2.52 ;
    END
  END vdd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.045 0.915 1.465 1.015 ;
    END
  END A
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.475 -0.22 0.565 0.68 ;
        RECT 1.375 -0.22 1.465 0.68 ;
        RECT 0 -0.22 1.68 0 ;
    END
  END gnd!
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.18 0.915 0.6 1.015 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.92 1.79 1.02 1.89 ;
        RECT 0.92 1.59 1.02 1.69 ;
        RECT 0.92 1.39 1.02 1.49 ;
        RECT 0.92 0.55 1.02 0.65 ;
        RECT 0.92 0.35 1.02 0.45 ;
      LAYER ME1 ;
        RECT 0.91 0.32 1.03 0.68 ;
        RECT 0.92 1.36 1.02 1.92 ;
        RECT 0.925 1.32 1.015 1.92 ;
      LAYER ME2 ;
        RECT 0.92 0.32 1.02 1.92 ;
    END
  END Y
  OBS
    LAYER ME1 ;
      RECT 0.215 1.32 0.305 1.92 ;
      RECT 0.21 1.36 0.31 1.92 ;
      RECT 0.2 0.32 0.32 0.68 ;
      RECT 0.18 0.915 0.6 1.015 ;
      RECT 0.18 1.12 0.98 1.22 ;
      RECT 0.925 1.32 1.015 1.92 ;
      RECT 0.92 1.36 1.02 1.92 ;
      RECT 0.91 0.32 1.03 0.68 ;
      RECT 1.045 0.915 1.465 1.015 ;
      RECT 0.475 1.32 0.565 2.52 ;
      RECT 1.375 1.32 1.465 2.52 ;
      RECT 0 2.3 1.68 2.52 ;
      RECT 0 -0.22 1.68 0 ;
      RECT 0.475 -0.22 0.565 0.68 ;
      RECT 1.375 -0.22 1.465 0.68 ;
    LAYER VI1 ;
      RECT 0.21 1.79 0.31 1.89 ;
      RECT 0.21 1.59 0.31 1.69 ;
      RECT 0.21 1.39 0.31 1.49 ;
      RECT 0.21 1.12 0.31 1.22 ;
      RECT 0.21 0.55 0.31 0.65 ;
      RECT 0.21 0.35 0.31 0.45 ;
      RECT 0.92 1.79 1.02 1.89 ;
      RECT 0.92 1.59 1.02 1.69 ;
      RECT 0.92 1.39 1.02 1.49 ;
      RECT 0.92 0.55 1.02 0.65 ;
      RECT 0.92 0.35 1.02 0.45 ;
    LAYER ME2 ;
      RECT 0.21 0.32 0.31 1.92 ;
      RECT 0.92 0.32 1.02 1.92 ;
  END
END INVENX4

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN INVX1 0 -0.11 ;
  SIZE 0.56 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.105 0.98 0.465 1.1 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.36 1.85 0.46 1.95 ;
        RECT 0.36 1.65 0.46 1.75 ;
        RECT 0.36 0.4 0.46 0.5 ;
        RECT 0.36 0.2 0.46 0.3 ;
      LAYER ME1 ;
        RECT 0.35 0.17 0.47 0.53 ;
        RECT 0.35 1.62 0.47 1.98 ;
      LAYER ME2 ;
        RECT 0.36 0.17 0.46 1.98 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 -0.22 0.195 0.53 ;
        RECT 0 -0.22 0.56 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 1.62 0.195 2.52 ;
        RECT 0 2.3 0.56 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.105 0.98 0.465 1.1 ;
      RECT 0.35 1.62 0.47 1.98 ;
      RECT 0.35 0.17 0.47 0.53 ;
      RECT 0.105 1.62 0.195 2.52 ;
      RECT 0 2.3 0.56 2.52 ;
      RECT 0 -0.22 0.56 0 ;
      RECT 0.105 -0.22 0.195 0.53 ;
    LAYER VI1 ;
      RECT 0.36 1.85 0.46 1.95 ;
      RECT 0.36 1.65 0.46 1.75 ;
      RECT 0.36 0.4 0.46 0.5 ;
      RECT 0.36 0.2 0.46 0.3 ;
    LAYER ME2 ;
      RECT 0.36 0.17 0.46 1.98 ;
  END
END INVX1

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN INVX2 0 -0.11 ;
  SIZE 0.56 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.1 0.84 0.46 0.96 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.36 1.79 0.46 1.89 ;
        RECT 0.36 1.59 0.46 1.69 ;
        RECT 0.36 1.39 0.46 1.49 ;
        RECT 0.36 0.55 0.46 0.65 ;
        RECT 0.36 0.35 0.46 0.45 ;
      LAYER ME1 ;
        RECT 0.35 0.32 0.47 0.68 ;
        RECT 0.36 1.36 0.46 1.92 ;
        RECT 0.365 1.32 0.455 1.92 ;
      LAYER ME2 ;
        RECT 0.36 0.32 0.46 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 1.32 0.195 2.52 ;
        RECT 0 2.3 0.56 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 -0.22 0.195 0.68 ;
        RECT 0 -0.22 0.56 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.365 1.32 0.455 1.92 ;
      RECT 0.36 1.36 0.46 1.92 ;
      RECT 0.1 0.84 0.46 0.96 ;
      RECT 0.35 0.32 0.47 0.68 ;
      RECT 0.105 1.32 0.195 2.52 ;
      RECT 0 2.3 0.56 2.52 ;
      RECT 0 -0.22 0.56 0 ;
      RECT 0.105 -0.22 0.195 0.68 ;
    LAYER VI1 ;
      RECT 0.36 1.79 0.46 1.89 ;
      RECT 0.36 1.59 0.46 1.69 ;
      RECT 0.36 1.39 0.46 1.49 ;
      RECT 0.36 0.55 0.46 0.65 ;
      RECT 0.36 0.35 0.46 0.45 ;
    LAYER ME2 ;
      RECT 0.36 0.32 0.46 1.92 ;
  END
END INVX2

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN INVX4 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.145 0.835 0.565 0.935 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.37 1.79 0.47 1.89 ;
        RECT 0.37 1.59 0.47 1.69 ;
        RECT 0.37 1.39 0.47 1.49 ;
        RECT 0.37 0.55 0.47 0.65 ;
        RECT 0.37 0.35 0.47 0.45 ;
      LAYER ME1 ;
        RECT 0.36 0.32 0.48 0.68 ;
        RECT 0.37 1.36 0.47 1.92 ;
        RECT 0.375 1.32 0.465 1.92 ;
      LAYER ME2 ;
        RECT 0.37 0.32 0.47 1.92 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 -0.22 0.205 0.68 ;
        RECT 0.635 -0.22 0.725 0.68 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 1.32 0.205 2.52 ;
        RECT 0.635 1.32 0.725 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.375 1.32 0.465 1.92 ;
      RECT 0.37 1.36 0.47 1.92 ;
      RECT 0.36 0.32 0.48 0.68 ;
      RECT 0.145 0.835 0.565 0.935 ;
      RECT 0.115 1.32 0.205 2.52 ;
      RECT 0.635 1.32 0.725 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.115 -0.22 0.205 0.68 ;
      RECT 0.635 -0.22 0.725 0.68 ;
    LAYER VI1 ;
      RECT 0.37 1.79 0.47 1.89 ;
      RECT 0.37 1.59 0.47 1.69 ;
      RECT 0.37 1.39 0.47 1.49 ;
      RECT 0.37 0.55 0.47 0.65 ;
      RECT 0.37 0.35 0.47 0.45 ;
    LAYER ME2 ;
      RECT 0.37 0.32 0.47 1.92 ;
  END
END INVX4

MACRO MUX2BX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN MUX2BX1 0 -0.11 ;
  SIZE 1.68 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.3 0.915 1.13 1.015 ;
        RECT 0.8 0.9 1.13 1.03 ;
    END
  END S
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.475 1.62 0.565 2.52 ;
        RECT 1.375 1.62 1.465 2.52 ;
        RECT 0 2.3 1.68 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.475 -0.22 0.565 0.53 ;
        RECT 1.375 -0.22 1.465 0.53 ;
        RECT 0 -0.22 1.68 0 ;
    END
  END gnd!
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.33 1.145 0.75 1.245 ;
    END
  END D0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.92 1.72 1.02 1.82 ;
        RECT 0.92 0.4 1.02 0.5 ;
      LAYER ME1 ;
        RECT 0.89 0.23 1.05 0.53 ;
        RECT 0.89 1.62 1.05 1.92 ;
      LAYER ME2 ;
        RECT 0.92 0.37 1.02 1.92 ;
    END
  END Y
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.995 1.205 1.415 1.305 ;
    END
  END D1
  OBS
    LAYER ME1 ;
      RECT 0.18 1.62 0.34 1.92 ;
      RECT 0.18 0.23 0.34 0.53 ;
      RECT 0.33 1.145 0.75 1.245 ;
      RECT 0.18 1.39 0.94 1.49 ;
      RECT 0.89 1.62 1.05 1.92 ;
      RECT 0.89 0.23 1.05 0.53 ;
      RECT 0.3 0.915 1.13 1.015 ;
      RECT 0.8 0.9 1.13 1.03 ;
      RECT 0.18 0.645 1.16 0.745 ;
      RECT 0.995 1.205 1.415 1.305 ;
      RECT 0.475 1.62 0.565 2.52 ;
      RECT 1.375 1.62 1.465 2.52 ;
      RECT 0 2.3 1.68 2.52 ;
      RECT 0 -0.22 1.68 0 ;
      RECT 0.475 -0.22 0.565 0.53 ;
      RECT 1.375 -0.22 1.465 0.53 ;
    LAYER VI1 ;
      RECT 0.21 1.72 0.31 1.82 ;
      RECT 0.21 1.39 0.31 1.49 ;
      RECT 0.21 0.645 0.31 0.745 ;
      RECT 0.21 0.4 0.31 0.5 ;
      RECT 0.92 1.72 1.02 1.82 ;
      RECT 0.92 0.4 1.02 0.5 ;
    LAYER ME2 ;
      RECT 0.21 0.37 0.31 1.92 ;
      RECT 0.92 0.37 1.02 1.92 ;
  END
END MUX2BX1

MACRO MUX2X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN MUX2X1 0 -0.11 ;
  SIZE 1.96 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.26 0.915 1.14 1.015 ;
        RECT 0.81 0.9 1.14 1.03 ;
    END
  END S
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 1.62 0.575 2.52 ;
        RECT 1.385 1.62 1.475 2.52 ;
        RECT 0 2.3 1.96 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 -0.22 0.575 0.53 ;
        RECT 1.385 -0.22 1.475 0.53 ;
        RECT 0 -0.22 1.96 0 ;
    END
  END gnd!
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.34 1.145 0.76 1.245 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.21 1.205 1.63 1.305 ;
    END
  END D1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.64 1.72 1.74 1.82 ;
        RECT 1.64 0.4 1.74 0.5 ;
      LAYER ME1 ;
        RECT 1.61 0.23 1.77 0.53 ;
        RECT 1.61 1.62 1.77 1.92 ;
      LAYER ME2 ;
        RECT 1.64 0.23 1.74 1.92 ;
    END
  END Y
  OBS
    LAYER ME1 ;
      RECT 0.19 1.62 0.35 1.92 ;
      RECT 0.19 0.23 0.35 0.53 ;
      RECT 0.34 1.145 0.76 1.245 ;
      RECT 0.19 1.39 0.95 1.49 ;
      RECT 0.9 1.62 1.06 1.92 ;
      RECT 0.9 0.23 1.06 0.53 ;
      RECT 0.26 0.915 1.14 1.015 ;
      RECT 0.81 0.9 1.14 1.03 ;
      RECT 0.19 0.635 1.155 0.735 ;
      RECT 1.21 1.205 1.63 1.305 ;
      RECT 1.24 0.915 1.71 1.015 ;
      RECT 1.61 1.62 1.77 1.92 ;
      RECT 1.61 0.23 1.77 0.53 ;
      RECT 0.485 1.62 0.575 2.52 ;
      RECT 1.385 1.62 1.475 2.52 ;
      RECT 0 2.3 1.96 2.52 ;
      RECT 0 -0.22 1.96 0 ;
      RECT 0.485 -0.22 0.575 0.53 ;
      RECT 1.385 -0.22 1.475 0.53 ;
    LAYER VI1 ;
      RECT 0.22 1.72 0.32 1.82 ;
      RECT 0.22 1.39 0.32 1.49 ;
      RECT 0.22 0.635 0.32 0.735 ;
      RECT 0.22 0.4 0.32 0.5 ;
      RECT 0.93 1.72 1.03 1.82 ;
      RECT 0.93 0.4 1.03 0.5 ;
      RECT 1.345 0.915 1.445 1.015 ;
      RECT 1.64 1.72 1.74 1.82 ;
      RECT 1.64 0.4 1.74 0.5 ;
    LAYER ME2 ;
      RECT 0.22 0.37 0.32 1.92 ;
      RECT 0.93 0.915 1.475 1.015 ;
      RECT 0.93 0.37 1.03 1.92 ;
      RECT 1.64 0.23 1.74 1.92 ;
  END
END MUX2X1

MACRO MUX4X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN MUX4X1 0 -0.11 ;
  SIZE 3.64 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 2.095 0.88 2.345 1.05 ;
    END
  END D2
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 3.175 1.405 3.275 1.505 ;
        RECT 3.175 0.645 3.275 0.745 ;
      LAYER ME1 ;
        RECT 2.76 1.405 3.39 1.505 ;
        RECT 2.53 0.645 3.305 0.745 ;
      LAYER ME2 ;
        RECT 3.175 0.615 3.275 1.535 ;
    END
  END S1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.32 1.42 1.42 1.52 ;
        RECT 1.32 0.915 1.42 1.015 ;
      LAYER ME1 ;
        RECT 1.29 1.42 2.01 1.52 ;
        RECT 1.32 0.645 1.79 0.745 ;
        RECT 0.25 0.915 1.45 1.015 ;
        RECT 1.32 0.645 1.42 1.015 ;
        RECT 0.75 0.9 1.08 1.03 ;
      LAYER ME2 ;
        RECT 1.32 0.885 1.42 1.55 ;
    END
  END S0
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.425 1.62 0.515 2.52 ;
        RECT 1.325 1.62 1.415 2.52 ;
        RECT 2.225 1.62 2.315 2.52 ;
        RECT 3.125 1.62 3.215 2.52 ;
        RECT 0 2.3 3.64 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.425 -0.22 0.515 0.53 ;
        RECT 1.325 -0.22 1.415 0.53 ;
        RECT 2.225 -0.22 2.315 0.53 ;
        RECT 3.125 -0.22 3.215 0.53 ;
        RECT 0 -0.22 3.64 0 ;
    END
  END gnd!
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.44 1.15 1.53 1.32 ;
        RECT 1.44 1.185 1.86 1.285 ;
    END
  END D3
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.91 1.19 1.33 1.29 ;
    END
  END D0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 2.67 1.72 2.77 1.82 ;
        RECT 2.67 0.4 2.77 0.5 ;
      LAYER ME1 ;
        RECT 2.64 0.23 2.8 0.53 ;
        RECT 2.64 1.62 2.8 1.92 ;
      LAYER ME2 ;
        RECT 2.67 0.37 2.77 1.92 ;
    END
  END Y
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.28 1.145 0.7 1.245 ;
    END
  END D1
  OBS
    LAYER ME1 ;
      RECT 0.13 1.62 0.29 1.92 ;
      RECT 0.13 0.23 0.29 0.53 ;
      RECT 0.28 1.145 0.7 1.245 ;
      RECT 0.13 1.39 0.88 1.49 ;
      RECT 0.84 1.62 1 1.92 ;
      RECT 0.84 0.23 1 0.53 ;
      RECT 0.13 0.645 1.23 0.745 ;
      RECT 0.91 1.19 1.33 1.29 ;
      RECT 1.32 0.645 1.79 0.745 ;
      RECT 1.32 0.645 1.42 1.015 ;
      RECT 0.25 0.915 1.45 1.015 ;
      RECT 0.75 0.9 1.08 1.03 ;
      RECT 1.44 1.185 1.86 1.285 ;
      RECT 1.44 1.15 1.53 1.32 ;
      RECT 1.74 1.62 1.9 1.92 ;
      RECT 1.74 0.23 1.9 0.53 ;
      RECT 1.56 0.87 1.66 1.03 ;
      RECT 1.56 0.9 1.99 1.03 ;
      RECT 1.29 1.42 2.01 1.52 ;
      RECT 2.095 0.88 2.345 1.05 ;
      RECT 2.275 1.205 2.695 1.305 ;
      RECT 2.64 1.62 2.8 1.92 ;
      RECT 2.64 0.23 2.8 0.53 ;
      RECT 2.53 0.645 3.305 0.745 ;
      RECT 2.935 1.145 3.36 1.245 ;
      RECT 2.76 1.405 3.39 1.505 ;
      RECT 3.35 1.62 3.51 1.92 ;
      RECT 2.56 0.915 3.51 1.015 ;
      RECT 2.56 0.9 2.89 1.03 ;
      RECT 3.35 0.23 3.51 0.53 ;
      RECT 0.425 1.62 0.515 2.52 ;
      RECT 1.325 1.62 1.415 2.52 ;
      RECT 2.225 1.62 2.315 2.52 ;
      RECT 3.125 1.62 3.215 2.52 ;
      RECT 0 2.3 3.64 2.52 ;
      RECT 0 -0.22 3.64 0 ;
      RECT 0.425 -0.22 0.515 0.53 ;
      RECT 1.325 -0.22 1.415 0.53 ;
      RECT 2.225 -0.22 2.315 0.53 ;
      RECT 3.125 -0.22 3.215 0.53 ;
    LAYER VI1 ;
      RECT 0.16 1.72 0.26 1.82 ;
      RECT 0.16 1.39 0.26 1.49 ;
      RECT 0.16 0.645 0.26 0.745 ;
      RECT 0.16 0.4 0.26 0.5 ;
      RECT 0.87 1.72 0.97 1.82 ;
      RECT 0.87 0.4 0.97 0.5 ;
      RECT 1.1 0.645 1.2 0.745 ;
      RECT 1.32 1.42 1.42 1.52 ;
      RECT 1.32 0.915 1.42 1.015 ;
      RECT 1.56 0.9 1.66 1 ;
      RECT 1.77 1.72 1.87 1.82 ;
      RECT 1.77 0.4 1.87 0.5 ;
      RECT 2.335 1.205 2.435 1.305 ;
      RECT 2.67 1.72 2.77 1.82 ;
      RECT 2.67 0.4 2.77 0.5 ;
      RECT 2.965 1.145 3.065 1.245 ;
      RECT 3.175 1.405 3.275 1.505 ;
      RECT 3.175 0.645 3.275 0.745 ;
      RECT 3.38 1.72 3.48 1.82 ;
      RECT 3.38 0.915 3.48 1.015 ;
      RECT 3.38 0.4 3.48 0.5 ;
    LAYER ME2 ;
      RECT 0.16 0.37 0.26 1.92 ;
      RECT 1.32 0.885 1.42 1.55 ;
      RECT 1.07 0.645 1.66 0.745 ;
      RECT 1.56 0.645 1.66 1.03 ;
      RECT 1.77 1.205 2.465 1.305 ;
      RECT 1.77 0.37 1.87 1.92 ;
      RECT 2.67 0.37 2.77 1.92 ;
      RECT 0.87 0.16 3.065 0.26 ;
      RECT 2.965 0.16 3.065 1.275 ;
      RECT 0.87 0.16 0.97 1.92 ;
      RECT 3.175 0.615 3.275 1.535 ;
      RECT 3.38 0.37 3.48 1.92 ;
  END
END MUX4X1

MACRO NAND2ALTX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN NAND2ALTX1 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.275 1.07 0.695 1.17 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.225 0.83 0.645 0.93 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.11 1.85 0.21 1.95 ;
        RECT 0.11 1.65 0.21 1.75 ;
        RECT 0.63 1.85 0.73 1.95 ;
        RECT 0.63 1.65 0.73 1.75 ;
        RECT 0.63 0.4 0.73 0.5 ;
        RECT 0.63 0.2 0.73 0.3 ;
      LAYER ME1 ;
        RECT 0.62 0.17 0.74 0.53 ;
        RECT 0.63 1.62 0.73 2.04 ;
        RECT 0.11 1.62 0.21 2.04 ;
      LAYER ME2 ;
        RECT 0.11 1.88 0.73 1.98 ;
        RECT 0.63 0.17 0.73 1.98 ;
        RECT 0.11 1.62 0.21 1.98 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.375 1.62 0.465 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.185 -0.22 0.275 0.53 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.11 1.62 0.21 2.04 ;
      RECT 0.225 0.83 0.645 0.93 ;
      RECT 0.275 1.07 0.695 1.17 ;
      RECT 0.63 1.62 0.73 2.04 ;
      RECT 0.62 0.17 0.74 0.53 ;
      RECT 0.375 1.62 0.465 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.185 -0.22 0.275 0.53 ;
    LAYER VI1 ;
      RECT 0.11 1.85 0.21 1.95 ;
      RECT 0.11 1.65 0.21 1.75 ;
      RECT 0.63 1.85 0.73 1.95 ;
      RECT 0.63 1.65 0.73 1.75 ;
      RECT 0.63 0.4 0.73 0.5 ;
      RECT 0.63 0.2 0.73 0.3 ;
    LAYER ME2 ;
      RECT 0.11 1.62 0.21 1.98 ;
      RECT 0.63 0.17 0.73 1.98 ;
      RECT 0.11 1.88 0.73 1.98 ;
  END
END NAND2ALTX1

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN NAND2X1 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.205 1.07 0.625 1.17 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.155 0.83 0.575 0.93 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.37 1.85 0.47 1.95 ;
        RECT 0.37 1.65 0.47 1.75 ;
        RECT 0.56 0.4 0.66 0.5 ;
        RECT 0.56 0.2 0.66 0.3 ;
      LAYER ME1 ;
        RECT 0.55 0.17 0.67 0.53 ;
        RECT 0.36 1.62 0.48 1.98 ;
      LAYER ME2 ;
        RECT 0.37 1.62 0.66 1.72 ;
        RECT 0.56 0.17 0.66 1.72 ;
        RECT 0.37 1.62 0.47 1.98 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 1.62 0.205 2.52 ;
        RECT 0.635 1.62 0.725 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 -0.22 0.205 0.53 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.36 1.62 0.48 1.98 ;
      RECT 0.155 0.83 0.575 0.93 ;
      RECT 0.205 1.07 0.625 1.17 ;
      RECT 0.55 0.17 0.67 0.53 ;
      RECT 0.115 1.62 0.205 2.52 ;
      RECT 0.635 1.62 0.725 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.115 -0.22 0.205 0.53 ;
    LAYER VI1 ;
      RECT 0.37 1.85 0.47 1.95 ;
      RECT 0.37 1.65 0.47 1.75 ;
      RECT 0.56 0.4 0.66 0.5 ;
      RECT 0.56 0.2 0.66 0.3 ;
    LAYER ME2 ;
      RECT 0.56 0.17 0.66 1.72 ;
      RECT 0.37 1.62 0.66 1.72 ;
      RECT 0.37 1.62 0.47 1.98 ;
  END
END NAND2X1

MACRO NAND2X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN NAND2X2 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.23 1.065 0.65 1.165 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.18 0.805 0.6 0.905 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.37 1.79 0.47 1.89 ;
        RECT 0.37 1.59 0.47 1.69 ;
        RECT 0.37 1.39 0.47 1.49 ;
        RECT 0.56 0.55 0.66 0.65 ;
        RECT 0.56 0.35 0.66 0.45 ;
      LAYER ME1 ;
        RECT 0.55 0.32 0.67 0.68 ;
        RECT 0.37 1.36 0.47 1.92 ;
        RECT 0.375 1.32 0.465 1.92 ;
      LAYER ME2 ;
        RECT 0.37 1.36 0.66 1.46 ;
        RECT 0.56 0.32 0.66 1.46 ;
        RECT 0.37 1.36 0.47 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 1.32 0.205 2.52 ;
        RECT 0.635 1.32 0.725 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 -0.22 0.205 0.68 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.375 1.32 0.465 1.92 ;
      RECT 0.37 1.36 0.47 1.92 ;
      RECT 0.18 0.805 0.6 0.905 ;
      RECT 0.23 1.065 0.65 1.165 ;
      RECT 0.55 0.32 0.67 0.68 ;
      RECT 0.115 1.32 0.205 2.52 ;
      RECT 0.635 1.32 0.725 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.115 -0.22 0.205 0.68 ;
    LAYER VI1 ;
      RECT 0.37 1.79 0.47 1.89 ;
      RECT 0.37 1.59 0.47 1.69 ;
      RECT 0.37 1.39 0.47 1.49 ;
      RECT 0.56 0.55 0.66 0.65 ;
      RECT 0.56 0.35 0.66 0.45 ;
    LAYER ME2 ;
      RECT 0.56 0.32 0.66 1.46 ;
      RECT 0.37 1.36 0.66 1.46 ;
      RECT 0.37 1.36 0.47 1.92 ;
  END
END NAND2X2

MACRO NAND2X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN NAND2X4 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.635 1.045 1.055 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.2 0.805 0.62 0.905 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.39 1.79 0.49 1.89 ;
        RECT 0.39 1.59 0.49 1.69 ;
        RECT 0.39 1.39 0.49 1.49 ;
        RECT 0.58 0.55 0.68 0.65 ;
        RECT 0.58 0.35 0.68 0.45 ;
        RECT 0.91 1.79 1.01 1.89 ;
        RECT 0.91 1.59 1.01 1.69 ;
        RECT 0.91 1.39 1.01 1.49 ;
      LAYER ME1 ;
        RECT 0.91 1.36 1.01 1.92 ;
        RECT 0.915 1.32 1.005 1.92 ;
        RECT 0.57 0.32 0.69 0.68 ;
        RECT 0.39 1.36 0.49 1.92 ;
        RECT 0.395 1.32 0.485 1.92 ;
      LAYER ME2 ;
        RECT 0.91 0.58 1.01 1.92 ;
        RECT 0.39 1.585 1.01 1.695 ;
        RECT 0.58 0.58 1.01 0.68 ;
        RECT 0.58 0.32 0.68 0.68 ;
        RECT 0.39 1.36 0.49 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 1.32 0.225 2.52 ;
        RECT 0.655 1.32 0.745 2.52 ;
        RECT 1.175 1.32 1.265 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 -0.22 0.225 0.68 ;
        RECT 1.035 -0.22 1.125 0.68 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.395 1.32 0.485 1.92 ;
      RECT 0.39 1.36 0.49 1.92 ;
      RECT 0.2 0.805 0.62 0.905 ;
      RECT 0.57 0.32 0.69 0.68 ;
      RECT 0.915 1.32 1.005 1.92 ;
      RECT 0.91 1.36 1.01 1.92 ;
      RECT 0.635 1.045 1.055 1.145 ;
      RECT 0.135 1.32 0.225 2.52 ;
      RECT 0.655 1.32 0.745 2.52 ;
      RECT 1.175 1.32 1.265 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.135 -0.22 0.225 0.68 ;
      RECT 1.035 -0.22 1.125 0.68 ;
    LAYER VI1 ;
      RECT 0.39 1.79 0.49 1.89 ;
      RECT 0.39 1.59 0.49 1.69 ;
      RECT 0.39 1.39 0.49 1.49 ;
      RECT 0.58 0.55 0.68 0.65 ;
      RECT 0.58 0.35 0.68 0.45 ;
      RECT 0.91 1.79 1.01 1.89 ;
      RECT 0.91 1.59 1.01 1.69 ;
      RECT 0.91 1.39 1.01 1.49 ;
    LAYER ME2 ;
      RECT 0.58 0.32 0.68 0.68 ;
      RECT 0.58 0.58 1.01 0.68 ;
      RECT 0.39 1.585 1.01 1.695 ;
      RECT 0.39 1.36 0.49 1.92 ;
      RECT 0.91 0.58 1.01 1.92 ;
  END
END NAND2X4

MACRO NOR2ALTX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN NOR2ALTX1 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.18 0.83 0.6 0.93 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.23 1.07 0.65 1.17 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.11 0.4 0.21 0.5 ;
        RECT 0.11 0.2 0.21 0.3 ;
        RECT 0.63 1.85 0.73 1.95 ;
        RECT 0.63 1.65 0.73 1.75 ;
        RECT 0.63 0.4 0.73 0.5 ;
        RECT 0.63 0.2 0.73 0.3 ;
      LAYER ME1 ;
        RECT 0.62 0.17 0.74 0.53 ;
        RECT 0.62 1.62 0.74 1.98 ;
        RECT 0.1 0.17 0.22 0.53 ;
      LAYER ME2 ;
        RECT 0.63 0.17 0.73 1.98 ;
        RECT 0.11 0.43 0.73 0.53 ;
        RECT 0.11 0.17 0.21 0.53 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.185 1.62 0.275 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.375 -0.22 0.465 0.53 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.1 0.17 0.22 0.53 ;
      RECT 0.18 0.83 0.6 0.93 ;
      RECT 0.23 1.07 0.65 1.17 ;
      RECT 0.62 1.62 0.74 1.98 ;
      RECT 0.62 0.17 0.74 0.53 ;
      RECT 0.185 1.62 0.275 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.375 -0.22 0.465 0.53 ;
    LAYER VI1 ;
      RECT 0.11 0.4 0.21 0.5 ;
      RECT 0.11 0.2 0.21 0.3 ;
      RECT 0.63 1.85 0.73 1.95 ;
      RECT 0.63 1.65 0.73 1.75 ;
      RECT 0.63 0.4 0.73 0.5 ;
      RECT 0.63 0.2 0.73 0.3 ;
    LAYER ME2 ;
      RECT 0.11 0.17 0.21 0.53 ;
      RECT 0.11 0.43 0.73 0.53 ;
      RECT 0.63 0.17 0.73 1.98 ;
  END
END NOR2ALTX1

MACRO NOR2X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN NOR2X1 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.18 0.83 0.6 0.93 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.23 1.07 0.65 1.17 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.37 0.4 0.47 0.5 ;
        RECT 0.37 0.2 0.47 0.3 ;
        RECT 0.56 1.85 0.66 1.95 ;
        RECT 0.56 1.65 0.66 1.75 ;
      LAYER ME1 ;
        RECT 0.55 1.62 0.67 1.98 ;
        RECT 0.36 0.17 0.48 0.53 ;
      LAYER ME2 ;
        RECT 0.56 0.43 0.66 1.98 ;
        RECT 0.37 0.43 0.66 0.53 ;
        RECT 0.37 0.17 0.47 0.53 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 1.62 0.205 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 -0.22 0.205 0.53 ;
        RECT 0.635 -0.22 0.725 0.53 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.36 0.17 0.48 0.53 ;
      RECT 0.18 0.83 0.6 0.93 ;
      RECT 0.23 1.07 0.65 1.17 ;
      RECT 0.55 1.62 0.67 1.98 ;
      RECT 0.115 1.62 0.205 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.115 -0.22 0.205 0.53 ;
      RECT 0.635 -0.22 0.725 0.53 ;
    LAYER VI1 ;
      RECT 0.37 0.4 0.47 0.5 ;
      RECT 0.37 0.2 0.47 0.3 ;
      RECT 0.56 1.85 0.66 1.95 ;
      RECT 0.56 1.65 0.66 1.75 ;
    LAYER ME2 ;
      RECT 0.37 0.17 0.47 0.53 ;
      RECT 0.37 0.43 0.66 0.53 ;
      RECT 0.56 0.43 0.66 1.98 ;
  END
END NOR2X1

MACRO NOR2X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN NOR2X2 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.805 0.58 0.905 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.21 1.055 0.63 1.155 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.37 0.55 0.47 0.65 ;
        RECT 0.37 0.35 0.47 0.45 ;
        RECT 0.56 1.79 0.66 1.89 ;
        RECT 0.56 1.59 0.66 1.69 ;
        RECT 0.56 1.39 0.66 1.49 ;
      LAYER ME1 ;
        RECT 0.56 1.36 0.66 1.92 ;
        RECT 0.565 1.32 0.655 1.92 ;
        RECT 0.36 0.32 0.48 0.68 ;
      LAYER ME2 ;
        RECT 0.56 0.58 0.66 1.92 ;
        RECT 0.37 0.58 0.66 0.68 ;
        RECT 0.37 0.32 0.47 0.68 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 1.32 0.205 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 -0.22 0.205 0.68 ;
        RECT 0.635 -0.22 0.725 0.68 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.36 0.32 0.48 0.68 ;
      RECT 0.16 0.805 0.58 0.905 ;
      RECT 0.21 1.055 0.63 1.155 ;
      RECT 0.565 1.32 0.655 1.92 ;
      RECT 0.56 1.36 0.66 1.92 ;
      RECT 0.115 1.32 0.205 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.115 -0.22 0.205 0.68 ;
      RECT 0.635 -0.22 0.725 0.68 ;
    LAYER VI1 ;
      RECT 0.37 0.55 0.47 0.65 ;
      RECT 0.37 0.35 0.47 0.45 ;
      RECT 0.56 1.79 0.66 1.89 ;
      RECT 0.56 1.59 0.66 1.69 ;
      RECT 0.56 1.39 0.66 1.49 ;
    LAYER ME2 ;
      RECT 0.37 0.32 0.47 0.68 ;
      RECT 0.37 0.58 0.66 0.68 ;
      RECT 0.56 0.58 0.66 1.92 ;
  END
END NOR2X2

MACRO NOR2X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN NOR2X4 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.2 0.805 0.62 0.905 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.62 1.045 1.04 1.145 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.39 0.55 0.49 0.65 ;
        RECT 0.39 0.35 0.49 0.45 ;
        RECT 0.58 1.79 0.68 1.89 ;
        RECT 0.58 1.59 0.68 1.69 ;
        RECT 0.58 1.39 0.68 1.49 ;
        RECT 0.91 0.55 1.01 0.65 ;
        RECT 0.91 0.35 1.01 0.45 ;
      LAYER ME1 ;
        RECT 0.9 0.32 1.02 0.68 ;
        RECT 0.58 1.36 0.68 1.92 ;
        RECT 0.585 1.32 0.675 1.92 ;
        RECT 0.38 0.32 0.5 0.68 ;
      LAYER ME2 ;
        RECT 0.39 0.58 1.01 0.68 ;
        RECT 0.91 0.32 1.01 0.68 ;
        RECT 0.58 0.58 0.68 1.92 ;
        RECT 0.39 0.32 0.49 0.68 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 1.32 0.225 2.52 ;
        RECT 1.035 1.32 1.125 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 -0.22 0.225 0.68 ;
        RECT 0.655 -0.22 0.745 0.68 ;
        RECT 1.175 -0.22 1.265 0.68 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.38 0.32 0.5 0.68 ;
      RECT 0.2 0.805 0.62 0.905 ;
      RECT 0.585 1.32 0.675 1.92 ;
      RECT 0.58 1.36 0.68 1.92 ;
      RECT 0.9 0.32 1.02 0.68 ;
      RECT 0.62 1.045 1.04 1.145 ;
      RECT 0.135 1.32 0.225 2.52 ;
      RECT 1.035 1.32 1.125 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.135 -0.22 0.225 0.68 ;
      RECT 0.655 -0.22 0.745 0.68 ;
      RECT 1.175 -0.22 1.265 0.68 ;
    LAYER VI1 ;
      RECT 0.39 0.55 0.49 0.65 ;
      RECT 0.39 0.35 0.49 0.45 ;
      RECT 0.58 1.79 0.68 1.89 ;
      RECT 0.58 1.59 0.68 1.69 ;
      RECT 0.58 1.39 0.68 1.49 ;
      RECT 0.91 0.55 1.01 0.65 ;
      RECT 0.91 0.35 1.01 0.45 ;
    LAYER ME2 ;
      RECT 0.39 0.32 0.49 0.68 ;
      RECT 0.91 0.32 1.01 0.68 ;
      RECT 0.39 0.58 1.01 0.68 ;
      RECT 0.58 0.58 0.68 1.92 ;
  END
END NOR2X4

MACRO OAI211X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI211X1 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.275 0.83 0.695 0.93 ;
    END
  END A2
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.17 1.62 0.26 2.52 ;
        RECT 0.88 1.62 0.97 2.52 ;
        RECT 0 2.3 1.54 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.43 -0.22 0.52 0.53 ;
        RECT -0.14 -0.22 1.54 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.195 1.235 0.615 1.335 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.685 1.06 1.105 1.16 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.135 1.85 1.235 1.95 ;
        RECT 1.135 1.65 1.235 1.75 ;
        RECT 1.135 0.61 1.235 0.71 ;
        RECT 1.135 0.41 1.235 0.51 ;
      LAYER ME1 ;
        RECT 1.125 0.38 1.245 0.74 ;
        RECT 1.125 1.62 1.245 1.98 ;
        RECT 1.14 1.44 1.23 1.98 ;
        RECT 0.62 1.44 1.23 1.53 ;
        RECT 0.62 1.44 0.71 1.92 ;
      LAYER ME2 ;
        RECT 1.135 0.38 1.235 1.98 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.815 0.83 1.235 0.93 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.195 1.235 0.615 1.335 ;
      RECT 0.275 0.83 0.695 0.93 ;
      RECT 0.17 0.38 0.26 0.71 ;
      RECT 0.69 0.38 0.78 0.71 ;
      RECT 0.17 0.62 0.78 0.71 ;
      RECT 0.685 1.06 1.105 1.16 ;
      RECT 0.815 0.83 1.235 0.93 ;
      RECT 0.62 1.44 1.23 1.53 ;
      RECT 1.14 1.44 1.23 1.98 ;
      RECT 0.62 1.44 0.71 1.92 ;
      RECT 1.125 1.62 1.245 1.98 ;
      RECT 1.125 0.38 1.245 0.74 ;
      RECT 0.17 1.62 0.26 2.52 ;
      RECT 0.88 1.62 0.97 2.52 ;
      RECT 0 2.3 1.54 2.52 ;
      RECT -0.14 -0.22 1.54 0 ;
      RECT 0.43 -0.22 0.52 0.53 ;
    LAYER VI1 ;
      RECT 1.135 1.85 1.235 1.95 ;
      RECT 1.135 1.65 1.235 1.75 ;
      RECT 1.135 0.61 1.235 0.71 ;
      RECT 1.135 0.41 1.235 0.51 ;
    LAYER ME2 ;
      RECT 1.135 0.38 1.235 1.98 ;
  END
END OAI211X1

MACRO OAI211X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI211X2 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.225 1.07 0.645 1.17 ;
    END
  END A2
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.17 1.32 0.26 2.52 ;
        RECT 0.88 1.32 0.97 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.43 -0.22 0.52 0.68 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.17 0.83 0.59 0.93 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.755 0.83 1.175 0.93 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.61 2.03 0.71 2.13 ;
        RECT 1.1 2.03 1.2 2.13 ;
        RECT 1.135 1.79 1.235 1.89 ;
        RECT 1.135 1.59 1.235 1.69 ;
        RECT 1.135 1.39 1.235 1.49 ;
        RECT 1.135 0.55 1.235 0.65 ;
        RECT 1.135 0.35 1.235 0.45 ;
      LAYER ME1 ;
        RECT 1.125 0.32 1.245 0.68 ;
        RECT 1.135 1.36 1.235 1.92 ;
        RECT 1.07 2.03 1.23 2.13 ;
        RECT 1.14 1.32 1.23 2.13 ;
        RECT 0.58 2.03 0.74 2.13 ;
        RECT 0.62 1.32 0.71 2.13 ;
      LAYER ME2 ;
        RECT 1.135 0.32 1.235 1.92 ;
        RECT 0.58 2.03 1.23 2.13 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.765 1.07 1.185 1.17 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.17 0.19 0.33 0.29 ;
      RECT 0.17 0.19 0.26 0.68 ;
      RECT 0.17 0.83 0.59 0.93 ;
      RECT 0.225 1.07 0.645 1.17 ;
      RECT 0.62 1.32 0.71 2.13 ;
      RECT 0.58 2.03 0.74 2.13 ;
      RECT 0.66 0.19 0.82 0.29 ;
      RECT 0.69 0.19 0.78 0.68 ;
      RECT 0.755 0.83 1.175 0.93 ;
      RECT 0.765 1.07 1.185 1.17 ;
      RECT 1.135 1.36 1.235 1.92 ;
      RECT 1.14 1.32 1.23 2.13 ;
      RECT 1.07 2.03 1.23 2.13 ;
      RECT 1.125 0.32 1.245 0.68 ;
      RECT 0.17 1.32 0.26 2.52 ;
      RECT 0.88 1.32 0.97 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.43 -0.22 0.52 0.68 ;
    LAYER VI1 ;
      RECT 0.2 0.19 0.3 0.29 ;
      RECT 0.61 2.03 0.71 2.13 ;
      RECT 0.69 0.19 0.79 0.29 ;
      RECT 1.1 2.03 1.2 2.13 ;
      RECT 1.135 1.79 1.235 1.89 ;
      RECT 1.135 1.59 1.235 1.69 ;
      RECT 1.135 1.39 1.235 1.49 ;
      RECT 1.135 0.55 1.235 0.65 ;
      RECT 1.135 0.35 1.235 0.45 ;
    LAYER ME2 ;
      RECT 0.17 0.19 0.82 0.29 ;
      RECT 0.58 2.03 1.23 2.13 ;
      RECT 1.135 0.32 1.235 1.92 ;
  END
END OAI211X2

MACRO OAI211X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI211X4 0 -0.11 ;
  SIZE 2.52 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.235 1.075 0.655 1.175 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.68 1.79 0.78 1.89 ;
        RECT 0.68 1.59 0.78 1.69 ;
        RECT 0.68 1.39 0.78 1.49 ;
        RECT 1.39 1.79 1.49 1.89 ;
        RECT 1.39 1.59 1.49 1.69 ;
        RECT 1.39 1.39 1.49 1.49 ;
        RECT 1.46 0.55 1.56 0.65 ;
        RECT 1.46 0.35 1.56 0.45 ;
        RECT 1.91 1.79 2.01 1.89 ;
        RECT 1.91 1.59 2.01 1.69 ;
        RECT 1.91 1.39 2.01 1.49 ;
      LAYER ME1 ;
        RECT 1.91 1.36 2.01 1.92 ;
        RECT 1.915 1.32 2.005 1.92 ;
        RECT 1.45 0.32 1.57 0.68 ;
        RECT 1.39 1.36 1.49 1.92 ;
        RECT 1.395 1.32 1.485 1.92 ;
        RECT 0.68 1.36 0.78 1.92 ;
        RECT 0.685 1.32 0.775 1.92 ;
      LAYER ME2 ;
        RECT 1.91 1.36 2.01 1.92 ;
        RECT 0.68 1.59 2.01 1.69 ;
        RECT 1.39 1.36 1.56 1.92 ;
        RECT 1.46 0.32 1.56 1.92 ;
        RECT 0.68 1.36 0.78 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.235 1.32 0.325 2.52 ;
        RECT 1.135 1.32 1.225 2.52 ;
        RECT 1.655 1.32 1.745 2.52 ;
        RECT 2.175 1.32 2.265 2.52 ;
        RECT 0 2.3 2.52 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.235 -0.22 0.325 0.68 ;
        RECT 0.755 -0.22 0.845 0.68 ;
        RECT 2.175 -0.22 2.265 0.68 ;
        RECT 0 -0.22 2.52 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.82 0.825 2.15 0.925 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.055 1.075 1.475 1.175 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.735 1.075 2.155 1.175 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.48 0.32 0.6 0.68 ;
      RECT 0.235 1.075 0.655 1.175 ;
      RECT 0.685 1.32 0.775 1.92 ;
      RECT 0.68 1.36 0.78 1.92 ;
      RECT 1.055 1.075 1.475 1.175 ;
      RECT 1.395 1.32 1.485 1.92 ;
      RECT 1.39 1.36 1.49 1.92 ;
      RECT 1.45 0.32 1.57 0.68 ;
      RECT 1.015 0.14 2.005 0.23 ;
      RECT 1.015 0.14 1.105 0.68 ;
      RECT 1.01 0.32 1.11 0.68 ;
      RECT 1.915 0.14 2.005 0.68 ;
      RECT 1.915 1.32 2.005 1.92 ;
      RECT 1.91 1.36 2.01 1.92 ;
      RECT 0.82 0.825 2.15 0.925 ;
      RECT 1.735 1.075 2.155 1.175 ;
      RECT 0.235 1.32 0.325 2.52 ;
      RECT 1.135 1.32 1.225 2.52 ;
      RECT 1.655 1.32 1.745 2.52 ;
      RECT 2.175 1.32 2.265 2.52 ;
      RECT 0 2.3 2.52 2.52 ;
      RECT 0 -0.22 2.52 0 ;
      RECT 0.235 -0.22 0.325 0.68 ;
      RECT 0.755 -0.22 0.845 0.68 ;
      RECT 2.175 -0.22 2.265 0.68 ;
    LAYER VI1 ;
      RECT 0.49 0.55 0.59 0.65 ;
      RECT 0.49 0.35 0.59 0.45 ;
      RECT 0.68 1.79 0.78 1.89 ;
      RECT 0.68 1.59 0.78 1.69 ;
      RECT 0.68 1.39 0.78 1.49 ;
      RECT 1.01 0.55 1.11 0.65 ;
      RECT 1.01 0.35 1.11 0.45 ;
      RECT 1.39 1.79 1.49 1.89 ;
      RECT 1.39 1.59 1.49 1.69 ;
      RECT 1.39 1.39 1.49 1.49 ;
      RECT 1.46 0.55 1.56 0.65 ;
      RECT 1.46 0.35 1.56 0.45 ;
      RECT 1.91 1.79 2.01 1.89 ;
      RECT 1.91 1.59 2.01 1.69 ;
      RECT 1.91 1.39 2.01 1.49 ;
    LAYER ME2 ;
      RECT 0.49 0.51 1.11 0.61 ;
      RECT 0.49 0.32 0.59 0.68 ;
      RECT 1.01 0.32 1.11 0.68 ;
      RECT 0.68 1.59 2.01 1.69 ;
      RECT 0.68 1.36 0.78 1.92 ;
      RECT 1.46 0.32 1.56 1.92 ;
      RECT 1.39 1.36 1.56 1.92 ;
      RECT 1.91 1.36 2.01 1.92 ;
  END
END OAI211X4

MACRO OAI21X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI21X1 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.45 0.825 0.87 0.925 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.83 1.85 0.93 1.95 ;
        RECT 0.83 1.65 0.93 1.75 ;
        RECT 0.9 0.4 1 0.5 ;
        RECT 0.9 0.2 1 0.3 ;
      LAYER ME1 ;
        RECT 0.89 0.17 1.01 0.53 ;
        RECT 0.82 1.62 0.94 1.98 ;
        RECT 0.835 1.44 0.925 1.98 ;
        RECT 0.125 1.44 0.925 1.53 ;
        RECT 0.125 1.44 0.215 1.92 ;
      LAYER ME2 ;
        RECT 0.83 0.17 1 0.53 ;
        RECT 0.83 0.17 0.93 1.98 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.575 1.62 0.665 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.385 -0.22 0.475 0.53 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.16 1.025 0.58 1.125 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.51 1.225 0.93 1.325 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.16 1.025 0.58 1.125 ;
      RECT 0.125 0.38 0.215 0.71 ;
      RECT 0.645 0.38 0.735 0.71 ;
      RECT 0.125 0.62 0.735 0.71 ;
      RECT 0.45 0.825 0.87 0.925 ;
      RECT 0.51 1.225 0.93 1.325 ;
      RECT 0.125 1.44 0.925 1.53 ;
      RECT 0.835 1.44 0.925 1.98 ;
      RECT 0.125 1.44 0.215 1.92 ;
      RECT 0.82 1.62 0.94 1.98 ;
      RECT 0.89 0.17 1.01 0.53 ;
      RECT 0.575 1.62 0.665 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.385 -0.22 0.475 0.53 ;
    LAYER VI1 ;
      RECT 0.83 1.85 0.93 1.95 ;
      RECT 0.83 1.65 0.93 1.75 ;
      RECT 0.9 0.4 1 0.5 ;
      RECT 0.9 0.2 1 0.3 ;
    LAYER ME2 ;
      RECT 0.83 0.17 1 0.53 ;
      RECT 0.83 0.17 0.93 1.98 ;
  END
END OAI21X1

MACRO OAI21X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI21X2 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.45 0.795 0.87 0.895 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.155 2.03 0.255 2.13 ;
        RECT 0.83 1.79 0.93 1.89 ;
        RECT 0.83 1.59 0.93 1.69 ;
        RECT 0.83 1.39 0.93 1.49 ;
        RECT 0.9 0.48 1 0.58 ;
      LAYER ME1 ;
        RECT 0.88 0.38 1.02 0.68 ;
        RECT 0.83 1.36 0.93 1.92 ;
        RECT 0.835 1.32 0.925 1.92 ;
        RECT 0.125 2.03 0.285 2.13 ;
        RECT 0.125 1.32 0.215 2.13 ;
      LAYER ME2 ;
        RECT 0.83 0.38 1 0.68 ;
        RECT 0.125 2.03 0.93 2.13 ;
        RECT 0.83 0.38 0.93 2.13 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.575 1.32 0.665 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.385 -0.22 0.475 0.68 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.125 0.96 0.375 1.13 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.575 1.105 0.995 1.205 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.125 1.32 0.215 2.13 ;
      RECT 0.125 2.03 0.285 2.13 ;
      RECT 0.125 0.19 0.285 0.29 ;
      RECT 0.125 0.19 0.215 0.68 ;
      RECT 0.125 0.96 0.375 1.13 ;
      RECT 0.615 0.19 0.775 0.29 ;
      RECT 0.645 0.19 0.735 0.68 ;
      RECT 0.45 0.795 0.87 0.895 ;
      RECT 0.835 1.32 0.925 1.92 ;
      RECT 0.83 1.36 0.93 1.92 ;
      RECT 0.575 1.105 0.995 1.205 ;
      RECT 0.88 0.38 1.02 0.68 ;
      RECT 0.575 1.32 0.665 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.385 -0.22 0.475 0.68 ;
    LAYER VI1 ;
      RECT 0.155 2.03 0.255 2.13 ;
      RECT 0.155 0.19 0.255 0.29 ;
      RECT 0.645 0.19 0.745 0.29 ;
      RECT 0.83 1.79 0.93 1.89 ;
      RECT 0.83 1.59 0.93 1.69 ;
      RECT 0.83 1.39 0.93 1.49 ;
      RECT 0.9 0.48 1 0.58 ;
    LAYER ME2 ;
      RECT 0.125 0.19 0.775 0.29 ;
      RECT 0.83 0.38 1 0.68 ;
      RECT 0.83 0.38 0.93 2.13 ;
      RECT 0.125 2.03 0.93 2.13 ;
  END
END OAI21X2

MACRO OAI21X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI21X4 0 -0.11 ;
  SIZE 1.96 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.49 1.105 0.91 1.205 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.67 1.79 0.77 1.89 ;
        RECT 0.67 1.59 0.77 1.69 ;
        RECT 0.67 1.39 0.77 1.49 ;
        RECT 1.19 0.55 1.29 0.65 ;
        RECT 1.19 0.35 1.29 0.45 ;
        RECT 1.38 1.79 1.48 1.89 ;
        RECT 1.38 1.59 1.48 1.69 ;
        RECT 1.38 1.39 1.48 1.49 ;
      LAYER ME1 ;
        RECT 1.38 1.36 1.48 1.92 ;
        RECT 1.385 1.32 1.475 1.92 ;
        RECT 1.18 0.32 1.3 0.68 ;
        RECT 0.67 1.36 0.77 1.92 ;
        RECT 0.675 1.32 0.765 1.92 ;
      LAYER ME2 ;
        RECT 1.38 0.58 1.48 1.92 ;
        RECT 0.67 1.65 1.48 1.75 ;
        RECT 1.19 0.58 1.48 0.68 ;
        RECT 1.19 0.32 1.29 0.68 ;
        RECT 0.67 1.36 0.77 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.225 1.32 0.315 2.52 ;
        RECT 1.125 1.32 1.215 2.52 ;
        RECT 1.645 1.32 1.735 2.52 ;
        RECT 0 2.3 1.96 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.155 -0.22 0.245 0.68 ;
        RECT 0.675 -0.22 0.765 0.68 ;
        RECT 1.715 -0.22 1.805 0.68 ;
        RECT 0 -0.22 1.96 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.23 0.825 0.65 0.925 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.2 1.105 1.62 1.205 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.4 0.32 0.52 0.68 ;
      RECT 0.23 0.825 0.65 0.925 ;
      RECT 0.675 1.32 0.765 1.92 ;
      RECT 0.67 1.36 0.77 1.92 ;
      RECT 0.49 1.105 0.91 1.205 ;
      RECT 1.18 0.32 1.3 0.68 ;
      RECT 1.385 1.32 1.475 1.92 ;
      RECT 1.38 1.36 1.48 1.92 ;
      RECT 0.935 0.12 1.545 0.21 ;
      RECT 0.935 0.12 1.025 0.68 ;
      RECT 0.92 0.32 1.04 0.68 ;
      RECT 1.455 0.12 1.545 0.68 ;
      RECT 1.2 1.105 1.62 1.205 ;
      RECT 0.225 1.32 0.315 2.52 ;
      RECT 1.125 1.32 1.215 2.52 ;
      RECT 1.645 1.32 1.735 2.52 ;
      RECT 0 2.3 1.96 2.52 ;
      RECT 0 -0.22 1.96 0 ;
      RECT 0.155 -0.22 0.245 0.68 ;
      RECT 0.675 -0.22 0.765 0.68 ;
      RECT 1.715 -0.22 1.805 0.68 ;
    LAYER VI1 ;
      RECT 0.41 0.55 0.51 0.65 ;
      RECT 0.41 0.35 0.51 0.45 ;
      RECT 0.67 1.79 0.77 1.89 ;
      RECT 0.67 1.59 0.77 1.69 ;
      RECT 0.67 1.39 0.77 1.49 ;
      RECT 0.93 0.55 1.03 0.65 ;
      RECT 0.93 0.35 1.03 0.45 ;
      RECT 1.19 0.55 1.29 0.65 ;
      RECT 1.19 0.35 1.29 0.45 ;
      RECT 1.38 1.79 1.48 1.89 ;
      RECT 1.38 1.59 1.48 1.69 ;
      RECT 1.38 1.39 1.48 1.49 ;
    LAYER ME2 ;
      RECT 0.41 0.45 1.03 0.55 ;
      RECT 0.41 0.32 0.51 0.68 ;
      RECT 0.93 0.32 1.03 0.68 ;
      RECT 1.19 0.32 1.29 0.68 ;
      RECT 1.19 0.58 1.48 0.68 ;
      RECT 0.67 1.65 1.48 1.75 ;
      RECT 0.67 1.36 0.77 1.92 ;
      RECT 1.38 0.58 1.48 1.92 ;
  END
END OAI21X4

MACRO OAI22X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI22X1 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.19 1.125 0.61 1.225 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.755 1.125 1.175 1.225 ;
    END
  END B2
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 1.62 0.225 2.52 ;
        RECT 1.035 1.62 1.125 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.395 -0.22 0.485 0.53 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.19 0.84 0.61 0.94 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.72 0.84 1.14 0.94 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.58 1.85 0.68 1.95 ;
        RECT 0.58 1.65 0.68 1.75 ;
        RECT 0.91 0.41 1.01 0.51 ;
      LAYER ME1 ;
        RECT 0.9 0.38 1.02 0.74 ;
        RECT 0.57 1.62 0.69 1.98 ;
      LAYER ME2 ;
        RECT 0.91 0.38 1.01 0.54 ;
        RECT 0.58 0.41 1.01 0.51 ;
        RECT 0.58 0.41 0.68 1.98 ;
    END
  END Y
  OBS
    LAYER ME1 ;
      RECT 0.19 1.125 0.61 1.225 ;
      RECT 0.19 0.84 0.61 0.94 ;
      RECT 0.57 1.62 0.69 1.98 ;
      RECT 0.9 0.38 1.02 0.74 ;
      RECT 0.72 0.84 1.14 0.94 ;
      RECT 0.755 1.125 1.175 1.225 ;
      RECT 0.655 0.2 1.265 0.29 ;
      RECT 1.175 0.2 1.265 0.53 ;
      RECT 0.135 0.38 0.225 0.71 ;
      RECT 0.655 0.2 0.745 0.71 ;
      RECT 0.135 0.62 0.745 0.71 ;
      RECT 0.135 1.62 0.225 2.52 ;
      RECT 1.035 1.62 1.125 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.395 -0.22 0.485 0.53 ;
    LAYER VI1 ;
      RECT 0.58 1.85 0.68 1.95 ;
      RECT 0.58 1.65 0.68 1.75 ;
      RECT 0.91 0.41 1.01 0.51 ;
    LAYER ME2 ;
      RECT 0.58 0.41 1.01 0.51 ;
      RECT 0.91 0.38 1.01 0.54 ;
      RECT 0.58 0.41 0.68 1.98 ;
  END
END OAI22X1

MACRO OAI22X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI22X2 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.19 1.07 0.61 1.17 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.815 1.07 1.235 1.17 ;
    END
  END B2
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 1.32 0.225 2.52 ;
        RECT 1.035 1.32 1.125 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.395 -0.22 0.485 0.68 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.135 0.83 0.555 0.93 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.58 1.79 0.68 1.89 ;
        RECT 0.58 1.59 0.68 1.69 ;
        RECT 0.58 1.39 0.68 1.49 ;
        RECT 0.91 0.55 1.01 0.65 ;
        RECT 0.91 0.35 1.01 0.45 ;
      LAYER ME1 ;
        RECT 0.9 0.32 1.02 0.68 ;
        RECT 0.58 1.36 0.68 1.92 ;
        RECT 0.585 1.32 0.675 1.92 ;
      LAYER ME2 ;
        RECT 0.58 0.58 1.01 0.68 ;
        RECT 0.91 0.32 1.01 0.68 ;
        RECT 0.58 0.58 0.68 1.92 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.72 0.83 1.14 0.93 ;
    END
  END B1
  OBS
    LAYER ME1 ;
      RECT 0.135 0.13 0.295 0.23 ;
      RECT 0.135 0.13 0.225 0.68 ;
      RECT 0.135 0.83 0.555 0.93 ;
      RECT 0.19 1.07 0.61 1.17 ;
      RECT 0.585 1.32 0.675 1.92 ;
      RECT 0.58 1.36 0.68 1.92 ;
      RECT 0.9 0.32 1.02 0.68 ;
      RECT 0.72 0.83 1.14 0.93 ;
      RECT 0.815 1.07 1.235 1.17 ;
      RECT 0.62 0.135 1.265 0.225 ;
      RECT 0.62 0.13 0.78 0.23 ;
      RECT 0.655 0.13 0.745 0.68 ;
      RECT 1.175 0.135 1.265 0.68 ;
      RECT 0.135 1.32 0.225 2.52 ;
      RECT 1.035 1.32 1.125 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.395 -0.22 0.485 0.68 ;
    LAYER VI1 ;
      RECT 0.165 0.13 0.265 0.23 ;
      RECT 0.58 1.79 0.68 1.89 ;
      RECT 0.58 1.59 0.68 1.69 ;
      RECT 0.58 1.39 0.68 1.49 ;
      RECT 0.65 0.13 0.75 0.23 ;
      RECT 0.91 0.55 1.01 0.65 ;
      RECT 0.91 0.35 1.01 0.45 ;
    LAYER ME2 ;
      RECT 0.135 0.13 0.78 0.23 ;
      RECT 0.91 0.32 1.01 0.68 ;
      RECT 0.58 0.58 1.01 0.68 ;
      RECT 0.58 0.58 0.68 1.92 ;
  END
END OAI22X2

MACRO OAI22X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OAI22X4 0 -0.11 ;
  SIZE 2.52 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.62 1.75 0.72 1.85 ;
        RECT 0.62 1.55 0.72 1.65 ;
        RECT 0.62 1.35 0.72 1.45 ;
        RECT 1.47 0.755 1.57 0.855 ;
        RECT 1.52 1.75 1.62 1.85 ;
        RECT 1.52 1.55 1.62 1.65 ;
        RECT 1.52 1.35 1.62 1.45 ;
      LAYER ME2 ;
        RECT 1.47 1.32 1.62 1.88 ;
        RECT 1.47 0.725 1.57 1.88 ;
        RECT 0.62 1.745 1.62 1.855 ;
        RECT 0.62 1.32 0.72 1.88 ;
      LAYER ME1 ;
        RECT 1.995 0.14 2.085 0.68 ;
        RECT 1.475 0.14 2.085 0.23 ;
        RECT 1.47 0.68 1.57 0.885 ;
        RECT 1.475 0.14 1.565 0.885 ;
        RECT 1.52 1.32 1.62 1.88 ;
        RECT 1.525 1.32 1.615 1.92 ;
        RECT 0.62 1.32 0.72 1.88 ;
        RECT 0.625 1.32 0.715 1.92 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.74 0.83 2.16 0.93 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.155 1.07 0.575 1.185 ;
    END
  END A1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.175 1.32 0.265 2.52 ;
        RECT 1.075 1.32 1.165 2.52 ;
        RECT 1.975 1.32 2.065 2.52 ;
        RECT 0 2.3 2.52 2.52 ;
    END
  END vdd!
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.45 1.07 1.87 1.17 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.62 0.83 1.04 0.93 ;
    END
  END A2
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.435 -0.22 0.525 0.68 ;
        RECT 0.955 -0.22 1.045 0.68 ;
        RECT 0 -0.22 2.52 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.16 0.32 0.28 0.68 ;
      RECT 0.155 1.07 0.575 1.185 ;
      RECT 0.62 1.32 0.72 1.88 ;
      RECT 0.625 1.32 0.715 1.92 ;
      RECT 0.68 0.32 0.8 0.68 ;
      RECT 0.62 0.83 1.04 0.93 ;
      RECT 1.2 0.32 1.32 0.68 ;
      RECT 1.52 1.32 1.62 1.88 ;
      RECT 1.525 1.32 1.615 1.92 ;
      RECT 1.72 0.32 1.84 0.68 ;
      RECT 1.45 1.07 1.87 1.17 ;
      RECT 1.475 0.14 2.085 0.23 ;
      RECT 1.475 0.14 1.565 0.885 ;
      RECT 1.995 0.14 2.085 0.68 ;
      RECT 1.47 0.68 1.57 0.885 ;
      RECT 1.74 0.83 2.16 0.93 ;
      RECT 2.24 0.32 2.36 0.68 ;
      RECT 0.175 1.32 0.265 2.52 ;
      RECT 1.075 1.32 1.165 2.52 ;
      RECT 1.975 1.32 2.065 2.52 ;
      RECT 0 2.3 2.52 2.52 ;
      RECT 0 -0.22 2.52 0 ;
      RECT 0.435 -0.22 0.525 0.68 ;
      RECT 0.955 -0.22 1.045 0.68 ;
    LAYER VI1 ;
      RECT 0.17 0.55 0.27 0.65 ;
      RECT 0.17 0.35 0.27 0.45 ;
      RECT 0.62 1.75 0.72 1.85 ;
      RECT 0.62 1.55 0.72 1.65 ;
      RECT 0.62 1.35 0.72 1.45 ;
      RECT 0.69 0.55 0.79 0.65 ;
      RECT 0.69 0.35 0.79 0.45 ;
      RECT 1.21 0.55 1.31 0.65 ;
      RECT 1.21 0.35 1.31 0.45 ;
      RECT 1.47 0.755 1.57 0.855 ;
      RECT 1.52 1.75 1.62 1.85 ;
      RECT 1.52 1.55 1.62 1.65 ;
      RECT 1.52 1.35 1.62 1.45 ;
      RECT 1.73 0.55 1.83 0.65 ;
      RECT 1.73 0.35 1.83 0.45 ;
      RECT 2.25 0.55 2.35 0.65 ;
      RECT 2.25 0.35 2.35 0.45 ;
    LAYER ME2 ;
      RECT 1.47 0.725 1.57 1.88 ;
      RECT 0.62 1.745 1.62 1.855 ;
      RECT 0.62 1.32 0.72 1.88 ;
      RECT 1.47 1.32 1.62 1.88 ;
      RECT 0.17 0.445 2.35 0.555 ;
      RECT 0.17 0.32 0.27 0.68 ;
      RECT 0.69 0.32 0.79 0.68 ;
      RECT 1.21 0.32 1.31 0.68 ;
      RECT 1.73 0.32 1.83 0.68 ;
      RECT 2.25 0.32 2.35 0.68 ;
  END
END OAI22X4

MACRO OR2X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OR2X1 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.25 1.085 0.67 1.185 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.2 1.325 0.62 1.425 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.9 1.85 1 1.95 ;
        RECT 0.9 1.65 1 1.75 ;
        RECT 0.9 0.4 1 0.5 ;
        RECT 0.9 0.2 1 0.3 ;
      LAYER ME1 ;
        RECT 0.89 0.17 1.01 0.53 ;
        RECT 0.89 1.62 1.01 1.98 ;
      LAYER ME2 ;
        RECT 0.9 0.17 1 1.98 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.645 1.62 0.735 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.125 -0.22 0.215 0.53 ;
        RECT 0.645 -0.22 0.735 0.53 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.18 1.62 0.3 1.98 ;
      RECT 0.37 0.17 0.49 0.53 ;
      RECT 0.2 1.325 0.62 1.425 ;
      RECT 0.25 1.085 0.67 1.185 ;
      RECT 0.16 0.78 0.88 0.87 ;
      RECT 0.16 0.775 0.32 0.875 ;
      RECT 0.89 1.62 1.01 1.98 ;
      RECT 0.89 0.17 1.01 0.53 ;
      RECT 0.645 1.62 0.735 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.125 -0.22 0.215 0.53 ;
      RECT 0.645 -0.22 0.735 0.53 ;
    LAYER VI1 ;
      RECT 0.19 1.85 0.29 1.95 ;
      RECT 0.19 1.65 0.29 1.75 ;
      RECT 0.19 0.775 0.29 0.875 ;
      RECT 0.38 0.4 0.48 0.5 ;
      RECT 0.38 0.2 0.48 0.3 ;
      RECT 0.9 1.85 1 1.95 ;
      RECT 0.9 1.65 1 1.75 ;
      RECT 0.9 0.4 1 0.5 ;
      RECT 0.9 0.2 1 0.3 ;
    LAYER ME2 ;
      RECT 0.38 0.17 0.48 0.53 ;
      RECT 0.19 0.43 0.48 0.53 ;
      RECT 0.19 0.43 0.29 1.98 ;
      RECT 0.9 0.17 1 1.98 ;
  END
END OR2X1

MACRO OR2X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OR2X2 0 -0.11 ;
  SIZE 1.12 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.5 1.075 0.92 1.175 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.13 1.03 0.41 1.18 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.9 1.79 1 1.89 ;
        RECT 0.9 1.59 1 1.69 ;
        RECT 0.9 1.39 1 1.49 ;
        RECT 0.9 0.55 1 0.65 ;
        RECT 0.9 0.35 1 0.45 ;
      LAYER ME1 ;
        RECT 0.89 0.32 1.01 0.68 ;
        RECT 0.9 1.36 1 1.92 ;
        RECT 0.905 1.32 0.995 1.92 ;
      LAYER ME2 ;
        RECT 0.9 0.32 1 1.92 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.645 1.32 0.735 2.52 ;
        RECT 0 2.3 1.12 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.125 -0.22 0.215 0.68 ;
        RECT 0.645 -0.22 0.735 0.68 ;
        RECT 0 -0.22 1.12 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.195 1.32 0.285 1.92 ;
      RECT 0.19 1.36 0.29 1.92 ;
      RECT 0.13 1.03 0.41 1.18 ;
      RECT 0.37 0.32 0.49 0.68 ;
      RECT 0.35 0.785 0.88 0.875 ;
      RECT 0.35 0.78 0.51 0.88 ;
      RECT 0.5 1.075 0.92 1.175 ;
      RECT 0.905 1.32 0.995 1.92 ;
      RECT 0.9 1.36 1 1.92 ;
      RECT 0.89 0.32 1.01 0.68 ;
      RECT 0.645 1.32 0.735 2.52 ;
      RECT 0 2.3 1.12 2.52 ;
      RECT 0 -0.22 1.12 0 ;
      RECT 0.125 -0.22 0.215 0.68 ;
      RECT 0.645 -0.22 0.735 0.68 ;
    LAYER VI1 ;
      RECT 0.19 1.79 0.29 1.89 ;
      RECT 0.19 1.59 0.29 1.69 ;
      RECT 0.19 1.39 0.29 1.49 ;
      RECT 0.38 0.78 0.48 0.88 ;
      RECT 0.38 0.55 0.48 0.65 ;
      RECT 0.38 0.35 0.48 0.45 ;
      RECT 0.9 1.79 1 1.89 ;
      RECT 0.9 1.59 1 1.69 ;
      RECT 0.9 1.39 1 1.49 ;
      RECT 0.9 0.55 1 0.65 ;
      RECT 0.9 0.35 1 0.45 ;
    LAYER ME2 ;
      RECT 0.38 0.32 0.48 1.46 ;
      RECT 0.19 1.36 0.48 1.46 ;
      RECT 0.19 1.36 0.29 1.92 ;
      RECT 0.9 0.32 1 1.92 ;
  END
END OR2X2

MACRO OR2X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN OR2X4 0 -0.11 ;
  SIZE 1.4 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.91 1.79 1.01 1.89 ;
        RECT 0.91 1.59 1.01 1.69 ;
        RECT 0.91 1.39 1.01 1.49 ;
        RECT 0.91 0.55 1.01 0.65 ;
        RECT 0.91 0.35 1.01 0.45 ;
      LAYER ME2 ;
        RECT 0.91 0.32 1.01 1.92 ;
      LAYER ME1 ;
        RECT 0.9 0.32 1.02 0.68 ;
        RECT 0.91 1.36 1.01 1.92 ;
        RECT 0.915 1.32 1.005 1.92 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.135 -0.22 0.225 0.68 ;
        RECT 0.655 -0.22 0.745 0.68 ;
        RECT 1.175 -0.22 1.265 0.68 ;
        RECT 0 -0.22 1.4 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.655 1.32 0.745 2.52 ;
        RECT 1.175 1.32 1.265 2.52 ;
        RECT 0 2.3 1.4 2.52 ;
    END
  END vdd!
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.005 0.42 1.155 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.51 1.055 0.93 1.155 ;
    END
  END A
  OBS
    LAYER ME1 ;
      RECT 0.205 1.32 0.295 1.92 ;
      RECT 0.2 1.36 0.3 1.92 ;
      RECT 0.14 1.005 0.42 1.155 ;
      RECT 0.38 0.32 0.5 0.68 ;
      RECT 0.51 1.055 0.93 1.155 ;
      RECT 0.915 1.32 1.005 1.92 ;
      RECT 0.91 1.36 1.01 1.92 ;
      RECT 0.9 0.32 1.02 0.68 ;
      RECT 0.36 0.8 1.12 0.89 ;
      RECT 0.36 0.795 0.52 0.895 ;
      RECT 0.655 1.32 0.745 2.52 ;
      RECT 1.175 1.32 1.265 2.52 ;
      RECT 0 2.3 1.4 2.52 ;
      RECT 0 -0.22 1.4 0 ;
      RECT 0.135 -0.22 0.225 0.68 ;
      RECT 0.655 -0.22 0.745 0.68 ;
      RECT 1.175 -0.22 1.265 0.68 ;
    LAYER VI1 ;
      RECT 0.2 1.79 0.3 1.89 ;
      RECT 0.2 1.59 0.3 1.69 ;
      RECT 0.2 1.39 0.3 1.49 ;
      RECT 0.39 0.795 0.49 0.895 ;
      RECT 0.39 0.55 0.49 0.65 ;
      RECT 0.39 0.35 0.49 0.45 ;
      RECT 0.91 1.79 1.01 1.89 ;
      RECT 0.91 1.59 1.01 1.69 ;
      RECT 0.91 1.39 1.01 1.49 ;
      RECT 0.91 0.55 1.01 0.65 ;
      RECT 0.91 0.35 1.01 0.45 ;
    LAYER ME2 ;
      RECT 0.39 0.32 0.49 1.46 ;
      RECT 0.2 1.36 0.49 1.46 ;
      RECT 0.2 1.36 0.3 1.92 ;
      RECT 0.91 0.32 1.01 1.92 ;
  END
END OR2X4

MACRO QDFFCNSX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDFFCNSX1 0 -0.11 ;
  SIZE 4.2 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 1.91 1.15 3.21 1.25 ;
        RECT 2.88 1.135 3.21 1.265 ;
    END
  END CLK
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.405 1.62 0.495 2.52 ;
        RECT 1.305 1.62 1.395 2.52 ;
        RECT 2.055 1.62 2.145 2.52 ;
        RECT 2.545 1.62 2.635 2.52 ;
        RECT 3.445 1.62 3.535 2.52 ;
        RECT 3.965 1.62 4.055 2.52 ;
        RECT 0 2.3 4.2 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.405 -0.22 0.495 0.53 ;
        RECT 1.305 -0.22 1.395 0.53 ;
        RECT 2.055 -0.22 2.145 0.53 ;
        RECT 2.545 -0.22 2.635 0.53 ;
        RECT 3.445 -0.22 3.535 0.53 ;
        RECT 0 -0.22 4.2 0 ;
    END
  END gnd!
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 3.57 1.18 3.99 1.28 ;
    END
  END SETB
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.335 1.195 0.755 1.295 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 3.7 1.72 3.8 1.82 ;
        RECT 3.89 0.63 3.99 0.73 ;
        RECT 3.89 0.4 3.99 0.5 ;
      LAYER ME1 ;
        RECT 3.86 0.23 4.02 0.53 ;
        RECT 3.32 0.63 4.02 0.73 ;
        RECT 3.67 1.62 3.83 1.92 ;
      LAYER ME2 ;
        RECT 3.7 1.62 3.99 1.72 ;
        RECT 3.89 0.37 3.99 1.72 ;
        RECT 3.7 1.62 3.8 1.92 ;
    END
  END Q
  OBS
    LAYER ME1 ;
      RECT 0.11 1.62 0.27 1.92 ;
      RECT 0.11 0.23 0.27 0.53 ;
      RECT 0.335 1.195 0.755 1.295 ;
      RECT 0.49 1.42 0.96 1.52 ;
      RECT 0.82 1.62 0.98 1.92 ;
      RECT 0.82 0.23 0.98 0.53 ;
      RECT 0.58 0.63 1.08 0.73 ;
      RECT 1.06 1.42 1.54 1.52 ;
      RECT 1.52 1.62 1.68 1.92 ;
      RECT 1.52 0.23 1.68 0.53 ;
      RECT 0.23 0.945 1.92 1.045 ;
      RECT 0.74 0.93 1.07 1.06 ;
      RECT 1.77 1.62 1.93 1.92 ;
      RECT 1.77 0.23 1.93 0.53 ;
      RECT 2.25 1.62 2.41 1.92 ;
      RECT 2.25 0.23 2.41 0.53 ;
      RECT 1.17 0.63 2.12 0.73 ;
      RECT 2.02 0.63 2.12 0.93 ;
      RECT 2.02 0.83 2.78 0.93 ;
      RECT 2.63 1.42 3.1 1.52 ;
      RECT 2.96 1.62 3.12 1.92 ;
      RECT 2.96 0.23 3.12 0.53 ;
      RECT 1.91 1.15 3.21 1.25 ;
      RECT 2.88 1.135 3.21 1.265 ;
      RECT 2.72 0.63 3.22 0.73 ;
      RECT 3.2 1.42 3.68 1.52 ;
      RECT 3.67 1.62 3.83 1.92 ;
      RECT 3.57 1.18 3.99 1.28 ;
      RECT 3.32 0.63 4.02 0.73 ;
      RECT 3.86 0.23 4.02 0.53 ;
      RECT 0.405 1.62 0.495 2.52 ;
      RECT 1.305 1.62 1.395 2.52 ;
      RECT 2.055 1.62 2.145 2.52 ;
      RECT 2.545 1.62 2.635 2.52 ;
      RECT 3.445 1.62 3.535 2.52 ;
      RECT 3.965 1.62 4.055 2.52 ;
      RECT 0 2.3 4.2 2.52 ;
      RECT 0 -0.22 4.2 0 ;
      RECT 0.405 -0.22 0.495 0.53 ;
      RECT 1.305 -0.22 1.395 0.53 ;
      RECT 2.055 -0.22 2.145 0.53 ;
      RECT 2.545 -0.22 2.635 0.53 ;
      RECT 3.445 -0.22 3.535 0.53 ;
    LAYER VI1 ;
      RECT 0.14 1.72 0.24 1.82 ;
      RECT 0.14 0.4 0.24 0.5 ;
      RECT 0.61 1.42 0.71 1.52 ;
      RECT 0.61 0.63 0.71 0.73 ;
      RECT 0.85 1.72 0.95 1.82 ;
      RECT 0.85 0.4 0.95 0.5 ;
      RECT 1.09 1.42 1.19 1.52 ;
      RECT 1.56 1.72 1.66 1.82 ;
      RECT 1.56 0.63 1.66 0.73 ;
      RECT 1.56 0.4 1.66 0.5 ;
      RECT 1.79 1.72 1.89 1.82 ;
      RECT 1.79 0.945 1.89 1.045 ;
      RECT 1.79 0.4 1.89 0.5 ;
      RECT 2.28 1.72 2.38 1.82 ;
      RECT 2.28 0.4 2.38 0.5 ;
      RECT 2.75 1.42 2.85 1.52 ;
      RECT 2.75 0.63 2.85 0.73 ;
      RECT 2.99 1.72 3.09 1.82 ;
      RECT 2.99 0.4 3.09 0.5 ;
      RECT 3.23 1.42 3.33 1.52 ;
      RECT 3.7 1.72 3.8 1.82 ;
      RECT 3.89 0.63 3.99 0.73 ;
      RECT 3.89 0.4 3.99 0.5 ;
    LAYER ME2 ;
      RECT 0.14 0.63 0.74 0.73 ;
      RECT 0.14 1.42 0.74 1.52 ;
      RECT 0.14 0.37 0.24 1.92 ;
      RECT 0.85 1.42 1.22 1.52 ;
      RECT 0.85 0.37 0.95 1.92 ;
      RECT 1.56 0.37 1.66 1.92 ;
      RECT 1.79 0.37 1.89 1.92 ;
      RECT 2.28 0.63 2.88 0.73 ;
      RECT 2.28 1.42 2.88 1.52 ;
      RECT 2.28 0.37 2.38 1.92 ;
      RECT 2.99 1.42 3.36 1.52 ;
      RECT 2.99 0.37 3.09 1.92 ;
      RECT 3.89 0.37 3.99 1.72 ;
      RECT 3.7 1.62 3.99 1.72 ;
      RECT 3.7 1.62 3.8 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDFFCNSX1

MACRO QDFFCRX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDFFCRX1 0 -0.11 ;
  SIZE 4.2 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 1.91 1.15 3.21 1.25 ;
        RECT 2.88 1.135 3.21 1.265 ;
    END
  END CLK
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.405 1.62 0.495 2.52 ;
        RECT 1.305 1.62 1.395 2.52 ;
        RECT 2.055 1.62 2.145 2.52 ;
        RECT 2.545 1.62 2.635 2.52 ;
        RECT 3.445 1.62 3.535 2.52 ;
        RECT 0 2.3 4.2 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.405 -0.22 0.495 0.53 ;
        RECT 1.305 -0.22 1.395 0.53 ;
        RECT 2.055 -0.22 2.145 0.53 ;
        RECT 2.545 -0.22 2.635 0.53 ;
        RECT 3.445 -0.22 3.535 0.53 ;
        RECT 3.965 -0.22 4.055 0.53 ;
        RECT 0 -0.22 4.2 0 ;
    END
  END gnd!
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 3.57 1.185 3.99 1.285 ;
    END
  END RST
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.22 1.19 0.64 1.29 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 3.7 0.4 3.8 0.5 ;
        RECT 3.89 1.72 3.99 1.82 ;
        RECT 3.89 0.63 3.99 0.73 ;
      LAYER ME1 ;
        RECT 3.32 0.63 4.02 0.73 ;
        RECT 3.86 1.62 4.02 1.92 ;
        RECT 3.67 0.23 3.83 0.53 ;
      LAYER ME2 ;
        RECT 3.89 0.43 3.99 1.92 ;
        RECT 3.7 0.43 3.99 0.53 ;
        RECT 3.7 0.37 3.8 0.53 ;
    END
  END Q
  OBS
    LAYER ME1 ;
      RECT 0.11 1.62 0.27 1.92 ;
      RECT 0.11 0.23 0.27 0.53 ;
      RECT 0.22 1.19 0.64 1.29 ;
      RECT 0.49 1.42 0.96 1.52 ;
      RECT 0.82 1.62 0.98 1.92 ;
      RECT 0.82 0.23 0.98 0.53 ;
      RECT 0.58 0.63 1.08 0.73 ;
      RECT 1.06 1.15 1.54 1.25 ;
      RECT 1.52 1.62 1.68 1.92 ;
      RECT 1.52 0.23 1.68 0.53 ;
      RECT 0.23 0.945 1.92 1.045 ;
      RECT 0.74 0.93 1.07 1.06 ;
      RECT 1.77 1.62 1.93 1.92 ;
      RECT 1.77 0.23 1.93 0.53 ;
      RECT 2.25 1.62 2.41 1.92 ;
      RECT 2.25 0.23 2.41 0.53 ;
      RECT 1.17 0.63 2.12 0.73 ;
      RECT 2.02 0.63 2.12 0.93 ;
      RECT 2.02 0.83 2.78 0.93 ;
      RECT 2.25 1.42 3.1 1.52 ;
      RECT 2.96 1.62 3.12 1.92 ;
      RECT 2.96 0.23 3.12 0.53 ;
      RECT 1.91 1.15 3.21 1.25 ;
      RECT 2.88 1.135 3.21 1.265 ;
      RECT 2.25 0.63 3.22 0.73 ;
      RECT 3.2 1.42 3.68 1.52 ;
      RECT 3.67 0.23 3.83 0.53 ;
      RECT 3.57 1.185 3.99 1.285 ;
      RECT 3.86 1.62 4.02 1.92 ;
      RECT 3.32 0.63 4.02 0.73 ;
      RECT 0.405 1.62 0.495 2.52 ;
      RECT 1.305 1.62 1.395 2.52 ;
      RECT 2.055 1.62 2.145 2.52 ;
      RECT 2.545 1.62 2.635 2.52 ;
      RECT 3.445 1.62 3.535 2.52 ;
      RECT 0 2.3 4.2 2.52 ;
      RECT 0 -0.22 4.2 0 ;
      RECT 0.405 -0.22 0.495 0.53 ;
      RECT 1.305 -0.22 1.395 0.53 ;
      RECT 2.055 -0.22 2.145 0.53 ;
      RECT 2.545 -0.22 2.635 0.53 ;
      RECT 3.445 -0.22 3.535 0.53 ;
      RECT 3.965 -0.22 4.055 0.53 ;
    LAYER VI1 ;
      RECT 0.14 1.72 0.24 1.82 ;
      RECT 0.14 0.4 0.24 0.5 ;
      RECT 0.61 1.42 0.71 1.52 ;
      RECT 0.61 0.63 0.71 0.73 ;
      RECT 0.85 1.72 0.95 1.82 ;
      RECT 0.85 0.4 0.95 0.5 ;
      RECT 1.09 1.15 1.19 1.25 ;
      RECT 1.56 1.72 1.66 1.82 ;
      RECT 1.56 0.63 1.66 0.73 ;
      RECT 1.56 0.4 1.66 0.5 ;
      RECT 1.79 1.72 1.89 1.82 ;
      RECT 1.79 0.945 1.89 1.045 ;
      RECT 1.79 0.4 1.89 0.5 ;
      RECT 2.28 1.72 2.38 1.82 ;
      RECT 2.28 1.42 2.38 1.52 ;
      RECT 2.28 0.63 2.38 0.73 ;
      RECT 2.28 0.4 2.38 0.5 ;
      RECT 2.99 1.72 3.09 1.82 ;
      RECT 2.99 0.4 3.09 0.5 ;
      RECT 3.23 1.42 3.33 1.52 ;
      RECT 3.7 0.4 3.8 0.5 ;
      RECT 3.89 1.72 3.99 1.82 ;
      RECT 3.89 0.63 3.99 0.73 ;
    LAYER ME2 ;
      RECT 0.14 0.63 0.74 0.73 ;
      RECT 0.14 1.42 0.74 1.52 ;
      RECT 0.14 0.37 0.24 1.92 ;
      RECT 0.85 1.15 1.22 1.25 ;
      RECT 0.85 0.37 0.95 1.92 ;
      RECT 1.56 0.37 1.66 1.92 ;
      RECT 1.79 0.37 1.89 1.92 ;
      RECT 2.28 0.37 2.38 1.92 ;
      RECT 2.99 1.42 3.36 1.52 ;
      RECT 2.99 0.37 3.09 1.92 ;
      RECT 3.7 0.37 3.8 0.53 ;
      RECT 3.7 0.43 3.99 0.53 ;
      RECT 3.89 0.43 3.99 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDFFCRX1

MACRO QDFFCSRX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDFFCSRX1 0 -0.11 ;
  SIZE 5.32 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.46 1.62 0.55 2.52 ;
        RECT 1.36 1.62 1.45 2.52 ;
        RECT 2.11 1.62 2.2 2.52 ;
        RECT 2.6 1.62 2.69 2.52 ;
        RECT 3.5 1.62 3.59 2.52 ;
        RECT 4.77 1.62 4.86 2.52 ;
        RECT 0 2.3 5.32 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.46 -0.22 0.55 0.53 ;
        RECT 1.36 -0.22 1.45 0.53 ;
        RECT 2.11 -0.22 2.2 0.53 ;
        RECT 2.6 -0.22 2.69 0.53 ;
        RECT 3.5 -0.22 3.59 0.53 ;
        RECT 4.02 -0.22 4.11 0.53 ;
        RECT 4.25 -0.22 4.34 0.53 ;
        RECT 4.77 -0.22 4.86 0.53 ;
        RECT 0 -0.22 5.32 0 ;
    END
  END gnd!
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 3.625 0.915 4.045 1.015 ;
    END
  END RST
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.41 1.18 0.83 1.28 ;
    END
  END D
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 4.375 1.085 4.795 1.185 ;
    END
  END SET
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 4.745 0.63 4.845 0.73 ;
        RECT 5.025 1.72 5.125 1.82 ;
        RECT 5.025 0.4 5.125 0.5 ;
      LAYER ME1 ;
        RECT 4.995 1.62 5.155 1.92 ;
        RECT 4.975 0.23 5.135 0.53 ;
        RECT 3.375 0.63 4.875 0.73 ;
      LAYER ME2 ;
        RECT 5.025 0.23 5.125 1.92 ;
        RECT 4.715 0.63 5.125 0.73 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 1.965 0.915 3.265 1.015 ;
        RECT 2.935 0.9 3.265 1.03 ;
    END
  END CLK
  OBS
    LAYER ME1 ;
      RECT 0.165 1.62 0.325 1.92 ;
      RECT 0.165 0.23 0.325 0.53 ;
      RECT 0.41 1.18 0.83 1.28 ;
      RECT 0.545 1.42 1.015 1.52 ;
      RECT 0.875 1.62 1.035 1.92 ;
      RECT 0.875 0.23 1.035 0.53 ;
      RECT 0.635 0.63 1.135 0.73 ;
      RECT 1.115 1.42 1.595 1.52 ;
      RECT 1.575 1.62 1.735 1.92 ;
      RECT 1.575 0.23 1.735 0.53 ;
      RECT 1.685 0.685 1.975 0.785 ;
      RECT 1.685 0.685 1.785 1.015 ;
      RECT 0.285 0.915 1.785 1.015 ;
      RECT 0.795 0.9 1.125 1.03 ;
      RECT 1.825 1.62 1.985 1.92 ;
      RECT 1.825 0.23 1.985 0.53 ;
      RECT 2.305 1.62 2.465 1.92 ;
      RECT 2.305 0.23 2.465 0.53 ;
      RECT 1.225 1.13 2.835 1.23 ;
      RECT 2.685 1.42 3.155 1.52 ;
      RECT 3.015 1.62 3.175 1.92 ;
      RECT 3.015 0.23 3.175 0.53 ;
      RECT 1.965 0.915 3.265 1.015 ;
      RECT 2.935 0.9 3.265 1.03 ;
      RECT 2.775 0.63 3.275 0.73 ;
      RECT 3.255 1.42 3.735 1.52 ;
      RECT 3.725 0.23 3.885 0.53 ;
      RECT 3.625 0.915 4.045 1.015 ;
      RECT 3.915 1.62 4.075 1.92 ;
      RECT 4.285 1.62 4.445 1.92 ;
      RECT 3.915 1.325 4.535 1.425 ;
      RECT 4.475 0.23 4.635 0.53 ;
      RECT 4.375 1.085 4.795 1.185 ;
      RECT 3.375 0.63 4.875 0.73 ;
      RECT 4.285 0.835 5.005 0.925 ;
      RECT 4.285 0.83 4.445 0.93 ;
      RECT 4.975 0.23 5.135 0.53 ;
      RECT 4.995 1.62 5.155 1.92 ;
      RECT 0.46 1.62 0.55 2.52 ;
      RECT 1.36 1.62 1.45 2.52 ;
      RECT 2.11 1.62 2.2 2.52 ;
      RECT 2.6 1.62 2.69 2.52 ;
      RECT 3.5 1.62 3.59 2.52 ;
      RECT 4.77 1.62 4.86 2.52 ;
      RECT 0 2.3 5.32 2.52 ;
      RECT 0 -0.22 5.32 0 ;
      RECT 0.46 -0.22 0.55 0.53 ;
      RECT 1.36 -0.22 1.45 0.53 ;
      RECT 2.11 -0.22 2.2 0.53 ;
      RECT 2.6 -0.22 2.69 0.53 ;
      RECT 3.5 -0.22 3.59 0.53 ;
      RECT 4.02 -0.22 4.11 0.53 ;
      RECT 4.25 -0.22 4.34 0.53 ;
      RECT 4.77 -0.22 4.86 0.53 ;
    LAYER VI1 ;
      RECT 0.195 1.72 0.295 1.82 ;
      RECT 0.195 0.4 0.295 0.5 ;
      RECT 0.665 1.42 0.765 1.52 ;
      RECT 0.665 0.63 0.765 0.73 ;
      RECT 0.905 1.72 1.005 1.82 ;
      RECT 0.905 0.4 1.005 0.5 ;
      RECT 1.145 1.42 1.245 1.52 ;
      RECT 1.615 1.72 1.715 1.82 ;
      RECT 1.615 1.13 1.715 1.23 ;
      RECT 1.615 0.4 1.715 0.5 ;
      RECT 1.845 1.72 1.945 1.82 ;
      RECT 1.845 0.685 1.945 0.785 ;
      RECT 1.845 0.4 1.945 0.5 ;
      RECT 2.335 1.72 2.435 1.82 ;
      RECT 2.335 0.4 2.435 0.5 ;
      RECT 2.805 1.42 2.905 1.52 ;
      RECT 2.805 0.63 2.905 0.73 ;
      RECT 3.045 1.72 3.145 1.82 ;
      RECT 3.045 0.4 3.145 0.5 ;
      RECT 3.285 1.42 3.385 1.52 ;
      RECT 3.755 0.4 3.855 0.5 ;
      RECT 3.945 1.72 4.045 1.82 ;
      RECT 3.945 1.325 4.045 1.425 ;
      RECT 4.315 1.72 4.415 1.82 ;
      RECT 4.315 0.83 4.415 0.93 ;
      RECT 4.505 0.4 4.605 0.5 ;
      RECT 4.745 0.63 4.845 0.73 ;
      RECT 5.025 1.72 5.125 1.82 ;
      RECT 5.025 0.4 5.125 0.5 ;
    LAYER ME2 ;
      RECT 0.195 0.63 0.795 0.73 ;
      RECT 0.195 1.42 0.795 1.52 ;
      RECT 0.195 0.37 0.295 1.92 ;
      RECT 0.905 1.42 1.275 1.52 ;
      RECT 0.905 0.37 1.005 1.92 ;
      RECT 1.615 0.23 1.715 1.92 ;
      RECT 1.845 0.37 1.945 1.92 ;
      RECT 2.335 0.63 2.935 0.73 ;
      RECT 2.335 1.42 2.935 1.52 ;
      RECT 2.335 0.37 2.435 1.92 ;
      RECT 3.045 1.42 3.415 1.52 ;
      RECT 3.045 0.37 3.145 1.92 ;
      RECT 3.755 0.37 3.855 0.53 ;
      RECT 3.755 0.43 4.045 0.53 ;
      RECT 3.945 0.43 4.045 1.92 ;
      RECT 4.505 0.37 4.605 0.53 ;
      RECT 4.315 0.43 4.605 0.53 ;
      RECT 4.315 0.43 4.415 1.92 ;
      RECT 4.715 0.63 5.125 0.73 ;
      RECT 5.025 0.23 5.125 1.92 ;
  END
END QDFFCSRX1

MACRO QDFFCX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDFFCX1 0 -0.11 ;
  SIZE 4.2 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.235 1.62 0.325 2.52 ;
        RECT 1.025 1.62 1.115 2.52 ;
        RECT 1.925 1.62 2.015 2.52 ;
        RECT 2.715 1.62 2.805 2.52 ;
        RECT 3.615 1.62 3.705 2.52 ;
        RECT 0 2.3 4.2 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.235 -0.22 0.325 0.53 ;
        RECT 1.025 -0.22 1.115 0.53 ;
        RECT 1.925 -0.22 2.015 0.53 ;
        RECT 2.715 -0.22 2.805 0.53 ;
        RECT 3.615 -0.22 3.705 0.53 ;
        RECT 0 -0.22 4.2 0 ;
    END
  END gnd!
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.23 0.83 2.66 0.93 ;
        RECT 1.845 0.915 3.39 1.015 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 3.87 1.72 3.97 1.82 ;
        RECT 3.87 0.63 3.97 0.73 ;
        RECT 3.87 0.4 3.97 0.5 ;
      LAYER ME1 ;
        RECT 3.84 0.23 4 0.53 ;
        RECT 3.49 0.63 4 0.73 ;
        RECT 3.84 1.62 4 1.92 ;
      LAYER ME2 ;
        RECT 3.87 0.37 3.97 1.92 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.23 1.225 1.26 1.325 ;
    END
  END D
  OBS
    LAYER ME1 ;
      RECT 0.46 1.62 0.62 1.92 ;
      RECT 0.46 0.23 0.62 0.53 ;
      RECT 0.73 1.62 0.89 1.92 ;
      RECT 0.73 0.23 0.89 0.53 ;
      RECT 0.23 1.225 1.26 1.325 ;
      RECT 1.16 1.425 1.58 1.525 ;
      RECT 1.44 1.62 1.6 1.92 ;
      RECT 1.44 0.23 1.6 0.53 ;
      RECT 0.46 1.025 1.7 1.125 ;
      RECT 1.2 0.63 1.71 0.73 ;
      RECT 1.68 1.425 2.16 1.525 ;
      RECT 2.15 1.62 2.31 1.92 ;
      RECT 1.8 0.63 2.31 0.73 ;
      RECT 2.15 0.23 2.31 0.53 ;
      RECT 2.42 1.62 2.58 1.92 ;
      RECT 2.42 0.23 2.58 0.53 ;
      RECT 2.15 1.13 2.95 1.23 ;
      RECT 2.85 1.425 3.27 1.525 ;
      RECT 3.13 1.62 3.29 1.92 ;
      RECT 3.13 0.23 3.29 0.53 ;
      RECT 0.23 0.83 2.66 0.93 ;
      RECT 1.845 0.915 3.39 1.015 ;
      RECT 2.89 0.63 3.4 0.73 ;
      RECT 3.37 1.12 3.85 1.22 ;
      RECT 3.84 1.62 4 1.92 ;
      RECT 3.49 0.63 4 0.73 ;
      RECT 3.84 0.23 4 0.53 ;
      RECT 0.235 1.62 0.325 2.52 ;
      RECT 1.025 1.62 1.115 2.52 ;
      RECT 1.925 1.62 2.015 2.52 ;
      RECT 2.715 1.62 2.805 2.52 ;
      RECT 3.615 1.62 3.705 2.52 ;
      RECT 0 2.3 4.2 2.52 ;
      RECT 0 -0.22 4.2 0 ;
      RECT 0.235 -0.22 0.325 0.53 ;
      RECT 1.025 -0.22 1.115 0.53 ;
      RECT 1.925 -0.22 2.015 0.53 ;
      RECT 2.715 -0.22 2.805 0.53 ;
      RECT 3.615 -0.22 3.705 0.53 ;
    LAYER VI1 ;
      RECT 0.49 1.72 0.59 1.82 ;
      RECT 0.49 1.025 0.59 1.125 ;
      RECT 0.49 0.4 0.59 0.5 ;
      RECT 0.76 1.72 0.86 1.82 ;
      RECT 0.76 0.4 0.86 0.5 ;
      RECT 1.23 1.425 1.33 1.525 ;
      RECT 1.23 0.63 1.33 0.73 ;
      RECT 1.47 1.72 1.57 1.82 ;
      RECT 1.47 0.4 1.57 0.5 ;
      RECT 1.71 1.425 1.81 1.525 ;
      RECT 2.18 1.72 2.28 1.82 ;
      RECT 2.18 1.13 2.28 1.23 ;
      RECT 2.18 0.63 2.28 0.73 ;
      RECT 2.18 0.4 2.28 0.5 ;
      RECT 2.45 1.72 2.55 1.82 ;
      RECT 2.45 0.4 2.55 0.5 ;
      RECT 2.92 1.425 3.02 1.525 ;
      RECT 2.92 0.63 3.02 0.73 ;
      RECT 3.16 1.72 3.26 1.82 ;
      RECT 3.16 0.4 3.26 0.5 ;
      RECT 3.4 1.12 3.5 1.22 ;
      RECT 3.87 1.72 3.97 1.82 ;
      RECT 3.87 0.63 3.97 0.73 ;
      RECT 3.87 0.4 3.97 0.5 ;
    LAYER ME2 ;
      RECT 0.49 0.37 0.59 1.92 ;
      RECT 0.76 0.63 1.36 0.73 ;
      RECT 0.76 1.425 1.36 1.525 ;
      RECT 0.76 0.37 0.86 1.92 ;
      RECT 1.47 1.425 1.84 1.525 ;
      RECT 1.47 0.37 1.57 1.92 ;
      RECT 2.18 0.37 2.28 1.92 ;
      RECT 2.45 0.63 3.05 0.73 ;
      RECT 2.45 1.425 3.05 1.525 ;
      RECT 2.45 0.37 2.55 1.92 ;
      RECT 3.16 1.12 3.53 1.22 ;
      RECT 3.16 0.37 3.26 1.92 ;
      RECT 3.87 0.37 3.97 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDFFCX1

MACRO QDFFNCNSX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDFFNCNSX1 0 -0.11 ;
  SIZE 4.2 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 3.57 1.42 3.99 1.52 ;
    END
  END SETB
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.405 1.62 0.495 2.52 ;
        RECT 1.305 1.62 1.395 2.52 ;
        RECT 2.055 1.62 2.145 2.52 ;
        RECT 2.545 1.62 2.635 2.52 ;
        RECT 3.445 1.62 3.535 2.52 ;
        RECT 3.965 1.62 4.055 2.52 ;
        RECT 0 2.3 4.2 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.405 -0.22 0.495 0.53 ;
        RECT 1.305 -0.22 1.395 0.53 ;
        RECT 2.055 -0.22 2.145 0.53 ;
        RECT 2.545 -0.22 2.635 0.53 ;
        RECT 3.445 -0.22 3.535 0.53 ;
        RECT 0 -0.22 4.2 0 ;
    END
  END gnd!
  PIN CLKB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 1.91 1.15 3.21 1.25 ;
        RECT 2.88 1.135 3.21 1.265 ;
    END
  END CLKB
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.335 1.19 0.755 1.29 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 3.7 1.72 3.8 1.82 ;
        RECT 3.89 0.63 3.99 0.73 ;
        RECT 3.89 0.4 3.99 0.5 ;
      LAYER ME1 ;
        RECT 3.86 0.23 4.02 0.53 ;
        RECT 3.31 0.63 4.02 0.73 ;
        RECT 3.67 1.62 3.83 1.92 ;
      LAYER ME2 ;
        RECT 3.7 1.62 3.99 1.72 ;
        RECT 3.89 0.37 3.99 1.72 ;
        RECT 3.7 1.62 3.8 1.92 ;
    END
  END Q
  OBS
    LAYER ME1 ;
      RECT 0.11 1.62 0.27 1.92 ;
      RECT 0.11 0.23 0.27 0.53 ;
      RECT 0.335 1.19 0.755 1.29 ;
      RECT 0.45 0.63 0.87 0.73 ;
      RECT 0.82 1.62 0.98 1.92 ;
      RECT 0.82 0.23 0.98 0.53 ;
      RECT 0.49 1.42 1.09 1.52 ;
      RECT 1.23 1.42 1.65 1.52 ;
      RECT 1.52 1.62 1.68 1.92 ;
      RECT 1.52 0.23 1.68 0.53 ;
      RECT 0.23 0.945 1.92 1.045 ;
      RECT 0.74 0.93 1.07 1.06 ;
      RECT 1.77 1.62 1.93 1.92 ;
      RECT 1.77 0.23 1.93 0.53 ;
      RECT 2.25 1.62 2.41 1.92 ;
      RECT 2.25 0.23 2.41 0.53 ;
      RECT 1.17 0.63 2.12 0.73 ;
      RECT 2.02 0.63 2.12 0.93 ;
      RECT 2.02 0.83 2.78 0.93 ;
      RECT 2.25 0.63 3.01 0.73 ;
      RECT 2.96 1.62 3.12 1.92 ;
      RECT 2.96 0.23 3.12 0.53 ;
      RECT 1.91 1.15 3.21 1.25 ;
      RECT 2.88 1.135 3.21 1.265 ;
      RECT 2.25 1.42 3.23 1.52 ;
      RECT 3.2 0.89 3.68 0.99 ;
      RECT 3.67 1.62 3.83 1.92 ;
      RECT 3.57 1.42 3.99 1.52 ;
      RECT 3.31 0.63 4.02 0.73 ;
      RECT 3.86 0.23 4.02 0.53 ;
      RECT 0.405 1.62 0.495 2.52 ;
      RECT 1.305 1.62 1.395 2.52 ;
      RECT 2.055 1.62 2.145 2.52 ;
      RECT 2.545 1.62 2.635 2.52 ;
      RECT 3.445 1.62 3.535 2.52 ;
      RECT 3.965 1.62 4.055 2.52 ;
      RECT 0 2.3 4.2 2.52 ;
      RECT 0 -0.22 4.2 0 ;
      RECT 0.405 -0.22 0.495 0.53 ;
      RECT 1.305 -0.22 1.395 0.53 ;
      RECT 2.055 -0.22 2.145 0.53 ;
      RECT 2.545 -0.22 2.635 0.53 ;
      RECT 3.445 -0.22 3.535 0.53 ;
    LAYER VI1 ;
      RECT 0.14 1.72 0.24 1.82 ;
      RECT 0.14 0.4 0.24 0.5 ;
      RECT 0.48 0.63 0.58 0.73 ;
      RECT 0.61 1.42 0.71 1.52 ;
      RECT 0.85 1.72 0.95 1.82 ;
      RECT 0.85 0.4 0.95 0.5 ;
      RECT 1.26 1.42 1.36 1.52 ;
      RECT 1.56 1.72 1.66 1.82 ;
      RECT 1.56 0.63 1.66 0.73 ;
      RECT 1.56 0.4 1.66 0.5 ;
      RECT 1.79 1.72 1.89 1.82 ;
      RECT 1.79 0.945 1.89 1.045 ;
      RECT 1.79 0.4 1.89 0.5 ;
      RECT 2.28 1.72 2.38 1.82 ;
      RECT 2.28 1.42 2.38 1.52 ;
      RECT 2.28 0.63 2.38 0.73 ;
      RECT 2.28 0.4 2.38 0.5 ;
      RECT 2.99 1.72 3.09 1.82 ;
      RECT 2.99 0.4 3.09 0.5 ;
      RECT 3.23 0.89 3.33 0.99 ;
      RECT 3.7 1.72 3.8 1.82 ;
      RECT 3.89 0.63 3.99 0.73 ;
      RECT 3.89 0.4 3.99 0.5 ;
    LAYER ME2 ;
      RECT 0.14 0.63 0.61 0.73 ;
      RECT 0.14 1.42 0.74 1.52 ;
      RECT 0.14 0.37 0.24 1.92 ;
      RECT 0.85 1.42 1.39 1.52 ;
      RECT 0.85 0.37 0.95 1.92 ;
      RECT 1.56 0.37 1.66 1.92 ;
      RECT 1.79 0.37 1.89 1.92 ;
      RECT 2.28 0.37 2.38 1.92 ;
      RECT 2.99 0.89 3.36 0.99 ;
      RECT 2.99 0.37 3.09 1.92 ;
      RECT 3.89 0.37 3.99 1.72 ;
      RECT 3.7 1.62 3.99 1.72 ;
      RECT 3.7 1.62 3.8 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDFFNCNSX1

MACRO QDFFNCRX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDFFNCRX1 0 -0.11 ;
  SIZE 4.2 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 3.7 0.4 3.8 0.5 ;
        RECT 3.89 1.72 3.99 1.82 ;
        RECT 3.89 0.63 3.99 0.73 ;
      LAYER ME2 ;
        RECT 3.89 0.43 3.99 1.92 ;
        RECT 3.7 0.43 3.99 0.53 ;
        RECT 3.7 0.37 3.8 0.53 ;
      LAYER ME1 ;
        RECT 3.32 0.63 4.02 0.73 ;
        RECT 3.86 1.62 4.02 1.92 ;
        RECT 3.67 0.23 3.83 0.53 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.405 1.62 0.495 2.52 ;
        RECT 1.305 1.62 1.395 2.52 ;
        RECT 2.055 1.62 2.145 2.52 ;
        RECT 2.545 1.62 2.635 2.52 ;
        RECT 3.445 1.62 3.535 2.52 ;
        RECT 0 2.3 4.2 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.405 -0.22 0.495 0.53 ;
        RECT 1.305 -0.22 1.395 0.53 ;
        RECT 2.055 -0.22 2.145 0.53 ;
        RECT 2.545 -0.22 2.635 0.53 ;
        RECT 3.445 -0.22 3.535 0.53 ;
        RECT 3.965 -0.22 4.055 0.53 ;
        RECT 0 -0.22 4.2 0 ;
    END
  END gnd!
  PIN CLKB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 1.91 1.15 3.21 1.25 ;
        RECT 2.88 1.135 3.21 1.265 ;
    END
  END CLKB
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.345 1.17 0.765 1.27 ;
    END
  END D
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 3.57 1.185 3.99 1.285 ;
    END
  END RST
  OBS
    LAYER ME1 ;
      RECT 0.11 1.62 0.27 1.92 ;
      RECT 0.11 0.23 0.27 0.53 ;
      RECT 0.345 1.17 0.765 1.27 ;
      RECT 0.45 0.63 0.87 0.73 ;
      RECT 0.82 1.62 0.98 1.92 ;
      RECT 0.82 0.23 0.98 0.53 ;
      RECT 0.49 1.42 1.09 1.52 ;
      RECT 1.23 1.42 1.65 1.52 ;
      RECT 1.52 1.62 1.68 1.92 ;
      RECT 1.52 0.23 1.68 0.53 ;
      RECT 0.23 0.945 1.92 1.045 ;
      RECT 0.74 0.93 1.07 1.06 ;
      RECT 1.77 1.62 1.93 1.92 ;
      RECT 1.77 0.23 1.93 0.53 ;
      RECT 2.25 1.62 2.41 1.92 ;
      RECT 2.25 0.23 2.41 0.53 ;
      RECT 1.17 0.63 2.12 0.73 ;
      RECT 2.02 0.63 2.12 0.93 ;
      RECT 2.02 0.83 2.78 0.93 ;
      RECT 2.25 0.63 3.01 0.73 ;
      RECT 2.96 1.62 3.12 1.92 ;
      RECT 2.96 0.23 3.12 0.53 ;
      RECT 1.91 1.15 3.21 1.25 ;
      RECT 2.88 1.135 3.21 1.265 ;
      RECT 2.25 1.42 3.23 1.52 ;
      RECT 3.37 1.42 3.79 1.52 ;
      RECT 3.67 0.23 3.83 0.53 ;
      RECT 3.57 1.185 3.99 1.285 ;
      RECT 3.86 1.62 4.02 1.92 ;
      RECT 3.32 0.63 4.02 0.73 ;
      RECT 0.405 1.62 0.495 2.52 ;
      RECT 1.305 1.62 1.395 2.52 ;
      RECT 2.055 1.62 2.145 2.52 ;
      RECT 2.545 1.62 2.635 2.52 ;
      RECT 3.445 1.62 3.535 2.52 ;
      RECT 0 2.3 4.2 2.52 ;
      RECT 0 -0.22 4.2 0 ;
      RECT 0.405 -0.22 0.495 0.53 ;
      RECT 1.305 -0.22 1.395 0.53 ;
      RECT 2.055 -0.22 2.145 0.53 ;
      RECT 2.545 -0.22 2.635 0.53 ;
      RECT 3.445 -0.22 3.535 0.53 ;
      RECT 3.965 -0.22 4.055 0.53 ;
    LAYER VI1 ;
      RECT 0.14 1.72 0.24 1.82 ;
      RECT 0.14 0.4 0.24 0.5 ;
      RECT 0.48 0.63 0.58 0.73 ;
      RECT 0.61 1.42 0.71 1.52 ;
      RECT 0.85 1.72 0.95 1.82 ;
      RECT 0.85 0.4 0.95 0.5 ;
      RECT 1.26 1.42 1.36 1.52 ;
      RECT 1.56 1.72 1.66 1.82 ;
      RECT 1.56 0.63 1.66 0.73 ;
      RECT 1.56 0.4 1.66 0.5 ;
      RECT 1.79 1.72 1.89 1.82 ;
      RECT 1.79 0.945 1.89 1.045 ;
      RECT 1.79 0.4 1.89 0.5 ;
      RECT 2.28 1.72 2.38 1.82 ;
      RECT 2.28 1.42 2.38 1.52 ;
      RECT 2.28 0.63 2.38 0.73 ;
      RECT 2.28 0.4 2.38 0.5 ;
      RECT 2.99 1.72 3.09 1.82 ;
      RECT 2.99 0.4 3.09 0.5 ;
      RECT 3.4 1.42 3.5 1.52 ;
      RECT 3.7 0.4 3.8 0.5 ;
      RECT 3.89 1.72 3.99 1.82 ;
      RECT 3.89 0.63 3.99 0.73 ;
    LAYER ME2 ;
      RECT 0.14 0.63 0.61 0.73 ;
      RECT 0.14 1.42 0.74 1.52 ;
      RECT 0.14 0.37 0.24 1.92 ;
      RECT 0.85 1.42 1.39 1.52 ;
      RECT 0.85 0.37 0.95 1.92 ;
      RECT 1.56 0.37 1.66 1.92 ;
      RECT 1.79 0.37 1.89 1.92 ;
      RECT 2.28 0.37 2.38 1.92 ;
      RECT 2.99 1.42 3.53 1.52 ;
      RECT 2.99 0.37 3.09 1.92 ;
      RECT 3.7 0.37 3.8 0.53 ;
      RECT 3.7 0.43 3.99 0.53 ;
      RECT 3.89 0.43 3.99 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDFFNCRX1

MACRO QDFFNCSRX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDFFNCSRX1 0 -0.11 ;
  SIZE 5.32 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.46 1.62 0.55 2.52 ;
        RECT 1.36 1.62 1.45 2.52 ;
        RECT 2.11 1.62 2.2 2.52 ;
        RECT 2.6 1.62 2.69 2.52 ;
        RECT 3.5 1.62 3.59 2.52 ;
        RECT 4.77 1.62 4.86 2.52 ;
        RECT 0 2.3 5.32 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.46 -0.22 0.55 0.53 ;
        RECT 1.36 -0.22 1.45 0.53 ;
        RECT 2.11 -0.22 2.2 0.53 ;
        RECT 2.6 -0.22 2.69 0.53 ;
        RECT 3.5 -0.22 3.59 0.53 ;
        RECT 4.02 -0.22 4.11 0.53 ;
        RECT 4.25 -0.22 4.34 0.53 ;
        RECT 4.77 -0.22 4.86 0.53 ;
        RECT 0 -0.22 5.32 0 ;
    END
  END gnd!
  PIN CLKB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 1.965 1.15 3.265 1.25 ;
        RECT 2.935 1.135 3.265 1.265 ;
    END
  END CLKB
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 3.625 0.915 4.045 1.015 ;
    END
  END RST
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 4.375 1.085 4.795 1.185 ;
    END
  END SET
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 4.745 0.63 4.845 0.73 ;
        RECT 5.025 1.72 5.125 1.82 ;
        RECT 5.025 0.4 5.125 0.5 ;
      LAYER ME1 ;
        RECT 4.995 1.62 5.155 1.92 ;
        RECT 4.975 0.23 5.135 0.53 ;
        RECT 3.375 0.63 4.875 0.73 ;
      LAYER ME2 ;
        RECT 5.025 0.23 5.125 1.92 ;
        RECT 4.715 0.63 5.125 0.73 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.375 1.17 0.795 1.27 ;
    END
  END D
  OBS
    LAYER ME1 ;
      RECT 0.165 1.62 0.325 1.92 ;
      RECT 0.165 0.23 0.325 0.53 ;
      RECT 0.375 1.17 0.795 1.27 ;
      RECT 0.165 0.63 0.925 0.73 ;
      RECT 0.875 1.62 1.035 1.92 ;
      RECT 0.875 0.23 1.035 0.53 ;
      RECT 0.165 1.42 1.135 1.52 ;
      RECT 1.115 1.175 1.595 1.275 ;
      RECT 1.575 1.62 1.735 1.92 ;
      RECT 1.575 0.23 1.735 0.53 ;
      RECT 0.285 0.945 1.975 1.045 ;
      RECT 0.795 0.93 1.125 1.06 ;
      RECT 1.825 1.62 1.985 1.92 ;
      RECT 1.825 0.23 1.985 0.53 ;
      RECT 2.305 1.62 2.465 1.92 ;
      RECT 2.305 0.23 2.465 0.53 ;
      RECT 1.215 0.63 2.18 0.73 ;
      RECT 2.08 0.63 2.18 0.975 ;
      RECT 2.08 0.875 2.835 0.975 ;
      RECT 2.305 0.63 3.065 0.73 ;
      RECT 3.015 1.62 3.175 1.92 ;
      RECT 3.015 0.23 3.175 0.53 ;
      RECT 1.965 1.15 3.265 1.25 ;
      RECT 2.935 1.135 3.265 1.265 ;
      RECT 2.305 1.42 3.285 1.52 ;
      RECT 3.39 1.42 3.81 1.52 ;
      RECT 3.725 0.23 3.885 0.53 ;
      RECT 3.625 0.915 4.045 1.015 ;
      RECT 3.915 1.62 4.075 1.92 ;
      RECT 4.285 1.62 4.445 1.92 ;
      RECT 3.915 1.325 4.535 1.425 ;
      RECT 4.475 0.23 4.635 0.53 ;
      RECT 4.375 1.085 4.795 1.185 ;
      RECT 3.375 0.63 4.875 0.73 ;
      RECT 4.285 0.835 5.005 0.925 ;
      RECT 4.285 0.83 4.445 0.93 ;
      RECT 4.975 0.23 5.135 0.53 ;
      RECT 4.995 1.62 5.155 1.92 ;
      RECT 0.46 1.62 0.55 2.52 ;
      RECT 1.36 1.62 1.45 2.52 ;
      RECT 2.11 1.62 2.2 2.52 ;
      RECT 2.6 1.62 2.69 2.52 ;
      RECT 3.5 1.62 3.59 2.52 ;
      RECT 4.77 1.62 4.86 2.52 ;
      RECT 0 2.3 5.32 2.52 ;
      RECT 0 -0.22 5.32 0 ;
      RECT 0.46 -0.22 0.55 0.53 ;
      RECT 1.36 -0.22 1.45 0.53 ;
      RECT 2.11 -0.22 2.2 0.53 ;
      RECT 2.6 -0.22 2.69 0.53 ;
      RECT 3.5 -0.22 3.59 0.53 ;
      RECT 4.02 -0.22 4.11 0.53 ;
      RECT 4.25 -0.22 4.34 0.53 ;
      RECT 4.77 -0.22 4.86 0.53 ;
    LAYER VI1 ;
      RECT 0.195 1.72 0.295 1.82 ;
      RECT 0.195 1.42 0.295 1.52 ;
      RECT 0.195 0.63 0.295 0.73 ;
      RECT 0.195 0.4 0.295 0.5 ;
      RECT 0.905 1.72 1.005 1.82 ;
      RECT 0.905 0.4 1.005 0.5 ;
      RECT 1.145 1.175 1.245 1.275 ;
      RECT 1.615 1.72 1.715 1.82 ;
      RECT 1.615 0.63 1.715 0.73 ;
      RECT 1.615 0.4 1.715 0.5 ;
      RECT 1.845 1.72 1.945 1.82 ;
      RECT 1.845 0.945 1.945 1.045 ;
      RECT 1.845 0.4 1.945 0.5 ;
      RECT 2.335 1.72 2.435 1.82 ;
      RECT 2.335 1.42 2.435 1.52 ;
      RECT 2.335 0.63 2.435 0.73 ;
      RECT 2.335 0.4 2.435 0.5 ;
      RECT 3.045 1.72 3.145 1.82 ;
      RECT 3.045 0.4 3.145 0.5 ;
      RECT 3.42 1.42 3.52 1.52 ;
      RECT 3.755 0.4 3.855 0.5 ;
      RECT 3.945 1.72 4.045 1.82 ;
      RECT 3.945 1.325 4.045 1.425 ;
      RECT 4.315 1.72 4.415 1.82 ;
      RECT 4.315 0.83 4.415 0.93 ;
      RECT 4.505 0.4 4.605 0.5 ;
      RECT 4.745 0.63 4.845 0.73 ;
      RECT 5.025 1.72 5.125 1.82 ;
      RECT 5.025 0.4 5.125 0.5 ;
    LAYER ME2 ;
      RECT 0.195 0.37 0.295 1.92 ;
      RECT 0.905 1.175 1.275 1.275 ;
      RECT 0.905 0.37 1.005 1.92 ;
      RECT 1.615 0.37 1.715 1.92 ;
      RECT 1.845 0.37 1.945 1.92 ;
      RECT 2.335 0.37 2.435 1.92 ;
      RECT 3.045 1.42 3.55 1.52 ;
      RECT 3.045 0.37 3.145 1.92 ;
      RECT 3.755 0.37 3.855 0.53 ;
      RECT 3.755 0.43 4.045 0.53 ;
      RECT 3.945 0.43 4.045 1.92 ;
      RECT 4.505 0.37 4.605 0.53 ;
      RECT 4.315 0.43 4.605 0.53 ;
      RECT 4.315 0.43 4.415 1.92 ;
      RECT 4.715 0.63 5.125 0.73 ;
      RECT 5.025 0.23 5.125 1.92 ;
  END
END QDFFNCSRX1

MACRO QDFFNCX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDFFNCX1 0 -0.11 ;
  SIZE 4.2 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.235 1.62 0.325 2.52 ;
        RECT 1.025 1.62 1.115 2.52 ;
        RECT 1.925 1.62 2.015 2.52 ;
        RECT 2.715 1.62 2.805 2.52 ;
        RECT 3.615 1.62 3.705 2.52 ;
        RECT 0 2.3 4.2 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.235 -0.22 0.325 0.53 ;
        RECT 1.025 -0.22 1.115 0.53 ;
        RECT 1.925 -0.22 2.015 0.53 ;
        RECT 2.715 -0.22 2.805 0.53 ;
        RECT 3.615 -0.22 3.705 0.53 ;
        RECT 0 -0.22 4.2 0 ;
    END
  END gnd!
  PIN CLKB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.23 0.83 2.31 0.93 ;
        RECT 1.845 0.915 3.39 1.015 ;
    END
  END CLKB
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 3.87 1.72 3.97 1.82 ;
        RECT 3.87 0.63 3.97 0.73 ;
        RECT 3.87 0.4 3.97 0.5 ;
      LAYER ME1 ;
        RECT 3.84 0.23 4 0.53 ;
        RECT 3.47 0.63 4 0.73 ;
        RECT 3.84 1.62 4 1.92 ;
      LAYER ME2 ;
        RECT 3.87 0.37 3.97 1.92 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.23 1.225 1.26 1.325 ;
    END
  END D
  OBS
    LAYER ME1 ;
      RECT 0.46 1.62 0.62 1.92 ;
      RECT 0.46 0.23 0.62 0.53 ;
      RECT 0.73 1.62 0.89 1.92 ;
      RECT 0.73 0.23 0.89 0.53 ;
      RECT 0.23 1.225 1.26 1.325 ;
      RECT 0.72 0.635 1.49 0.725 ;
      RECT 0.72 0.63 1.48 0.73 ;
      RECT 1.44 1.62 1.6 1.92 ;
      RECT 1.44 0.23 1.6 0.53 ;
      RECT 0.46 1.025 1.7 1.125 ;
      RECT 0.73 1.425 1.71 1.525 ;
      RECT 1.835 1.425 2.295 1.525 ;
      RECT 2.15 1.62 2.31 1.92 ;
      RECT 2.15 0.23 2.31 0.53 ;
      RECT 1.78 0.63 2.32 0.73 ;
      RECT 2.42 1.62 2.58 1.92 ;
      RECT 2.42 0.23 2.58 0.53 ;
      RECT 2.15 1.135 2.95 1.225 ;
      RECT 2.15 1.13 2.93 1.23 ;
      RECT 2.42 0.63 3.18 0.73 ;
      RECT 3.13 1.62 3.29 1.92 ;
      RECT 3.13 0.23 3.29 0.53 ;
      RECT 0.23 0.83 2.31 0.93 ;
      RECT 1.845 0.915 3.39 1.015 ;
      RECT 2.42 1.425 3.4 1.525 ;
      RECT 3.36 1.12 3.85 1.22 ;
      RECT 3.84 1.62 4 1.92 ;
      RECT 3.47 0.63 4 0.73 ;
      RECT 3.84 0.23 4 0.53 ;
      RECT 0.235 1.62 0.325 2.52 ;
      RECT 1.025 1.62 1.115 2.52 ;
      RECT 1.925 1.62 2.015 2.52 ;
      RECT 2.715 1.62 2.805 2.52 ;
      RECT 3.615 1.62 3.705 2.52 ;
      RECT 0 2.3 4.2 2.52 ;
      RECT 0 -0.22 4.2 0 ;
      RECT 0.235 -0.22 0.325 0.53 ;
      RECT 1.025 -0.22 1.115 0.53 ;
      RECT 1.925 -0.22 2.015 0.53 ;
      RECT 2.715 -0.22 2.805 0.53 ;
      RECT 3.615 -0.22 3.705 0.53 ;
    LAYER VI1 ;
      RECT 0.49 1.72 0.59 1.82 ;
      RECT 0.49 1.025 0.59 1.125 ;
      RECT 0.49 0.4 0.59 0.5 ;
      RECT 0.76 1.72 0.86 1.82 ;
      RECT 0.76 1.425 0.86 1.525 ;
      RECT 0.76 0.63 0.86 0.73 ;
      RECT 0.76 0.4 0.86 0.5 ;
      RECT 1.47 1.72 1.57 1.82 ;
      RECT 1.47 0.4 1.57 0.5 ;
      RECT 1.9 1.425 2 1.525 ;
      RECT 2.18 1.72 2.28 1.82 ;
      RECT 2.18 1.13 2.28 1.23 ;
      RECT 2.18 0.63 2.28 0.73 ;
      RECT 2.18 0.4 2.28 0.5 ;
      RECT 2.45 1.72 2.55 1.82 ;
      RECT 2.45 1.425 2.55 1.525 ;
      RECT 2.45 0.63 2.55 0.73 ;
      RECT 2.45 0.4 2.55 0.5 ;
      RECT 3.16 1.72 3.26 1.82 ;
      RECT 3.16 0.4 3.26 0.5 ;
      RECT 3.4 1.12 3.5 1.22 ;
      RECT 3.87 1.72 3.97 1.82 ;
      RECT 3.87 0.63 3.97 0.73 ;
      RECT 3.87 0.4 3.97 0.5 ;
    LAYER ME2 ;
      RECT 0.49 0.37 0.59 1.92 ;
      RECT 0.76 0.63 1.36 0.73 ;
      RECT 0.76 0.37 0.86 1.92 ;
      RECT 1.47 1.425 2.03 1.525 ;
      RECT 1.47 0.37 1.57 1.92 ;
      RECT 2.18 0.37 2.28 1.92 ;
      RECT 2.45 0.37 2.55 1.92 ;
      RECT 3.16 1.12 3.53 1.22 ;
      RECT 3.16 0.37 3.26 1.92 ;
      RECT 3.87 0.37 3.97 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDFFNCX1

MACRO QDLATENSX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDLATENSX1 0 -0.11 ;
  SIZE 2.24 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.31 1.13 0.73 1.23 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.29 0.915 1.16 1.015 ;
        RECT 0.83 0.9 1.16 1.03 ;
    END
  END G
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.52 0.915 1.94 1.015 ;
    END
  END SETB
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.495 -0.22 0.585 0.53 ;
        RECT 1.395 -0.22 1.485 0.53 ;
        RECT 0 -0.22 2.24 0 ;
    END
  END gnd!
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.56 0.63 1.66 0.73 ;
        RECT 1.65 1.72 1.75 1.82 ;
        RECT 1.84 0.4 1.94 0.5 ;
      LAYER ME1 ;
        RECT 1.81 0.23 1.97 0.53 ;
        RECT 1.62 1.62 1.78 1.92 ;
        RECT 1.27 0.63 1.77 0.73 ;
      LAYER ME2 ;
        RECT 1.65 1.62 1.94 1.72 ;
        RECT 1.84 0.37 1.94 1.72 ;
        RECT 1.53 0.63 1.94 0.73 ;
        RECT 1.65 1.62 1.75 1.92 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.495 1.62 0.585 2.52 ;
        RECT 1.395 1.62 1.485 2.52 ;
        RECT 1.915 1.62 2.005 2.52 ;
        RECT 0 2.3 2.24 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.2 1.62 0.36 1.92 ;
      RECT 0.2 0.23 0.36 0.53 ;
      RECT 0.31 1.13 0.73 1.23 ;
      RECT 0.58 1.42 1.05 1.52 ;
      RECT 0.91 1.62 1.07 1.92 ;
      RECT 0.91 0.23 1.07 0.53 ;
      RECT 0.29 0.915 1.16 1.015 ;
      RECT 0.83 0.9 1.16 1.03 ;
      RECT 0.67 0.63 1.17 0.73 ;
      RECT 1.15 1.42 1.63 1.52 ;
      RECT 1.27 0.63 1.77 0.73 ;
      RECT 1.62 1.62 1.78 1.92 ;
      RECT 1.52 0.915 1.94 1.015 ;
      RECT 1.81 0.23 1.97 0.53 ;
      RECT 0.495 1.62 0.585 2.52 ;
      RECT 1.395 1.62 1.485 2.52 ;
      RECT 1.915 1.62 2.005 2.52 ;
      RECT 0 2.3 2.24 2.52 ;
      RECT 0 -0.22 2.24 0 ;
      RECT 0.495 -0.22 0.585 0.53 ;
      RECT 1.395 -0.22 1.485 0.53 ;
    LAYER VI1 ;
      RECT 0.23 1.72 0.33 1.82 ;
      RECT 0.23 0.4 0.33 0.5 ;
      RECT 0.7 1.42 0.8 1.52 ;
      RECT 0.7 0.63 0.8 0.73 ;
      RECT 0.94 1.72 1.04 1.82 ;
      RECT 0.94 0.4 1.04 0.5 ;
      RECT 1.18 1.42 1.28 1.52 ;
      RECT 1.56 0.63 1.66 0.73 ;
      RECT 1.65 1.72 1.75 1.82 ;
      RECT 1.84 0.4 1.94 0.5 ;
    LAYER ME2 ;
      RECT 0.23 0.63 0.83 0.73 ;
      RECT 0.23 1.42 0.83 1.52 ;
      RECT 0.23 0.37 0.33 1.92 ;
      RECT 0.94 1.42 1.31 1.52 ;
      RECT 0.94 0.37 1.04 1.92 ;
      RECT 1.53 0.63 1.94 0.73 ;
      RECT 1.84 0.37 1.94 1.72 ;
      RECT 1.65 1.62 1.94 1.72 ;
      RECT 1.65 1.62 1.75 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDLATENSX1

MACRO QDLATERX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDLATERX1 0 -0.11 ;
  SIZE 2.24 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.31 1.13 0.73 1.23 ;
    END
  END D
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.52 0.915 1.94 1.015 ;
    END
  END RST
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.495 -0.22 0.585 0.53 ;
        RECT 1.395 -0.22 1.485 0.53 ;
        RECT 1.915 -0.22 2.005 0.53 ;
        RECT 0 -0.22 2.24 0 ;
    END
  END gnd!
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.56 0.63 1.66 0.73 ;
        RECT 1.65 0.4 1.75 0.5 ;
        RECT 1.84 1.72 1.94 1.82 ;
      LAYER ME1 ;
        RECT 1.81 1.62 1.97 1.92 ;
        RECT 1.62 0.23 1.78 0.53 ;
        RECT 1.27 0.63 1.77 0.73 ;
      LAYER ME2 ;
        RECT 1.84 0.43 1.94 1.92 ;
        RECT 1.53 0.63 1.94 0.73 ;
        RECT 1.65 0.43 1.94 0.53 ;
        RECT 1.65 0.37 1.75 0.53 ;
    END
  END Q
  PIN G
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.29 0.915 1.16 1.015 ;
        RECT 0.83 0.9 1.16 1.03 ;
    END
  END G
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.495 1.62 0.585 2.52 ;
        RECT 1.395 1.62 1.485 2.52 ;
        RECT 0 2.3 2.24 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.2 1.62 0.36 1.92 ;
      RECT 0.2 0.23 0.36 0.53 ;
      RECT 0.31 1.13 0.73 1.23 ;
      RECT 0.58 1.42 1.05 1.52 ;
      RECT 0.91 1.62 1.07 1.92 ;
      RECT 0.91 0.23 1.07 0.53 ;
      RECT 0.29 0.915 1.16 1.015 ;
      RECT 0.83 0.9 1.16 1.03 ;
      RECT 0.67 0.63 1.17 0.73 ;
      RECT 1.15 1.42 1.63 1.52 ;
      RECT 1.27 0.63 1.77 0.73 ;
      RECT 1.62 0.23 1.78 0.53 ;
      RECT 1.52 0.915 1.94 1.015 ;
      RECT 1.81 1.62 1.97 1.92 ;
      RECT 0.495 1.62 0.585 2.52 ;
      RECT 1.395 1.62 1.485 2.52 ;
      RECT 0 2.3 2.24 2.52 ;
      RECT 0 -0.22 2.24 0 ;
      RECT 0.495 -0.22 0.585 0.53 ;
      RECT 1.395 -0.22 1.485 0.53 ;
      RECT 1.915 -0.22 2.005 0.53 ;
    LAYER VI1 ;
      RECT 0.23 1.72 0.33 1.82 ;
      RECT 0.23 0.4 0.33 0.5 ;
      RECT 0.7 1.42 0.8 1.52 ;
      RECT 0.7 0.63 0.8 0.73 ;
      RECT 0.94 1.72 1.04 1.82 ;
      RECT 0.94 0.4 1.04 0.5 ;
      RECT 1.18 1.42 1.28 1.52 ;
      RECT 1.56 0.63 1.66 0.73 ;
      RECT 1.65 0.4 1.75 0.5 ;
      RECT 1.84 1.72 1.94 1.82 ;
    LAYER ME2 ;
      RECT 0.23 0.63 0.83 0.73 ;
      RECT 0.23 1.42 0.83 1.52 ;
      RECT 0.23 0.37 0.33 1.92 ;
      RECT 0.94 1.42 1.31 1.52 ;
      RECT 0.94 0.37 1.04 1.92 ;
      RECT 1.65 0.37 1.75 0.53 ;
      RECT 1.65 0.43 1.94 0.53 ;
      RECT 1.53 0.63 1.94 0.73 ;
      RECT 1.84 0.43 1.94 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDLATERX1

MACRO QDLATESRX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDLATESRX1 0 -0.11 ;
  SIZE 3.08 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.225 1.13 0.645 1.23 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.205 0.915 1.075 1.015 ;
        RECT 0.745 0.9 1.075 1.03 ;
    END
  END G
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.435 0.915 1.855 1.015 ;
    END
  END RST
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.41 -0.22 0.5 0.53 ;
        RECT 1.31 -0.22 1.4 0.53 ;
        RECT 1.83 -0.22 1.92 0.53 ;
        RECT 2.06 -0.22 2.15 0.53 ;
        RECT 2.58 -0.22 2.67 0.53 ;
        RECT 0 -0.22 3.08 0 ;
    END
  END gnd!
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 2.555 0.63 2.655 0.73 ;
        RECT 2.835 1.72 2.935 1.82 ;
        RECT 2.835 0.4 2.935 0.5 ;
      LAYER ME1 ;
        RECT 2.805 1.62 2.965 1.92 ;
        RECT 2.785 0.23 2.945 0.53 ;
        RECT 1.185 0.63 2.685 0.73 ;
      LAYER ME2 ;
        RECT 2.835 0.23 2.935 1.92 ;
        RECT 2.525 0.63 2.935 0.73 ;
    END
  END Q
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 2.185 1.085 2.605 1.185 ;
    END
  END SET
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.41 1.62 0.5 2.52 ;
        RECT 1.31 1.62 1.4 2.52 ;
        RECT 2.58 1.62 2.67 2.52 ;
        RECT 0 2.3 3.08 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.115 1.62 0.275 1.92 ;
      RECT 0.115 0.23 0.275 0.53 ;
      RECT 0.225 1.13 0.645 1.23 ;
      RECT 0.495 1.42 0.965 1.52 ;
      RECT 0.825 1.62 0.985 1.92 ;
      RECT 0.825 0.23 0.985 0.53 ;
      RECT 0.205 0.915 1.075 1.015 ;
      RECT 0.745 0.9 1.075 1.03 ;
      RECT 0.585 0.63 1.085 0.73 ;
      RECT 1.065 1.42 1.545 1.52 ;
      RECT 1.535 0.23 1.695 0.53 ;
      RECT 1.435 0.915 1.855 1.015 ;
      RECT 1.725 1.62 1.885 1.92 ;
      RECT 2.095 1.62 2.255 1.92 ;
      RECT 1.725 1.325 2.345 1.425 ;
      RECT 2.285 0.23 2.445 0.53 ;
      RECT 2.185 1.085 2.605 1.185 ;
      RECT 1.185 0.63 2.685 0.73 ;
      RECT 2.095 0.835 2.815 0.925 ;
      RECT 2.095 0.83 2.255 0.93 ;
      RECT 2.785 0.23 2.945 0.53 ;
      RECT 2.805 1.62 2.965 1.92 ;
      RECT 0.41 1.62 0.5 2.52 ;
      RECT 1.31 1.62 1.4 2.52 ;
      RECT 2.58 1.62 2.67 2.52 ;
      RECT 0 2.3 3.08 2.52 ;
      RECT 0 -0.22 3.08 0 ;
      RECT 0.41 -0.22 0.5 0.53 ;
      RECT 1.31 -0.22 1.4 0.53 ;
      RECT 1.83 -0.22 1.92 0.53 ;
      RECT 2.06 -0.22 2.15 0.53 ;
      RECT 2.58 -0.22 2.67 0.53 ;
    LAYER VI1 ;
      RECT 0.145 1.72 0.245 1.82 ;
      RECT 0.145 0.4 0.245 0.5 ;
      RECT 0.615 1.42 0.715 1.52 ;
      RECT 0.615 0.63 0.715 0.73 ;
      RECT 0.855 1.72 0.955 1.82 ;
      RECT 0.855 0.4 0.955 0.5 ;
      RECT 1.095 1.42 1.195 1.52 ;
      RECT 1.565 0.4 1.665 0.5 ;
      RECT 1.755 1.72 1.855 1.82 ;
      RECT 1.755 1.325 1.855 1.425 ;
      RECT 2.125 1.72 2.225 1.82 ;
      RECT 2.125 0.83 2.225 0.93 ;
      RECT 2.315 0.4 2.415 0.5 ;
      RECT 2.555 0.63 2.655 0.73 ;
      RECT 2.835 1.72 2.935 1.82 ;
      RECT 2.835 0.4 2.935 0.5 ;
    LAYER ME2 ;
      RECT 0.145 0.63 0.745 0.73 ;
      RECT 0.145 1.42 0.745 1.52 ;
      RECT 0.145 0.37 0.245 1.92 ;
      RECT 0.855 1.42 1.225 1.52 ;
      RECT 0.855 0.37 0.955 1.92 ;
      RECT 1.565 0.37 1.665 0.53 ;
      RECT 1.565 0.43 1.855 0.53 ;
      RECT 1.755 0.43 1.855 1.92 ;
      RECT 2.315 0.37 2.415 0.53 ;
      RECT 2.125 0.43 2.415 0.53 ;
      RECT 2.125 0.43 2.225 1.92 ;
      RECT 2.525 0.63 2.935 0.73 ;
      RECT 2.835 0.23 2.935 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDLATESRX1

MACRO QDLATEX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDLATEX1 0 -0.11 ;
  SIZE 1.96 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.3 0.83 0.72 0.93 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.31 1.045 1.15 1.145 ;
        RECT 0.82 1.03 1.15 1.16 ;
    END
  END G
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 -0.22 0.575 0.53 ;
        RECT 1.385 -0.22 1.475 0.53 ;
        RECT 0 -0.22 1.96 0 ;
    END
  END gnd!
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.64 1.72 1.74 1.82 ;
        RECT 1.64 0.63 1.74 0.73 ;
        RECT 1.64 0.4 1.74 0.5 ;
      LAYER ME1 ;
        RECT 1.61 0.23 1.77 0.53 ;
        RECT 1.25 0.63 1.77 0.73 ;
        RECT 1.61 1.62 1.77 1.92 ;
      LAYER ME2 ;
        RECT 1.64 0.23 1.74 1.92 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 1.62 0.575 2.52 ;
        RECT 1.385 1.62 1.475 2.52 ;
        RECT 0 2.3 1.96 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.19 1.62 0.35 1.92 ;
      RECT 0.19 0.23 0.35 0.53 ;
      RECT 0.3 0.83 0.72 0.93 ;
      RECT 0.57 1.42 1.04 1.52 ;
      RECT 0.9 1.62 1.06 1.92 ;
      RECT 0.9 0.23 1.06 0.53 ;
      RECT 0.31 1.045 1.15 1.145 ;
      RECT 0.82 1.03 1.15 1.16 ;
      RECT 0.66 0.63 1.16 0.73 ;
      RECT 1.14 1.42 1.62 1.52 ;
      RECT 1.61 1.62 1.77 1.92 ;
      RECT 1.25 0.63 1.77 0.73 ;
      RECT 1.61 0.23 1.77 0.53 ;
      RECT 0.485 1.62 0.575 2.52 ;
      RECT 1.385 1.62 1.475 2.52 ;
      RECT 0 2.3 1.96 2.52 ;
      RECT 0 -0.22 1.96 0 ;
      RECT 0.485 -0.22 0.575 0.53 ;
      RECT 1.385 -0.22 1.475 0.53 ;
    LAYER VI1 ;
      RECT 0.22 1.72 0.32 1.82 ;
      RECT 0.22 0.4 0.32 0.5 ;
      RECT 0.69 1.42 0.79 1.52 ;
      RECT 0.69 0.63 0.79 0.73 ;
      RECT 0.93 1.72 1.03 1.82 ;
      RECT 0.93 0.4 1.03 0.5 ;
      RECT 1.17 1.42 1.27 1.52 ;
      RECT 1.64 1.72 1.74 1.82 ;
      RECT 1.64 0.63 1.74 0.73 ;
      RECT 1.64 0.4 1.74 0.5 ;
    LAYER ME2 ;
      RECT 0.22 0.63 0.82 0.73 ;
      RECT 0.22 1.42 0.82 1.52 ;
      RECT 0.22 0.37 0.32 1.92 ;
      RECT 0.93 1.42 1.3 1.52 ;
      RECT 0.93 0.37 1.03 1.92 ;
      RECT 1.64 0.23 1.74 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDLATEX1

MACRO QDLATNENSX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDLATNENSX1 0 -0.11 ;
  SIZE 2.24 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.31 0.83 0.73 0.93 ;
    END
  END D
  PIN GB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.29 1.045 1.16 1.145 ;
        RECT 0.83 1.03 1.16 1.16 ;
    END
  END GB
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.52 1.42 1.94 1.52 ;
    END
  END SETB
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.495 -0.22 0.585 0.53 ;
        RECT 1.395 -0.22 1.485 0.53 ;
        RECT 0 -0.22 2.24 0 ;
    END
  END gnd!
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.56 0.63 1.66 0.73 ;
        RECT 1.65 1.72 1.75 1.82 ;
        RECT 1.84 0.4 1.94 0.5 ;
      LAYER ME1 ;
        RECT 1.81 0.23 1.97 0.53 ;
        RECT 1.62 1.62 1.78 1.92 ;
        RECT 1.22 0.63 1.69 0.73 ;
      LAYER ME2 ;
        RECT 1.65 1.62 1.94 1.72 ;
        RECT 1.84 0.37 1.94 1.72 ;
        RECT 1.53 0.63 1.94 0.73 ;
        RECT 1.65 1.62 1.75 1.92 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.495 1.62 0.585 2.52 ;
        RECT 1.395 1.62 1.485 2.52 ;
        RECT 1.915 1.62 2.005 2.52 ;
        RECT 0 2.3 2.24 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.2 1.62 0.36 1.92 ;
      RECT 0.2 0.23 0.36 0.53 ;
      RECT 0.31 0.83 0.73 0.93 ;
      RECT 0.2 0.63 0.96 0.73 ;
      RECT 0.91 1.62 1.07 1.92 ;
      RECT 0.91 0.23 1.07 0.53 ;
      RECT 0.29 1.045 1.16 1.145 ;
      RECT 0.83 1.03 1.16 1.16 ;
      RECT 0.2 1.42 1.18 1.52 ;
      RECT 1.15 0.83 1.63 0.93 ;
      RECT 1.22 0.63 1.69 0.73 ;
      RECT 1.62 1.62 1.78 1.92 ;
      RECT 1.52 1.42 1.94 1.52 ;
      RECT 1.81 0.23 1.97 0.53 ;
      RECT 0.495 1.62 0.585 2.52 ;
      RECT 1.395 1.62 1.485 2.52 ;
      RECT 1.915 1.62 2.005 2.52 ;
      RECT 0 2.3 2.24 2.52 ;
      RECT 0 -0.22 2.24 0 ;
      RECT 0.495 -0.22 0.585 0.53 ;
      RECT 1.395 -0.22 1.485 0.53 ;
    LAYER VI1 ;
      RECT 0.23 1.72 0.33 1.82 ;
      RECT 0.23 1.42 0.33 1.52 ;
      RECT 0.23 0.63 0.33 0.73 ;
      RECT 0.23 0.4 0.33 0.5 ;
      RECT 0.94 1.72 1.04 1.82 ;
      RECT 0.94 0.4 1.04 0.5 ;
      RECT 1.18 0.83 1.28 0.93 ;
      RECT 1.56 0.63 1.66 0.73 ;
      RECT 1.65 1.72 1.75 1.82 ;
      RECT 1.84 0.4 1.94 0.5 ;
    LAYER ME2 ;
      RECT 0.23 0.37 0.33 1.92 ;
      RECT 0.94 0.83 1.31 0.93 ;
      RECT 0.94 0.37 1.04 1.92 ;
      RECT 1.53 0.63 1.94 0.73 ;
      RECT 1.84 0.37 1.94 1.72 ;
      RECT 1.65 1.62 1.94 1.72 ;
      RECT 1.65 1.62 1.75 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDLATNENSX1

MACRO QDLATNERX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDLATNERX1 0 -0.11 ;
  SIZE 2.24 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.31 0.83 0.73 0.93 ;
    END
  END D
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.48 1.42 1.9 1.52 ;
    END
  END RST
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.495 -0.22 0.585 0.53 ;
        RECT 1.395 -0.22 1.485 0.53 ;
        RECT 1.915 -0.22 2.005 0.53 ;
        RECT 0 -0.22 2.24 0 ;
    END
  END gnd!
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.56 0.63 1.66 0.73 ;
        RECT 1.65 0.4 1.75 0.5 ;
        RECT 1.84 1.72 1.94 1.82 ;
      LAYER ME1 ;
        RECT 1.81 1.62 1.97 1.92 ;
        RECT 1.62 0.23 1.78 0.53 ;
        RECT 1.22 0.63 1.69 0.73 ;
      LAYER ME2 ;
        RECT 1.84 0.43 1.94 1.92 ;
        RECT 1.53 0.63 1.94 0.73 ;
        RECT 1.65 0.43 1.94 0.53 ;
        RECT 1.65 0.37 1.75 0.53 ;
    END
  END Q
  PIN GB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.29 1.045 1.16 1.145 ;
        RECT 0.83 1.03 1.16 1.16 ;
    END
  END GB
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.495 1.62 0.585 2.52 ;
        RECT 1.395 1.62 1.485 2.52 ;
        RECT 0 2.3 2.24 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.2 1.62 0.36 1.92 ;
      RECT 0.2 0.23 0.36 0.53 ;
      RECT 0.31 0.83 0.73 0.93 ;
      RECT 0.2 0.63 0.96 0.73 ;
      RECT 0.91 1.62 1.07 1.92 ;
      RECT 0.91 0.23 1.07 0.53 ;
      RECT 0.29 1.045 1.16 1.145 ;
      RECT 0.83 1.03 1.16 1.16 ;
      RECT 0.2 1.42 1.18 1.52 ;
      RECT 1.15 0.83 1.63 0.93 ;
      RECT 1.22 0.63 1.69 0.73 ;
      RECT 1.62 0.23 1.78 0.53 ;
      RECT 1.48 1.42 1.9 1.52 ;
      RECT 1.81 1.62 1.97 1.92 ;
      RECT 0.495 1.62 0.585 2.52 ;
      RECT 1.395 1.62 1.485 2.52 ;
      RECT 0 2.3 2.24 2.52 ;
      RECT 0 -0.22 2.24 0 ;
      RECT 0.495 -0.22 0.585 0.53 ;
      RECT 1.395 -0.22 1.485 0.53 ;
      RECT 1.915 -0.22 2.005 0.53 ;
    LAYER VI1 ;
      RECT 0.23 1.72 0.33 1.82 ;
      RECT 0.23 1.42 0.33 1.52 ;
      RECT 0.23 0.63 0.33 0.73 ;
      RECT 0.23 0.4 0.33 0.5 ;
      RECT 0.94 1.72 1.04 1.82 ;
      RECT 0.94 0.4 1.04 0.5 ;
      RECT 1.18 0.83 1.28 0.93 ;
      RECT 1.56 0.63 1.66 0.73 ;
      RECT 1.65 0.4 1.75 0.5 ;
      RECT 1.84 1.72 1.94 1.82 ;
    LAYER ME2 ;
      RECT 0.23 0.37 0.33 1.92 ;
      RECT 0.94 0.83 1.31 0.93 ;
      RECT 0.94 0.37 1.04 1.92 ;
      RECT 1.65 0.37 1.75 0.53 ;
      RECT 1.65 0.43 1.94 0.53 ;
      RECT 1.53 0.63 1.94 0.73 ;
      RECT 1.84 0.43 1.94 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDLATNERX1

MACRO QDLATNESRX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDLATNESRX1 0 -0.11 ;
  SIZE 3.08 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.225 1.13 0.645 1.23 ;
    END
  END D
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 1.435 0.915 1.855 1.015 ;
    END
  END RST
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.41 -0.22 0.5 0.53 ;
        RECT 1.31 -0.22 1.4 0.53 ;
        RECT 1.83 -0.22 1.92 0.53 ;
        RECT 2.06 -0.22 2.15 0.53 ;
        RECT 2.58 -0.22 2.67 0.53 ;
        RECT 0 -0.22 3.08 0 ;
    END
  END gnd!
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 2.555 0.63 2.655 0.73 ;
        RECT 2.835 1.72 2.935 1.82 ;
        RECT 2.835 0.4 2.935 0.5 ;
      LAYER ME1 ;
        RECT 2.805 1.62 2.965 1.92 ;
        RECT 2.785 0.23 2.945 0.53 ;
        RECT 1.185 0.63 2.685 0.73 ;
      LAYER ME2 ;
        RECT 2.835 0.23 2.935 1.92 ;
        RECT 2.525 0.63 2.935 0.73 ;
    END
  END Q
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 2.185 1.085 2.605 1.185 ;
    END
  END SET
  PIN GB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.205 0.915 1.075 1.015 ;
        RECT 0.745 0.9 1.075 1.03 ;
    END
  END GB
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.41 1.62 0.5 2.52 ;
        RECT 1.31 1.62 1.4 2.52 ;
        RECT 2.58 1.62 2.67 2.52 ;
        RECT 0 2.3 3.08 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.115 1.62 0.275 1.92 ;
      RECT 0.115 0.23 0.275 0.53 ;
      RECT 0.225 1.13 0.645 1.23 ;
      RECT 0.115 0.63 0.875 0.73 ;
      RECT 0.825 1.62 0.985 1.92 ;
      RECT 0.825 0.23 0.985 0.53 ;
      RECT 0.205 0.915 1.075 1.015 ;
      RECT 0.745 0.9 1.075 1.03 ;
      RECT 0.115 1.42 1.095 1.52 ;
      RECT 1.2 1.42 1.62 1.52 ;
      RECT 1.535 0.23 1.695 0.53 ;
      RECT 1.435 0.915 1.855 1.015 ;
      RECT 1.725 1.62 1.885 1.92 ;
      RECT 2.095 1.62 2.255 1.92 ;
      RECT 1.725 1.325 2.345 1.425 ;
      RECT 2.285 0.23 2.445 0.53 ;
      RECT 2.185 1.085 2.605 1.185 ;
      RECT 1.185 0.63 2.685 0.73 ;
      RECT 2.095 0.835 2.815 0.925 ;
      RECT 2.095 0.83 2.255 0.93 ;
      RECT 2.785 0.23 2.945 0.53 ;
      RECT 2.805 1.62 2.965 1.92 ;
      RECT 0.41 1.62 0.5 2.52 ;
      RECT 1.31 1.62 1.4 2.52 ;
      RECT 2.58 1.62 2.67 2.52 ;
      RECT 0 2.3 3.08 2.52 ;
      RECT 0 -0.22 3.08 0 ;
      RECT 0.41 -0.22 0.5 0.53 ;
      RECT 1.31 -0.22 1.4 0.53 ;
      RECT 1.83 -0.22 1.92 0.53 ;
      RECT 2.06 -0.22 2.15 0.53 ;
      RECT 2.58 -0.22 2.67 0.53 ;
    LAYER VI1 ;
      RECT 0.145 1.72 0.245 1.82 ;
      RECT 0.145 1.42 0.245 1.52 ;
      RECT 0.145 0.63 0.245 0.73 ;
      RECT 0.145 0.4 0.245 0.5 ;
      RECT 0.855 1.72 0.955 1.82 ;
      RECT 0.855 0.4 0.955 0.5 ;
      RECT 1.23 1.42 1.33 1.52 ;
      RECT 1.565 0.4 1.665 0.5 ;
      RECT 1.755 1.72 1.855 1.82 ;
      RECT 1.755 1.325 1.855 1.425 ;
      RECT 2.125 1.72 2.225 1.82 ;
      RECT 2.125 0.83 2.225 0.93 ;
      RECT 2.315 0.4 2.415 0.5 ;
      RECT 2.555 0.63 2.655 0.73 ;
      RECT 2.835 1.72 2.935 1.82 ;
      RECT 2.835 0.4 2.935 0.5 ;
    LAYER ME2 ;
      RECT 0.145 0.37 0.245 1.92 ;
      RECT 0.855 1.42 1.36 1.52 ;
      RECT 0.855 0.37 0.955 1.92 ;
      RECT 1.565 0.37 1.665 0.53 ;
      RECT 1.565 0.43 1.855 0.53 ;
      RECT 1.755 0.43 1.855 1.92 ;
      RECT 2.315 0.37 2.415 0.53 ;
      RECT 2.125 0.43 2.415 0.53 ;
      RECT 2.125 0.43 2.225 1.92 ;
      RECT 2.525 0.63 2.935 0.73 ;
      RECT 2.835 0.23 2.935 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDLATNESRX1

MACRO QDLATNEX1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN QDLATNEX1 0 -0.11 ;
  SIZE 1.96 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.3 0.83 0.72 0.93 ;
    END
  END D
  PIN GB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER ME1 ;
        RECT 0.31 1.045 1.15 1.145 ;
        RECT 0.82 1.03 1.15 1.16 ;
    END
  END GB
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 -0.22 0.575 0.53 ;
        RECT 1.385 -0.22 1.475 0.53 ;
        RECT 0 -0.22 1.96 0 ;
    END
  END gnd!
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.64 1.72 1.74 1.82 ;
        RECT 1.64 0.63 1.74 0.73 ;
        RECT 1.64 0.4 1.74 0.5 ;
      LAYER ME1 ;
        RECT 1.61 0.23 1.77 0.53 ;
        RECT 1.24 0.63 1.77 0.73 ;
        RECT 1.61 1.62 1.77 1.92 ;
      LAYER ME2 ;
        RECT 1.64 0.37 1.74 1.92 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 1.62 0.575 2.52 ;
        RECT 1.385 1.62 1.475 2.52 ;
        RECT 0 2.3 1.96 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.19 1.62 0.35 1.92 ;
      RECT 0.19 0.23 0.35 0.53 ;
      RECT 0.3 0.83 0.72 0.93 ;
      RECT 0.19 0.63 0.95 0.73 ;
      RECT 0.9 1.62 1.06 1.92 ;
      RECT 0.9 0.23 1.06 0.53 ;
      RECT 0.31 1.045 1.15 1.145 ;
      RECT 0.82 1.03 1.15 1.16 ;
      RECT 0.19 1.42 1.16 1.52 ;
      RECT 1.14 0.83 1.62 0.93 ;
      RECT 1.61 1.62 1.77 1.92 ;
      RECT 1.24 0.63 1.77 0.73 ;
      RECT 1.61 0.23 1.77 0.53 ;
      RECT 0.485 1.62 0.575 2.52 ;
      RECT 1.385 1.62 1.475 2.52 ;
      RECT 0 2.3 1.96 2.52 ;
      RECT 0 -0.22 1.96 0 ;
      RECT 0.485 -0.22 0.575 0.53 ;
      RECT 1.385 -0.22 1.475 0.53 ;
    LAYER VI1 ;
      RECT 0.22 1.72 0.32 1.82 ;
      RECT 0.22 1.42 0.32 1.52 ;
      RECT 0.22 0.63 0.32 0.73 ;
      RECT 0.22 0.4 0.32 0.5 ;
      RECT 0.93 1.72 1.03 1.82 ;
      RECT 0.93 0.4 1.03 0.5 ;
      RECT 1.17 0.83 1.27 0.93 ;
      RECT 1.64 1.72 1.74 1.82 ;
      RECT 1.64 0.63 1.74 0.73 ;
      RECT 1.64 0.4 1.74 0.5 ;
    LAYER ME2 ;
      RECT 0.22 0.37 0.32 1.92 ;
      RECT 0.93 0.83 1.3 0.93 ;
      RECT 0.93 0.37 1.03 1.92 ;
      RECT 1.64 0.37 1.74 1.92 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END QDLATNEX1

MACRO TIE0X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN TIE0X1 0 -0.11 ;
  SIZE 0.56 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.365 0.38 0.455 1.085 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 -0.22 0.195 0.53 ;
        RECT 0 -0.22 0.56 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 1.62 0.195 2.52 ;
        RECT 0 2.3 0.56 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.22 1.33 0.455 1.42 ;
      RECT 0.365 1.33 0.455 1.92 ;
      RECT 0.365 0.38 0.455 1.085 ;
      RECT 0.105 1.62 0.195 2.52 ;
      RECT 0 2.3 0.56 2.52 ;
      RECT 0 -0.22 0.56 0 ;
      RECT 0.105 -0.22 0.195 0.53 ;
  END
END TIE0X1

MACRO TIE0X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN TIE0X2 0 -0.11 ;
  SIZE 0.56 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.365 0.38 0.455 0.95 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 -0.22 0.195 0.68 ;
        RECT 0 -0.22 0.56 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 1.32 0.195 2.52 ;
        RECT 0 2.3 0.56 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.22 1.07 0.455 1.16 ;
      RECT 0.365 1.07 0.455 1.92 ;
      RECT 0.365 0.38 0.455 0.95 ;
      RECT 0.105 1.32 0.195 2.52 ;
      RECT 0 2.3 0.56 2.52 ;
      RECT 0 -0.22 0.56 0 ;
      RECT 0.105 -0.22 0.195 0.68 ;
  END
END TIE0X2

MACRO TIE0X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN TIE0X4 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 1.32 0.205 2.52 ;
        RECT 0.635 1.32 0.725 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.375 0.38 0.465 0.92 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 -0.22 0.205 0.68 ;
        RECT 0.635 -0.22 0.725 0.68 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.375 1.03 0.465 1.92 ;
      RECT 0.375 0.38 0.465 0.92 ;
      RECT 0.115 1.32 0.205 2.52 ;
      RECT 0.635 1.32 0.725 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.115 -0.22 0.205 0.68 ;
      RECT 0.635 -0.22 0.725 0.68 ;
  END
END TIE0X4

MACRO TIE1X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN TIE1X1 0 -0.11 ;
  SIZE 0.56 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.365 1.05 0.455 1.92 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 -0.22 0.195 0.53 ;
        RECT 0 -0.22 0.56 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 1.62 0.195 2.52 ;
        RECT 0 2.3 0.56 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.365 1.05 0.455 1.92 ;
      RECT 0.365 0.38 0.455 0.79 ;
      RECT 0.22 0.7 0.455 0.79 ;
      RECT 0.105 1.62 0.195 2.52 ;
      RECT 0 2.3 0.56 2.52 ;
      RECT 0 -0.22 0.56 0 ;
      RECT 0.105 -0.22 0.195 0.53 ;
  END
END TIE1X1

MACRO TIE1X2
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN TIE1X2 0 -0.11 ;
  SIZE 0.56 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.365 1.05 0.455 1.92 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 -0.22 0.195 0.68 ;
        RECT 0 -0.22 0.56 0 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.105 1.32 0.195 2.52 ;
        RECT 0 2.3 0.56 2.52 ;
    END
  END vdd!
  OBS
    LAYER ME1 ;
      RECT 0.365 1.05 0.455 1.92 ;
      RECT 0.365 0.38 0.455 0.93 ;
      RECT 0.22 0.84 0.455 0.93 ;
      RECT 0.105 1.32 0.195 2.52 ;
      RECT 0 2.3 0.56 2.52 ;
      RECT 0 -0.22 0.56 0 ;
      RECT 0.105 -0.22 0.195 0.68 ;
  END
END TIE1X2

MACRO TIE1X4
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN TIE1X4 0 -0.11 ;
  SIZE 0.84 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 1.32 0.205 2.52 ;
        RECT 0.635 1.32 0.725 2.52 ;
        RECT 0 2.3 0.84 2.52 ;
    END
  END vdd!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.375 1.08 0.465 1.92 ;
    END
  END Y
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.115 -0.22 0.205 0.68 ;
        RECT 0.635 -0.22 0.725 0.68 ;
        RECT 0 -0.22 0.84 0 ;
    END
  END gnd!
  OBS
    LAYER ME1 ;
      RECT 0.375 1.08 0.465 1.92 ;
      RECT 0.375 0.38 0.465 0.97 ;
      RECT 0.115 1.32 0.205 2.52 ;
      RECT 0.635 1.32 0.725 2.52 ;
      RECT 0 2.3 0.84 2.52 ;
      RECT 0 -0.22 0.84 0 ;
      RECT 0.115 -0.22 0.205 0.68 ;
      RECT 0.635 -0.22 0.725 0.68 ;
  END
END TIE1X4

MACRO XNOR2X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN XNOR2X1 0 -0.11 ;
  SIZE 1.96 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 1.62 0.575 2.52 ;
        RECT 1.385 1.62 1.475 2.52 ;
        RECT 0 2.3 1.96 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 -0.22 0.575 0.53 ;
        RECT 1.385 -0.22 1.475 0.53 ;
        RECT 0 -0.22 1.96 0 ;
    END
  END gnd!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.93 1.72 1.03 1.82 ;
        RECT 0.93 0.4 1.03 0.5 ;
      LAYER ME2 ;
        RECT 0.93 0.37 1.03 1.92 ;
      LAYER ME1 ;
        RECT 0.9 0.23 1.06 0.53 ;
        RECT 0.9 1.62 1.06 1.92 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.3 0.915 0.72 1.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.45 0.915 1.55 1.015 ;
      LAYER ME2 ;
        RECT 1.45 0.705 1.55 1.225 ;
      LAYER ME1 ;
        RECT 1.45 0.88 1.55 1.05 ;
        RECT 0.81 0.915 1.55 1.015 ;
        RECT 0.81 0.9 1.14 1.03 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.19 1.62 0.35 1.92 ;
      RECT 0.19 0.23 0.35 0.53 ;
      RECT 0.3 0.915 0.72 1.015 ;
      RECT 0.9 1.62 1.06 1.92 ;
      RECT 0.9 0.23 1.06 0.53 ;
      RECT 0.19 1.39 1.39 1.49 ;
      RECT 0.81 0.915 1.55 1.015 ;
      RECT 0.81 0.9 1.14 1.03 ;
      RECT 1.45 0.88 1.55 1.05 ;
      RECT 0.79 0.65 1.735 0.74 ;
      RECT 1.02 1.19 1.735 1.28 ;
      RECT 1.645 0.38 1.735 1.92 ;
      RECT 0.485 1.62 0.575 2.52 ;
      RECT 1.385 1.62 1.475 2.52 ;
      RECT 0 2.3 1.96 2.52 ;
      RECT 0 -0.22 1.96 0 ;
      RECT 0.485 -0.22 0.575 0.53 ;
      RECT 1.385 -0.22 1.475 0.53 ;
    LAYER VI1 ;
      RECT 0.22 1.72 0.32 1.82 ;
      RECT 0.22 1.39 0.32 1.49 ;
      RECT 0.22 0.4 0.32 0.5 ;
      RECT 0.93 1.72 1.03 1.82 ;
      RECT 0.93 0.4 1.03 0.5 ;
      RECT 1.45 0.915 1.55 1.015 ;
    LAYER ME2 ;
      RECT 0.22 0.37 0.32 1.92 ;
      RECT 0.93 0.37 1.03 1.92 ;
      RECT 1.45 0.705 1.55 1.225 ;
  END
END XNOR2X1

MACRO XOR2X1
  CLASS CORE ;
  ORIGIN 0 0.11 ;
  FOREIGN XOR2X1 0 -0.11 ;
  SIZE 1.96 BY 2.52 ;
  SYMMETRY X Y ;
  SITE Core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 1.62 0.575 2.52 ;
        RECT 1.385 1.62 1.475 2.52 ;
        RECT 0 2.3 1.96 2.52 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0.485 -0.22 0.575 0.53 ;
        RECT 1.385 -0.22 1.475 0.53 ;
        RECT 0 -0.22 1.96 0 ;
    END
  END gnd!
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 0.93 1.72 1.03 1.82 ;
        RECT 0.93 0.4 1.03 0.5 ;
      LAYER ME2 ;
        RECT 0.93 0.37 1.03 1.92 ;
      LAYER ME1 ;
        RECT 0.9 0.23 1.06 0.53 ;
        RECT 0.9 1.62 1.06 1.92 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0.24 0.915 0.71 1.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VI1 ;
        RECT 1.45 0.915 1.55 1.015 ;
      LAYER ME2 ;
        RECT 1.45 0.715 1.55 1.235 ;
      LAYER ME1 ;
        RECT 1.45 0.88 1.55 1.05 ;
        RECT 0.81 0.915 1.55 1.015 ;
        RECT 0.81 0.9 1.14 1.03 ;
    END
  END B
  OBS
    LAYER ME1 ;
      RECT 0.19 1.62 0.35 1.92 ;
      RECT 0.19 0.23 0.35 0.53 ;
      RECT 0.24 0.915 0.71 1.015 ;
      RECT 0.9 1.62 1.06 1.92 ;
      RECT 0.9 0.23 1.06 0.53 ;
      RECT 0.19 1.39 1.39 1.49 ;
      RECT 0.81 0.915 1.55 1.015 ;
      RECT 0.81 0.9 1.14 1.03 ;
      RECT 1.45 0.88 1.55 1.05 ;
      RECT 1.01 0.65 1.735 0.74 ;
      RECT 0.79 1.19 1.735 1.28 ;
      RECT 1.645 0.38 1.735 1.92 ;
      RECT 0.485 1.62 0.575 2.52 ;
      RECT 1.385 1.62 1.475 2.52 ;
      RECT 0 2.3 1.96 2.52 ;
      RECT 0 -0.22 1.96 0 ;
      RECT 0.485 -0.22 0.575 0.53 ;
      RECT 1.385 -0.22 1.475 0.53 ;
    LAYER VI1 ;
      RECT 0.22 1.72 0.32 1.82 ;
      RECT 0.22 1.39 0.32 1.49 ;
      RECT 0.22 0.4 0.32 0.5 ;
      RECT 0.93 1.72 1.03 1.82 ;
      RECT 0.93 0.4 1.03 0.5 ;
      RECT 1.45 0.915 1.55 1.015 ;
    LAYER ME2 ;
      RECT 0.22 0.37 0.32 1.92 ;
      RECT 0.93 0.37 1.03 1.92 ;
      RECT 1.45 0.715 1.55 1.235 ;
  END
END XOR2X1

END LIBRARY
