module voter(\A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] ,
     \A[7] , \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14]
     , \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] ,
     \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] ,
     \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] ,
     \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] ,
     \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] ,
     \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
     \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
     \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] ,
     \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] ,
     \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] ,
     \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] ,
     \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] ,
     \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] , \A[105]
     , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] , \A[111] ,
     \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
     \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
     \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] ,
     \A[130] , \A[131] , \A[132] , \A[133] , \A[134] , \A[135] ,
     \A[136] , \A[137] , \A[138] , \A[139] , \A[140] , \A[141] ,
     \A[142] , \A[143] , \A[144] , \A[145] , \A[146] , \A[147] ,
     \A[148] , \A[149] , \A[150] , \A[151] , \A[152] , \A[153] ,
     \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] ,
     \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] ,
     \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] ,
     \A[172] , \A[173] , \A[174] , \A[175] , \A[176] , \A[177] ,
     \A[178] , \A[179] , \A[180] , \A[181] , \A[182] , \A[183] ,
     \A[184] , \A[185] , \A[186] , \A[187] , \A[188] , \A[189] ,
     \A[190] , \A[191] , \A[192] , \A[193] , \A[194] , \A[195] ,
     \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] ,
     \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] ,
     \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] ,
     \A[214] , \A[215] , \A[216] , \A[217] , \A[218] , \A[219] ,
     \A[220] , \A[221] , \A[222] , \A[223] , \A[224] , \A[225] ,
     \A[226] , \A[227] , \A[228] , \A[229] , \A[230] , \A[231] ,
     \A[232] , \A[233] , \A[234] , \A[235] , \A[236] , \A[237] ,
     \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] ,
     \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] ,
     \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] ,
     \A[256] , \A[257] , \A[258] , \A[259] , \A[260] , \A[261] ,
     \A[262] , \A[263] , \A[264] , \A[265] , \A[266] , \A[267] ,
     \A[268] , \A[269] , \A[270] , \A[271] , \A[272] , \A[273] ,
     \A[274] , \A[275] , \A[276] , \A[277] , \A[278] , \A[279] ,
     \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] ,
     \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] ,
     \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] ,
     \A[298] , \A[299] , \A[300] , \A[301] , \A[302] , \A[303] ,
     \A[304] , \A[305] , \A[306] , \A[307] , \A[308] , \A[309] ,
     \A[310] , \A[311] , \A[312] , \A[313] , \A[314] , \A[315] ,
     \A[316] , \A[317] , \A[318] , \A[319] , \A[320] , \A[321] ,
     \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] ,
     \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] ,
     \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] ,
     \A[340] , \A[341] , \A[342] , \A[343] , \A[344] , \A[345] ,
     \A[346] , \A[347] , \A[348] , \A[349] , \A[350] , \A[351] ,
     \A[352] , \A[353] , \A[354] , \A[355] , \A[356] , \A[357] ,
     \A[358] , \A[359] , \A[360] , \A[361] , \A[362] , \A[363] ,
     \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] ,
     \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] ,
     \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] ,
     \A[382] , \A[383] , \A[384] , \A[385] , \A[386] , \A[387] ,
     \A[388] , \A[389] , \A[390] , \A[391] , \A[392] , \A[393] ,
     \A[394] , \A[395] , \A[396] , \A[397] , \A[398] , \A[399] ,
     \A[400] , \A[401] , \A[402] , \A[403] , \A[404] , \A[405] ,
     \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] ,
     \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] ,
     \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] ,
     \A[424] , \A[425] , \A[426] , \A[427] , \A[428] , \A[429] ,
     \A[430] , \A[431] , \A[432] , \A[433] , \A[434] , \A[435] ,
     \A[436] , \A[437] , \A[438] , \A[439] , \A[440] , \A[441] ,
     \A[442] , \A[443] , \A[444] , \A[445] , \A[446] , \A[447] ,
     \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] ,
     \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] ,
     \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] ,
     \A[466] , \A[467] , \A[468] , \A[469] , \A[470] , \A[471] ,
     \A[472] , \A[473] , \A[474] , \A[475] , \A[476] , \A[477] ,
     \A[478] , \A[479] , \A[480] , \A[481] , \A[482] , \A[483] ,
     \A[484] , \A[485] , \A[486] , \A[487] , \A[488] , \A[489] ,
     \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] ,
     \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] ,
     \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] ,
     \A[508] , \A[509] , \A[510] , \A[511] , \A[512] , \A[513] ,
     \A[514] , \A[515] , \A[516] , \A[517] , \A[518] , \A[519] ,
     \A[520] , \A[521] , \A[522] , \A[523] , \A[524] , \A[525] ,
     \A[526] , \A[527] , \A[528] , \A[529] , \A[530] , \A[531] ,
     \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] ,
     \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] ,
     \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] ,
     \A[550] , \A[551] , \A[552] , \A[553] , \A[554] , \A[555] ,
     \A[556] , \A[557] , \A[558] , \A[559] , \A[560] , \A[561] ,
     \A[562] , \A[563] , \A[564] , \A[565] , \A[566] , \A[567] ,
     \A[568] , \A[569] , \A[570] , \A[571] , \A[572] , \A[573] ,
     \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] ,
     \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] ,
     \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] ,
     \A[592] , \A[593] , \A[594] , \A[595] , \A[596] , \A[597] ,
     \A[598] , \A[599] , \A[600] , \A[601] , \A[602] , \A[603] ,
     \A[604] , \A[605] , \A[606] , \A[607] , \A[608] , \A[609] ,
     \A[610] , \A[611] , \A[612] , \A[613] , \A[614] , \A[615] ,
     \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] ,
     \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] ,
     \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] ,
     \A[634] , \A[635] , \A[636] , \A[637] , \A[638] , \A[639] ,
     \A[640] , \A[641] , \A[642] , \A[643] , \A[644] , \A[645] ,
     \A[646] , \A[647] , \A[648] , \A[649] , \A[650] , \A[651] ,
     \A[652] , \A[653] , \A[654] , \A[655] , \A[656] , \A[657] ,
     \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] ,
     \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] ,
     \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] ,
     \A[676] , \A[677] , \A[678] , \A[679] , \A[680] , \A[681] ,
     \A[682] , \A[683] , \A[684] , \A[685] , \A[686] , \A[687] ,
     \A[688] , \A[689] , \A[690] , \A[691] , \A[692] , \A[693] ,
     \A[694] , \A[695] , \A[696] , \A[697] , \A[698] , \A[699] ,
     \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] ,
     \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] ,
     \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] ,
     \A[718] , \A[719] , \A[720] , \A[721] , \A[722] , \A[723] ,
     \A[724] , \A[725] , \A[726] , \A[727] , \A[728] , \A[729] ,
     \A[730] , \A[731] , \A[732] , \A[733] , \A[734] , \A[735] ,
     \A[736] , \A[737] , \A[738] , \A[739] , \A[740] , \A[741] ,
     \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] ,
     \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] ,
     \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] ,
     \A[760] , \A[761] , \A[762] , \A[763] , \A[764] , \A[765] ,
     \A[766] , \A[767] , \A[768] , \A[769] , \A[770] , \A[771] ,
     \A[772] , \A[773] , \A[774] , \A[775] , \A[776] , \A[777] ,
     \A[778] , \A[779] , \A[780] , \A[781] , \A[782] , \A[783] ,
     \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] ,
     \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] ,
     \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] ,
     \A[802] , \A[803] , \A[804] , \A[805] , \A[806] , \A[807] ,
     \A[808] , \A[809] , \A[810] , \A[811] , \A[812] , \A[813] ,
     \A[814] , \A[815] , \A[816] , \A[817] , \A[818] , \A[819] ,
     \A[820] , \A[821] , \A[822] , \A[823] , \A[824] , \A[825] ,
     \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] ,
     \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] ,
     \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] ,
     \A[844] , \A[845] , \A[846] , \A[847] , \A[848] , \A[849] ,
     \A[850] , \A[851] , \A[852] , \A[853] , \A[854] , \A[855] ,
     \A[856] , \A[857] , \A[858] , \A[859] , \A[860] , \A[861] ,
     \A[862] , \A[863] , \A[864] , \A[865] , \A[866] , \A[867] ,
     \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] ,
     \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] ,
     \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] ,
     \A[886] , \A[887] , \A[888] , \A[889] , \A[890] , \A[891] ,
     \A[892] , \A[893] , \A[894] , \A[895] , \A[896] , \A[897] ,
     \A[898] , \A[899] , \A[900] , \A[901] , \A[902] , \A[903] ,
     \A[904] , \A[905] , \A[906] , \A[907] , \A[908] , \A[909] ,
     \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] ,
     \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] ,
     \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] ,
     \A[928] , \A[929] , \A[930] , \A[931] , \A[932] , \A[933] ,
     \A[934] , \A[935] , \A[936] , \A[937] , \A[938] , \A[939] ,
     \A[940] , \A[941] , \A[942] , \A[943] , \A[944] , \A[945] ,
     \A[946] , \A[947] , \A[948] , \A[949] , \A[950] , \A[951] ,
     \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] ,
     \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] ,
     \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] ,
     \A[970] , \A[971] , \A[972] , \A[973] , \A[974] , \A[975] ,
     \A[976] , \A[977] , \A[978] , \A[979] , \A[980] , \A[981] ,
     \A[982] , \A[983] , \A[984] , \A[985] , \A[986] , \A[987] ,
     \A[988] , \A[989] , \A[990] , \A[991] , \A[992] , \A[993] ,
     \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] ,
     \A[1000] , maj);
  input \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
       \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] ,
       \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] ,
       \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] ,
       \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] ,
       \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] ,
       \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] ,
       \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
       \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
       \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] ,
       \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] ,
       \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] ,
       \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] ,
       \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] ,
       \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] ,
       \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
       \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
       \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] ,
       \A[123] , \A[124] , \A[125] , \A[126] , \A[127] , \A[128] ,
       \A[129] , \A[130] , \A[131] , \A[132] , \A[133] , \A[134] ,
       \A[135] , \A[136] , \A[137] , \A[138] , \A[139] , \A[140] ,
       \A[141] , \A[142] , \A[143] , \A[144] , \A[145] , \A[146] ,
       \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
       \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
       \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] ,
       \A[165] , \A[166] , \A[167] , \A[168] , \A[169] , \A[170] ,
       \A[171] , \A[172] , \A[173] , \A[174] , \A[175] , \A[176] ,
       \A[177] , \A[178] , \A[179] , \A[180] , \A[181] , \A[182] ,
       \A[183] , \A[184] , \A[185] , \A[186] , \A[187] , \A[188] ,
       \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
       \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
       \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] ,
       \A[207] , \A[208] , \A[209] , \A[210] , \A[211] , \A[212] ,
       \A[213] , \A[214] , \A[215] , \A[216] , \A[217] , \A[218] ,
       \A[219] , \A[220] , \A[221] , \A[222] , \A[223] , \A[224] ,
       \A[225] , \A[226] , \A[227] , \A[228] , \A[229] , \A[230] ,
       \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
       \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
       \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] ,
       \A[249] , \A[250] , \A[251] , \A[252] , \A[253] , \A[254] ,
       \A[255] , \A[256] , \A[257] , \A[258] , \A[259] , \A[260] ,
       \A[261] , \A[262] , \A[263] , \A[264] , \A[265] , \A[266] ,
       \A[267] , \A[268] , \A[269] , \A[270] , \A[271] , \A[272] ,
       \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
       \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
       \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] ,
       \A[291] , \A[292] , \A[293] , \A[294] , \A[295] , \A[296] ,
       \A[297] , \A[298] , \A[299] , \A[300] , \A[301] , \A[302] ,
       \A[303] , \A[304] , \A[305] , \A[306] , \A[307] , \A[308] ,
       \A[309] , \A[310] , \A[311] , \A[312] , \A[313] , \A[314] ,
       \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
       \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
       \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] ,
       \A[333] , \A[334] , \A[335] , \A[336] , \A[337] , \A[338] ,
       \A[339] , \A[340] , \A[341] , \A[342] , \A[343] , \A[344] ,
       \A[345] , \A[346] , \A[347] , \A[348] , \A[349] , \A[350] ,
       \A[351] , \A[352] , \A[353] , \A[354] , \A[355] , \A[356] ,
       \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
       \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
       \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] ,
       \A[375] , \A[376] , \A[377] , \A[378] , \A[379] , \A[380] ,
       \A[381] , \A[382] , \A[383] , \A[384] , \A[385] , \A[386] ,
       \A[387] , \A[388] , \A[389] , \A[390] , \A[391] , \A[392] ,
       \A[393] , \A[394] , \A[395] , \A[396] , \A[397] , \A[398] ,
       \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
       \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
       \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] ,
       \A[417] , \A[418] , \A[419] , \A[420] , \A[421] , \A[422] ,
       \A[423] , \A[424] , \A[425] , \A[426] , \A[427] , \A[428] ,
       \A[429] , \A[430] , \A[431] , \A[432] , \A[433] , \A[434] ,
       \A[435] , \A[436] , \A[437] , \A[438] , \A[439] , \A[440] ,
       \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
       \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
       \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] ,
       \A[459] , \A[460] , \A[461] , \A[462] , \A[463] , \A[464] ,
       \A[465] , \A[466] , \A[467] , \A[468] , \A[469] , \A[470] ,
       \A[471] , \A[472] , \A[473] , \A[474] , \A[475] , \A[476] ,
       \A[477] , \A[478] , \A[479] , \A[480] , \A[481] , \A[482] ,
       \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
       \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
       \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] ,
       \A[501] , \A[502] , \A[503] , \A[504] , \A[505] , \A[506] ,
       \A[507] , \A[508] , \A[509] , \A[510] , \A[511] , \A[512] ,
       \A[513] , \A[514] , \A[515] , \A[516] , \A[517] , \A[518] ,
       \A[519] , \A[520] , \A[521] , \A[522] , \A[523] , \A[524] ,
       \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
       \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
       \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] ,
       \A[543] , \A[544] , \A[545] , \A[546] , \A[547] , \A[548] ,
       \A[549] , \A[550] , \A[551] , \A[552] , \A[553] , \A[554] ,
       \A[555] , \A[556] , \A[557] , \A[558] , \A[559] , \A[560] ,
       \A[561] , \A[562] , \A[563] , \A[564] , \A[565] , \A[566] ,
       \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
       \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
       \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] ,
       \A[585] , \A[586] , \A[587] , \A[588] , \A[589] , \A[590] ,
       \A[591] , \A[592] , \A[593] , \A[594] , \A[595] , \A[596] ,
       \A[597] , \A[598] , \A[599] , \A[600] , \A[601] , \A[602] ,
       \A[603] , \A[604] , \A[605] , \A[606] , \A[607] , \A[608] ,
       \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
       \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
       \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] ,
       \A[627] , \A[628] , \A[629] , \A[630] , \A[631] , \A[632] ,
       \A[633] , \A[634] , \A[635] , \A[636] , \A[637] , \A[638] ,
       \A[639] , \A[640] , \A[641] , \A[642] , \A[643] , \A[644] ,
       \A[645] , \A[646] , \A[647] , \A[648] , \A[649] , \A[650] ,
       \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
       \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
       \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] ,
       \A[669] , \A[670] , \A[671] , \A[672] , \A[673] , \A[674] ,
       \A[675] , \A[676] , \A[677] , \A[678] , \A[679] , \A[680] ,
       \A[681] , \A[682] , \A[683] , \A[684] , \A[685] , \A[686] ,
       \A[687] , \A[688] , \A[689] , \A[690] , \A[691] , \A[692] ,
       \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
       \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
       \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] ,
       \A[711] , \A[712] , \A[713] , \A[714] , \A[715] , \A[716] ,
       \A[717] , \A[718] , \A[719] , \A[720] , \A[721] , \A[722] ,
       \A[723] , \A[724] , \A[725] , \A[726] , \A[727] , \A[728] ,
       \A[729] , \A[730] , \A[731] , \A[732] , \A[733] , \A[734] ,
       \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
       \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
       \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] ,
       \A[753] , \A[754] , \A[755] , \A[756] , \A[757] , \A[758] ,
       \A[759] , \A[760] , \A[761] , \A[762] , \A[763] , \A[764] ,
       \A[765] , \A[766] , \A[767] , \A[768] , \A[769] , \A[770] ,
       \A[771] , \A[772] , \A[773] , \A[774] , \A[775] , \A[776] ,
       \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
       \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
       \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] ,
       \A[795] , \A[796] , \A[797] , \A[798] , \A[799] , \A[800] ,
       \A[801] , \A[802] , \A[803] , \A[804] , \A[805] , \A[806] ,
       \A[807] , \A[808] , \A[809] , \A[810] , \A[811] , \A[812] ,
       \A[813] , \A[814] , \A[815] , \A[816] , \A[817] , \A[818] ,
       \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
       \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
       \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] ,
       \A[837] , \A[838] , \A[839] , \A[840] , \A[841] , \A[842] ,
       \A[843] , \A[844] , \A[845] , \A[846] , \A[847] , \A[848] ,
       \A[849] , \A[850] , \A[851] , \A[852] , \A[853] , \A[854] ,
       \A[855] , \A[856] , \A[857] , \A[858] , \A[859] , \A[860] ,
       \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
       \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
       \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] ,
       \A[879] , \A[880] , \A[881] , \A[882] , \A[883] , \A[884] ,
       \A[885] , \A[886] , \A[887] , \A[888] , \A[889] , \A[890] ,
       \A[891] , \A[892] , \A[893] , \A[894] , \A[895] , \A[896] ,
       \A[897] , \A[898] , \A[899] , \A[900] , \A[901] , \A[902] ,
       \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
       \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
       \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] ,
       \A[921] , \A[922] , \A[923] , \A[924] , \A[925] , \A[926] ,
       \A[927] , \A[928] , \A[929] , \A[930] , \A[931] , \A[932] ,
       \A[933] , \A[934] , \A[935] , \A[936] , \A[937] , \A[938] ,
       \A[939] , \A[940] , \A[941] , \A[942] , \A[943] , \A[944] ,
       \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
       \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
       \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] ,
       \A[963] , \A[964] , \A[965] , \A[966] , \A[967] , \A[968] ,
       \A[969] , \A[970] , \A[971] , \A[972] , \A[973] , \A[974] ,
       \A[975] , \A[976] , \A[977] , \A[978] , \A[979] , \A[980] ,
       \A[981] , \A[982] , \A[983] , \A[984] , \A[985] , \A[986] ,
       \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
       \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
       \A[999] , \A[1000] ;
  output maj;
  wire \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
       \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] ,
       \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] ,
       \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] ,
       \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] ,
       \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] ,
       \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] ,
       \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
       \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
       \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] ,
       \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] ,
       \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] ,
       \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] ,
       \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] ,
       \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] ,
       \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
       \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
       \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] ,
       \A[123] , \A[124] , \A[125] , \A[126] , \A[127] , \A[128] ,
       \A[129] , \A[130] , \A[131] , \A[132] , \A[133] , \A[134] ,
       \A[135] , \A[136] , \A[137] , \A[138] , \A[139] , \A[140] ,
       \A[141] , \A[142] , \A[143] , \A[144] , \A[145] , \A[146] ,
       \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
       \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
       \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] ,
       \A[165] , \A[166] , \A[167] , \A[168] , \A[169] , \A[170] ,
       \A[171] , \A[172] , \A[173] , \A[174] , \A[175] , \A[176] ,
       \A[177] , \A[178] , \A[179] , \A[180] , \A[181] , \A[182] ,
       \A[183] , \A[184] , \A[185] , \A[186] , \A[187] , \A[188] ,
       \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
       \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
       \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] ,
       \A[207] , \A[208] , \A[209] , \A[210] , \A[211] , \A[212] ,
       \A[213] , \A[214] , \A[215] , \A[216] , \A[217] , \A[218] ,
       \A[219] , \A[220] , \A[221] , \A[222] , \A[223] , \A[224] ,
       \A[225] , \A[226] , \A[227] , \A[228] , \A[229] , \A[230] ,
       \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
       \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
       \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] ,
       \A[249] , \A[250] , \A[251] , \A[252] , \A[253] , \A[254] ,
       \A[255] , \A[256] , \A[257] , \A[258] , \A[259] , \A[260] ,
       \A[261] , \A[262] , \A[263] , \A[264] , \A[265] , \A[266] ,
       \A[267] , \A[268] , \A[269] , \A[270] , \A[271] , \A[272] ,
       \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
       \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
       \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] ,
       \A[291] , \A[292] , \A[293] , \A[294] , \A[295] , \A[296] ,
       \A[297] , \A[298] , \A[299] , \A[300] , \A[301] , \A[302] ,
       \A[303] , \A[304] , \A[305] , \A[306] , \A[307] , \A[308] ,
       \A[309] , \A[310] , \A[311] , \A[312] , \A[313] , \A[314] ,
       \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
       \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
       \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] ,
       \A[333] , \A[334] , \A[335] , \A[336] , \A[337] , \A[338] ,
       \A[339] , \A[340] , \A[341] , \A[342] , \A[343] , \A[344] ,
       \A[345] , \A[346] , \A[347] , \A[348] , \A[349] , \A[350] ,
       \A[351] , \A[352] , \A[353] , \A[354] , \A[355] , \A[356] ,
       \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
       \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
       \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] ,
       \A[375] , \A[376] , \A[377] , \A[378] , \A[379] , \A[380] ,
       \A[381] , \A[382] , \A[383] , \A[384] , \A[385] , \A[386] ,
       \A[387] , \A[388] , \A[389] , \A[390] , \A[391] , \A[392] ,
       \A[393] , \A[394] , \A[395] , \A[396] , \A[397] , \A[398] ,
       \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
       \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
       \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] ,
       \A[417] , \A[418] , \A[419] , \A[420] , \A[421] , \A[422] ,
       \A[423] , \A[424] , \A[425] , \A[426] , \A[427] , \A[428] ,
       \A[429] , \A[430] , \A[431] , \A[432] , \A[433] , \A[434] ,
       \A[435] , \A[436] , \A[437] , \A[438] , \A[439] , \A[440] ,
       \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
       \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
       \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] ,
       \A[459] , \A[460] , \A[461] , \A[462] , \A[463] , \A[464] ,
       \A[465] , \A[466] , \A[467] , \A[468] , \A[469] , \A[470] ,
       \A[471] , \A[472] , \A[473] , \A[474] , \A[475] , \A[476] ,
       \A[477] , \A[478] , \A[479] , \A[480] , \A[481] , \A[482] ,
       \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
       \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
       \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] ,
       \A[501] , \A[502] , \A[503] , \A[504] , \A[505] , \A[506] ,
       \A[507] , \A[508] , \A[509] , \A[510] , \A[511] , \A[512] ,
       \A[513] , \A[514] , \A[515] , \A[516] , \A[517] , \A[518] ,
       \A[519] , \A[520] , \A[521] , \A[522] , \A[523] , \A[524] ,
       \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
       \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
       \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] ,
       \A[543] , \A[544] , \A[545] , \A[546] , \A[547] , \A[548] ,
       \A[549] , \A[550] , \A[551] , \A[552] , \A[553] , \A[554] ,
       \A[555] , \A[556] , \A[557] , \A[558] , \A[559] , \A[560] ,
       \A[561] , \A[562] , \A[563] , \A[564] , \A[565] , \A[566] ,
       \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
       \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
       \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] ,
       \A[585] , \A[586] , \A[587] , \A[588] , \A[589] , \A[590] ,
       \A[591] , \A[592] , \A[593] , \A[594] , \A[595] , \A[596] ,
       \A[597] , \A[598] , \A[599] , \A[600] , \A[601] , \A[602] ,
       \A[603] , \A[604] , \A[605] , \A[606] , \A[607] , \A[608] ,
       \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
       \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
       \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] ,
       \A[627] , \A[628] , \A[629] , \A[630] , \A[631] , \A[632] ,
       \A[633] , \A[634] , \A[635] , \A[636] , \A[637] , \A[638] ,
       \A[639] , \A[640] , \A[641] , \A[642] , \A[643] , \A[644] ,
       \A[645] , \A[646] , \A[647] , \A[648] , \A[649] , \A[650] ,
       \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
       \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
       \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] ,
       \A[669] , \A[670] , \A[671] , \A[672] , \A[673] , \A[674] ,
       \A[675] , \A[676] , \A[677] , \A[678] , \A[679] , \A[680] ,
       \A[681] , \A[682] , \A[683] , \A[684] , \A[685] , \A[686] ,
       \A[687] , \A[688] , \A[689] , \A[690] , \A[691] , \A[692] ,
       \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
       \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
       \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] ,
       \A[711] , \A[712] , \A[713] , \A[714] , \A[715] , \A[716] ,
       \A[717] , \A[718] , \A[719] , \A[720] , \A[721] , \A[722] ,
       \A[723] , \A[724] , \A[725] , \A[726] , \A[727] , \A[728] ,
       \A[729] , \A[730] , \A[731] , \A[732] , \A[733] , \A[734] ,
       \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
       \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
       \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] ,
       \A[753] , \A[754] , \A[755] , \A[756] , \A[757] , \A[758] ,
       \A[759] , \A[760] , \A[761] , \A[762] , \A[763] , \A[764] ,
       \A[765] , \A[766] , \A[767] , \A[768] , \A[769] , \A[770] ,
       \A[771] , \A[772] , \A[773] , \A[774] , \A[775] , \A[776] ,
       \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
       \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
       \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] ,
       \A[795] , \A[796] , \A[797] , \A[798] , \A[799] , \A[800] ,
       \A[801] , \A[802] , \A[803] , \A[804] , \A[805] , \A[806] ,
       \A[807] , \A[808] , \A[809] , \A[810] , \A[811] , \A[812] ,
       \A[813] , \A[814] , \A[815] , \A[816] , \A[817] , \A[818] ,
       \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
       \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
       \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] ,
       \A[837] , \A[838] , \A[839] , \A[840] , \A[841] , \A[842] ,
       \A[843] , \A[844] , \A[845] , \A[846] , \A[847] , \A[848] ,
       \A[849] , \A[850] , \A[851] , \A[852] , \A[853] , \A[854] ,
       \A[855] , \A[856] , \A[857] , \A[858] , \A[859] , \A[860] ,
       \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
       \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
       \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] ,
       \A[879] , \A[880] , \A[881] , \A[882] , \A[883] , \A[884] ,
       \A[885] , \A[886] , \A[887] , \A[888] , \A[889] , \A[890] ,
       \A[891] , \A[892] , \A[893] , \A[894] , \A[895] , \A[896] ,
       \A[897] , \A[898] , \A[899] , \A[900] , \A[901] , \A[902] ,
       \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
       \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
       \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] ,
       \A[921] , \A[922] , \A[923] , \A[924] , \A[925] , \A[926] ,
       \A[927] , \A[928] , \A[929] , \A[930] , \A[931] , \A[932] ,
       \A[933] , \A[934] , \A[935] , \A[936] , \A[937] , \A[938] ,
       \A[939] , \A[940] , \A[941] , \A[942] , \A[943] , \A[944] ,
       \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
       \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
       \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] ,
       \A[963] , \A[964] , \A[965] , \A[966] , \A[967] , \A[968] ,
       \A[969] , \A[970] , \A[971] , \A[972] , \A[973] , \A[974] ,
       \A[975] , \A[976] , \A[977] , \A[978] , \A[979] , \A[980] ,
       \A[981] , \A[982] , \A[983] , \A[984] , \A[985] , \A[986] ,
       \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
       \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
       \A[999] , \A[1000] ;
  wire maj;
  wire n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010;
  wire n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  wire n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  wire n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  wire n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
  wire n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050;
  wire n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058;
  wire n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066;
  wire n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074;
  wire n1075, n1076, n1077, n1078, n1079, n1080, n1084, n1085;
  wire n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093;
  wire n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101;
  wire n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109;
  wire n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117;
  wire n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125;
  wire n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133;
  wire n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141;
  wire n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149;
  wire n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157;
  wire n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165;
  wire n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173;
  wire n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181;
  wire n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1192;
  wire n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200;
  wire n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208;
  wire n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216;
  wire n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224;
  wire n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232;
  wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240;
  wire n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248;
  wire n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256;
  wire n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264;
  wire n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272;
  wire n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;
  wire n1281, n1282, n1283, n1284, n1288, n1289, n1290, n1291;
  wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;
  wire n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307;
  wire n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;
  wire n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;
  wire n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331;
  wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
  wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
  wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
  wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
  wire n1364, n1365, n1366, n1367, n1368, n1369, n1373, n1374;
  wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
  wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
  wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
  wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
  wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
  wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
  wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
  wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
  wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
  wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
  wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
  wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
  wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
  wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
  wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
  wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
  wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
  wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
  wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
  wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
  wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
  wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
  wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
  wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
  wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
  wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
  wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
  wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
  wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
  wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
  wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
  wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
  wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
  wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
  wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
  wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
  wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
  wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
  wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
  wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
  wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
  wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
  wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
  wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
  wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
  wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
  wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1753;
  wire n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761;
  wire n1762, n1763, n1764, n1768, n1769, n1770, n1771, n1772;
  wire n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780;
  wire n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788;
  wire n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796;
  wire n1797, n1798, n1799, n1800, n1804, n1805, n1806, n1807;
  wire n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815;
  wire n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823;
  wire n1824, n1825, n1826, n1827, n1828, n1832, n1833, n1834;
  wire n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842;
  wire n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850;
  wire n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858;
  wire n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866;
  wire n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874;
  wire n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882;
  wire n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890;
  wire n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898;
  wire n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906;
  wire n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914;
  wire n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922;
  wire n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930;
  wire n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938;
  wire n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949;
  wire n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957;
  wire n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965;
  wire n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973;
  wire n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981;
  wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
  wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997;
  wire n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005;
  wire n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013;
  wire n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;
  wire n2022, n2023, n2027, n2028, n2029, n2030, n2031, n2032;
  wire n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040;
  wire n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048;
  wire n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056;
  wire n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064;
  wire n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072;
  wire n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080;
  wire n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088;
  wire n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096;
  wire n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104;
  wire n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112;
  wire n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120;
  wire n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128;
  wire n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136;
  wire n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144;
  wire n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152;
  wire n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160;
  wire n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168;
  wire n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176;
  wire n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184;
  wire n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192;
  wire n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200;
  wire n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208;
  wire n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216;
  wire n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224;
  wire n2225, n2229, n2230, n2231, n2232, n2233, n2234, n2235;
  wire n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243;
  wire n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251;
  wire n2252, n2253, n2257, n2258, n2259, n2260, n2261, n2262;
  wire n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270;
  wire n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278;
  wire n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286;
  wire n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294;
  wire n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
  wire n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310;
  wire n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318;
  wire n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326;
  wire n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334;
  wire n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342;
  wire n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
  wire n2351, n2352, n2356, n2357, n2358, n2359, n2360, n2361;
  wire n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369;
  wire n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377;
  wire n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385;
  wire n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393;
  wire n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401;
  wire n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409;
  wire n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417;
  wire n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425;
  wire n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433;
  wire n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441;
  wire n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449;
  wire n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457;
  wire n2458, n2459, n2460, n2464, n2465, n2466, n2467, n2468;
  wire n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476;
  wire n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484;
  wire n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492;
  wire n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500;
  wire n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508;
  wire n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516;
  wire n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524;
  wire n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532;
  wire n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540;
  wire n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548;
  wire n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556;
  wire n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567;
  wire n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575;
  wire n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583;
  wire n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591;
  wire n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599;
  wire n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607;
  wire n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615;
  wire n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623;
  wire n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631;
  wire n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639;
  wire n2640, n2641, n2645, n2646, n2647, n2648, n2649, n2650;
  wire n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658;
  wire n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666;
  wire n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674;
  wire n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682;
  wire n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690;
  wire n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698;
  wire n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706;
  wire n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714;
  wire n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722;
  wire n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730;
  wire n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738;
  wire n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746;
  wire n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754;
  wire n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762;
  wire n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770;
  wire n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778;
  wire n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786;
  wire n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794;
  wire n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802;
  wire n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810;
  wire n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818;
  wire n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826;
  wire n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834;
  wire n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842;
  wire n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850;
  wire n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858;
  wire n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866;
  wire n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874;
  wire n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882;
  wire n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890;
  wire n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898;
  wire n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906;
  wire n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914;
  wire n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922;
  wire n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930;
  wire n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938;
  wire n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946;
  wire n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954;
  wire n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962;
  wire n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970;
  wire n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978;
  wire n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986;
  wire n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994;
  wire n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002;
  wire n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010;
  wire n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018;
  wire n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026;
  wire n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034;
  wire n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042;
  wire n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050;
  wire n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058;
  wire n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066;
  wire n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074;
  wire n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082;
  wire n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090;
  wire n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098;
  wire n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106;
  wire n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114;
  wire n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122;
  wire n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130;
  wire n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138;
  wire n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146;
  wire n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154;
  wire n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162;
  wire n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170;
  wire n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178;
  wire n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186;
  wire n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194;
  wire n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202;
  wire n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210;
  wire n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218;
  wire n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226;
  wire n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234;
  wire n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242;
  wire n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250;
  wire n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258;
  wire n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266;
  wire n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274;
  wire n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282;
  wire n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290;
  wire n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298;
  wire n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306;
  wire n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314;
  wire n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322;
  wire n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330;
  wire n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338;
  wire n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346;
  wire n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354;
  wire n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362;
  wire n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370;
  wire n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378;
  wire n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386;
  wire n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394;
  wire n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402;
  wire n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410;
  wire n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418;
  wire n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426;
  wire n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434;
  wire n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442;
  wire n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450;
  wire n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458;
  wire n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466;
  wire n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474;
  wire n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482;
  wire n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490;
  wire n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498;
  wire n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506;
  wire n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514;
  wire n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522;
  wire n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530;
  wire n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538;
  wire n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546;
  wire n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554;
  wire n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562;
  wire n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570;
  wire n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578;
  wire n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586;
  wire n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594;
  wire n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602;
  wire n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610;
  wire n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618;
  wire n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626;
  wire n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634;
  wire n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642;
  wire n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650;
  wire n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658;
  wire n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666;
  wire n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674;
  wire n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682;
  wire n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690;
  wire n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698;
  wire n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706;
  wire n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714;
  wire n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722;
  wire n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730;
  wire n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738;
  wire n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746;
  wire n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754;
  wire n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762;
  wire n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770;
  wire n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778;
  wire n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786;
  wire n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794;
  wire n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802;
  wire n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810;
  wire n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818;
  wire n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826;
  wire n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834;
  wire n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842;
  wire n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850;
  wire n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858;
  wire n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866;
  wire n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874;
  wire n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882;
  wire n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890;
  wire n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898;
  wire n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906;
  wire n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914;
  wire n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922;
  wire n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930;
  wire n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938;
  wire n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946;
  wire n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954;
  wire n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962;
  wire n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970;
  wire n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978;
  wire n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986;
  wire n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3997;
  wire n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005;
  wire n4006, n4007, n4008, n4012, n4013, n4014, n4015, n4016;
  wire n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024;
  wire n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032;
  wire n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040;
  wire n4041, n4042, n4043, n4044, n4048, n4049, n4050, n4051;
  wire n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059;
  wire n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067;
  wire n4068, n4069, n4070, n4071, n4072, n4076, n4077, n4078;
  wire n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086;
  wire n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094;
  wire n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4105;
  wire n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113;
  wire n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121;
  wire n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129;
  wire n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140;
  wire n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148;
  wire n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4159;
  wire n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167;
  wire n4168, n4169, n4170, n4174, n4175, n4176, n4177, n4178;
  wire n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186;
  wire n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194;
  wire n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202;
  wire n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210;
  wire n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218;
  wire n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226;
  wire n4227, n4228, n4229, n4230, n4234, n4235, n4236, n4237;
  wire n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245;
  wire n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253;
  wire n4254, n4255, n4256, n4257, n4258, n4262, n4263, n4264;
  wire n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272;
  wire n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280;
  wire n4281, n4282, n4283, n4284, n4288, n4289, n4290, n4291;
  wire n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299;
  wire n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310;
  wire n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318;
  wire n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326;
  wire n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334;
  wire n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342;
  wire n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350;
  wire n4351, n4355, n4356, n4357, n4358, n4359, n4360, n4361;
  wire n4362, n4363, n4364, n4365, n4366, n4370, n4371, n4372;
  wire n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380;
  wire n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388;
  wire n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396;
  wire n4397, n4398, n4399, n4400, n4401, n4402, n4406, n4407;
  wire n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415;
  wire n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423;
  wire n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4434;
  wire n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442;
  wire n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450;
  wire n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458;
  wire n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466;
  wire n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474;
  wire n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482;
  wire n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490;
  wire n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498;
  wire n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506;
  wire n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514;
  wire n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522;
  wire n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530;
  wire n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538;
  wire n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546;
  wire n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554;
  wire n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565;
  wire n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573;
  wire n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581;
  wire n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589;
  wire n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597;
  wire n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605;
  wire n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613;
  wire n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621;
  wire n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629;
  wire n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637;
  wire n4638, n4639, n4643, n4644, n4645, n4646, n4647, n4648;
  wire n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656;
  wire n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664;
  wire n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672;
  wire n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680;
  wire n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688;
  wire n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696;
  wire n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704;
  wire n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712;
  wire n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720;
  wire n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728;
  wire n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736;
  wire n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744;
  wire n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752;
  wire n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760;
  wire n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768;
  wire n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776;
  wire n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784;
  wire n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792;
  wire n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800;
  wire n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808;
  wire n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816;
  wire n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824;
  wire n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832;
  wire n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840;
  wire n4841, n4845, n4846, n4847, n4848, n4849, n4850, n4851;
  wire n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859;
  wire n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867;
  wire n4868, n4869, n4873, n4874, n4875, n4876, n4877, n4878;
  wire n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886;
  wire n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894;
  wire n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902;
  wire n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910;
  wire n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918;
  wire n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926;
  wire n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934;
  wire n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942;
  wire n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950;
  wire n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958;
  wire n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966;
  wire n4967, n4968, n4969, n4970, n4971, n4972, n4976, n4977;
  wire n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985;
  wire n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993;
  wire n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001;
  wire n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009;
  wire n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017;
  wire n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025;
  wire n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033;
  wire n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041;
  wire n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049;
  wire n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057;
  wire n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068;
  wire n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076;
  wire n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084;
  wire n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092;
  wire n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100;
  wire n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108;
  wire n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116;
  wire n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124;
  wire n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132;
  wire n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140;
  wire n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148;
  wire n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156;
  wire n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164;
  wire n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172;
  wire n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180;
  wire n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188;
  wire n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196;
  wire n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204;
  wire n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212;
  wire n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220;
  wire n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228;
  wire n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236;
  wire n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244;
  wire n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252;
  wire n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260;
  wire n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268;
  wire n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276;
  wire n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284;
  wire n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292;
  wire n5293, n5294, n5295, n5296, n5300, n5301, n5302, n5303;
  wire n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311;
  wire n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319;
  wire n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327;
  wire n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335;
  wire n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343;
  wire n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351;
  wire n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359;
  wire n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367;
  wire n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375;
  wire n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383;
  wire n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391;
  wire n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399;
  wire n5400, n5401, n5402, n5403, n5404, n5408, n5409, n5410;
  wire n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418;
  wire n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426;
  wire n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434;
  wire n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442;
  wire n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450;
  wire n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458;
  wire n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466;
  wire n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474;
  wire n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482;
  wire n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490;
  wire n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498;
  wire n5499, n5500, n5504, n5505, n5506, n5507, n5508, n5509;
  wire n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517;
  wire n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525;
  wire n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533;
  wire n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541;
  wire n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549;
  wire n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557;
  wire n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565;
  wire n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573;
  wire n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581;
  wire n5582, n5583, n5584, n5585, n5589, n5590, n5591, n5592;
  wire n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600;
  wire n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608;
  wire n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616;
  wire n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624;
  wire n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632;
  wire n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640;
  wire n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648;
  wire n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656;
  wire n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664;
  wire n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672;
  wire n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680;
  wire n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688;
  wire n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696;
  wire n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704;
  wire n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712;
  wire n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720;
  wire n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728;
  wire n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736;
  wire n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744;
  wire n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752;
  wire n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760;
  wire n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768;
  wire n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776;
  wire n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784;
  wire n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792;
  wire n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800;
  wire n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808;
  wire n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816;
  wire n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824;
  wire n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832;
  wire n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840;
  wire n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848;
  wire n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856;
  wire n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864;
  wire n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872;
  wire n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880;
  wire n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888;
  wire n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896;
  wire n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904;
  wire n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912;
  wire n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920;
  wire n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928;
  wire n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936;
  wire n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944;
  wire n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952;
  wire n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960;
  wire n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968;
  wire n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976;
  wire n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984;
  wire n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992;
  wire n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000;
  wire n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008;
  wire n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016;
  wire n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024;
  wire n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032;
  wire n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040;
  wire n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048;
  wire n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056;
  wire n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064;
  wire n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072;
  wire n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080;
  wire n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088;
  wire n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096;
  wire n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104;
  wire n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112;
  wire n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120;
  wire n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128;
  wire n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136;
  wire n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144;
  wire n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152;
  wire n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160;
  wire n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168;
  wire n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176;
  wire n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184;
  wire n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192;
  wire n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200;
  wire n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208;
  wire n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216;
  wire n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224;
  wire n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232;
  wire n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240;
  wire n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248;
  wire n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256;
  wire n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264;
  wire n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272;
  wire n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280;
  wire n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288;
  wire n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296;
  wire n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304;
  wire n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6315;
  wire n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323;
  wire n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331;
  wire n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339;
  wire n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350;
  wire n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358;
  wire n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6369;
  wire n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377;
  wire n6378, n6379, n6380, n6384, n6385, n6386, n6387, n6388;
  wire n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396;
  wire n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404;
  wire n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412;
  wire n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420;
  wire n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428;
  wire n6429, n6430, n6431, n6432, n6436, n6437, n6438, n6439;
  wire n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447;
  wire n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458;
  wire n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466;
  wire n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474;
  wire n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482;
  wire n6483, n6487, n6488, n6489, n6490, n6491, n6492, n6493;
  wire n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501;
  wire n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509;
  wire n6510, n6511, n6515, n6516, n6517, n6518, n6519, n6520;
  wire n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528;
  wire n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536;
  wire n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544;
  wire n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552;
  wire n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560;
  wire n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568;
  wire n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576;
  wire n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584;
  wire n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592;
  wire n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600;
  wire n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608;
  wire n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616;
  wire n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624;
  wire n6625, n6626, n6627, n6628, n6632, n6633, n6634, n6635;
  wire n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643;
  wire n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651;
  wire n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659;
  wire n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667;
  wire n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675;
  wire n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683;
  wire n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691;
  wire n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699;
  wire n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707;
  wire n6708, n6709, n6710, n6711, n6712, n6713, n6717, n6718;
  wire n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726;
  wire n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734;
  wire n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742;
  wire n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750;
  wire n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758;
  wire n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766;
  wire n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774;
  wire n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782;
  wire n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790;
  wire n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798;
  wire n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806;
  wire n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814;
  wire n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822;
  wire n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830;
  wire n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838;
  wire n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846;
  wire n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854;
  wire n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862;
  wire n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870;
  wire n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878;
  wire n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886;
  wire n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894;
  wire n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902;
  wire n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910;
  wire n6911, n6912, n6913, n6914, n6915, n6919, n6920, n6921;
  wire n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929;
  wire n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937;
  wire n6938, n6939, n6940, n6941, n6942, n6943, n6947, n6948;
  wire n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956;
  wire n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964;
  wire n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972;
  wire n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980;
  wire n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988;
  wire n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996;
  wire n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004;
  wire n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012;
  wire n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020;
  wire n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028;
  wire n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036;
  wire n7037, n7038, n7039, n7040, n7041, n7042, n7046, n7047;
  wire n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055;
  wire n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063;
  wire n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071;
  wire n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079;
  wire n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087;
  wire n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095;
  wire n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103;
  wire n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111;
  wire n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119;
  wire n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127;
  wire n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135;
  wire n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143;
  wire n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7154;
  wire n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162;
  wire n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170;
  wire n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178;
  wire n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186;
  wire n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194;
  wire n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202;
  wire n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210;
  wire n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218;
  wire n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226;
  wire n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234;
  wire n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242;
  wire n7243, n7244, n7245, n7246, n7250, n7251, n7252, n7253;
  wire n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261;
  wire n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269;
  wire n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277;
  wire n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285;
  wire n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293;
  wire n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301;
  wire n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309;
  wire n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317;
  wire n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325;
  wire n7326, n7327, n7328, n7329, n7330, n7331, n7335, n7336;
  wire n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344;
  wire n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352;
  wire n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360;
  wire n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368;
  wire n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376;
  wire n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384;
  wire n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392;
  wire n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400;
  wire n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408;
  wire n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416;
  wire n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424;
  wire n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432;
  wire n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440;
  wire n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448;
  wire n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456;
  wire n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464;
  wire n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472;
  wire n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480;
  wire n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488;
  wire n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496;
  wire n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504;
  wire n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512;
  wire n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520;
  wire n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528;
  wire n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536;
  wire n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544;
  wire n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552;
  wire n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560;
  wire n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568;
  wire n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576;
  wire n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584;
  wire n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592;
  wire n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600;
  wire n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608;
  wire n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616;
  wire n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624;
  wire n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632;
  wire n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640;
  wire n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648;
  wire n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656;
  wire n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664;
  wire n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672;
  wire n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680;
  wire n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688;
  wire n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696;
  wire n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704;
  wire n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712;
  wire n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720;
  wire n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728;
  wire n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736;
  wire n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744;
  wire n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752;
  wire n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760;
  wire n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768;
  wire n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776;
  wire n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784;
  wire n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792;
  wire n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800;
  wire n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808;
  wire n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816;
  wire n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824;
  wire n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832;
  wire n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840;
  wire n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848;
  wire n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856;
  wire n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864;
  wire n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872;
  wire n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880;
  wire n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888;
  wire n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896;
  wire n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904;
  wire n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912;
  wire n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920;
  wire n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928;
  wire n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936;
  wire n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944;
  wire n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952;
  wire n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960;
  wire n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968;
  wire n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976;
  wire n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984;
  wire n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992;
  wire n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000;
  wire n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008;
  wire n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016;
  wire n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024;
  wire n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032;
  wire n8033, n8034, n8035, n8036, n8037, n8041, n8042, n8043;
  wire n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051;
  wire n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059;
  wire n8060, n8061, n8062, n8063, n8064, n8065, n8069, n8070;
  wire n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078;
  wire n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086;
  wire n8087, n8088, n8089, n8090, n8091, n8095, n8096, n8097;
  wire n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105;
  wire n8106, n8110, n8111, n8112, n8113, n8114, n8115, n8116;
  wire n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124;
  wire n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132;
  wire n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140;
  wire n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148;
  wire n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156;
  wire n8157, n8158, n8162, n8163, n8164, n8165, n8166, n8167;
  wire n8168, n8169, n8170, n8171, n8172, n8173, n8177, n8178;
  wire n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186;
  wire n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194;
  wire n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202;
  wire n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8213;
  wire n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221;
  wire n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229;
  wire n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237;
  wire n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248;
  wire n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256;
  wire n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264;
  wire n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272;
  wire n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280;
  wire n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288;
  wire n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296;
  wire n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304;
  wire n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312;
  wire n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320;
  wire n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328;
  wire n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336;
  wire n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344;
  wire n8345, n8346, n8347, n8348, n8349, n8350, n8354, n8355;
  wire n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363;
  wire n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371;
  wire n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379;
  wire n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387;
  wire n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395;
  wire n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403;
  wire n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411;
  wire n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419;
  wire n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427;
  wire n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435;
  wire n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443;
  wire n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451;
  wire n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8462;
  wire n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470;
  wire n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478;
  wire n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486;
  wire n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494;
  wire n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502;
  wire n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510;
  wire n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518;
  wire n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526;
  wire n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534;
  wire n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542;
  wire n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550;
  wire n8551, n8552, n8553, n8554, n8558, n8559, n8560, n8561;
  wire n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569;
  wire n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577;
  wire n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585;
  wire n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593;
  wire n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601;
  wire n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609;
  wire n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617;
  wire n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625;
  wire n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633;
  wire n8634, n8635, n8636, n8637, n8638, n8639, n8643, n8644;
  wire n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652;
  wire n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660;
  wire n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668;
  wire n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676;
  wire n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684;
  wire n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692;
  wire n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700;
  wire n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708;
  wire n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716;
  wire n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724;
  wire n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732;
  wire n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740;
  wire n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748;
  wire n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756;
  wire n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764;
  wire n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772;
  wire n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780;
  wire n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788;
  wire n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796;
  wire n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804;
  wire n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812;
  wire n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820;
  wire n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828;
  wire n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836;
  wire n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844;
  wire n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852;
  wire n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860;
  wire n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868;
  wire n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876;
  wire n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884;
  wire n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892;
  wire n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900;
  wire n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908;
  wire n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916;
  wire n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924;
  wire n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932;
  wire n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940;
  wire n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948;
  wire n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956;
  wire n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964;
  wire n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972;
  wire n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980;
  wire n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988;
  wire n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996;
  wire n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004;
  wire n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012;
  wire n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9023;
  wire n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031;
  wire n9032, n9033, n9034, n9038, n9039, n9040, n9041, n9042;
  wire n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050;
  wire n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058;
  wire n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066;
  wire n9067, n9068, n9069, n9070, n9074, n9075, n9076, n9077;
  wire n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085;
  wire n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093;
  wire n9094, n9095, n9096, n9097, n9098, n9102, n9103, n9104;
  wire n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112;
  wire n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120;
  wire n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128;
  wire n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136;
  wire n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144;
  wire n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152;
  wire n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160;
  wire n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168;
  wire n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176;
  wire n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184;
  wire n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192;
  wire n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200;
  wire n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208;
  wire n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219;
  wire n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227;
  wire n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235;
  wire n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243;
  wire n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251;
  wire n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259;
  wire n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267;
  wire n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275;
  wire n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283;
  wire n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291;
  wire n9292, n9293, n9297, n9298, n9299, n9300, n9301, n9302;
  wire n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310;
  wire n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318;
  wire n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326;
  wire n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334;
  wire n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342;
  wire n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350;
  wire n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358;
  wire n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366;
  wire n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374;
  wire n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382;
  wire n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390;
  wire n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398;
  wire n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406;
  wire n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414;
  wire n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422;
  wire n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430;
  wire n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438;
  wire n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446;
  wire n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454;
  wire n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462;
  wire n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470;
  wire n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478;
  wire n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486;
  wire n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494;
  wire n9495, n9499, n9500, n9501, n9502, n9503, n9504, n9505;
  wire n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513;
  wire n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521;
  wire n9522, n9523, n9527, n9528, n9529, n9530, n9531, n9532;
  wire n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540;
  wire n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548;
  wire n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556;
  wire n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564;
  wire n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572;
  wire n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580;
  wire n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588;
  wire n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596;
  wire n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604;
  wire n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612;
  wire n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620;
  wire n9621, n9622, n9626, n9627, n9628, n9629, n9630, n9631;
  wire n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639;
  wire n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647;
  wire n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655;
  wire n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663;
  wire n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671;
  wire n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679;
  wire n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687;
  wire n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695;
  wire n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703;
  wire n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711;
  wire n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719;
  wire n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727;
  wire n9728, n9729, n9730, n9734, n9735, n9736, n9737, n9738;
  wire n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746;
  wire n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754;
  wire n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762;
  wire n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770;
  wire n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778;
  wire n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786;
  wire n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794;
  wire n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802;
  wire n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810;
  wire n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818;
  wire n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826;
  wire n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837;
  wire n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845;
  wire n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853;
  wire n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861;
  wire n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869;
  wire n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877;
  wire n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885;
  wire n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893;
  wire n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901;
  wire n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909;
  wire n9910, n9911, n9915, n9916, n9917, n9918, n9919, n9920;
  wire n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928;
  wire n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936;
  wire n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944;
  wire n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952;
  wire n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960;
  wire n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968;
  wire n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976;
  wire n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984;
  wire n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992;
  wire n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000;
  wire n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008;
  wire n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016;
  wire n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024;
  wire n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032;
  wire n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040;
  wire n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048;
  wire n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056;
  wire n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064;
  wire n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072;
  wire n10073, n10074, n10077, n10078, n10079, n10080, n10081, n10082;
  wire n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090;
  wire n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100;
  wire n10101, n10102, n10103, n10104, n10107, n10108, n10109, n10110;
  wire n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118;
  wire n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126;
  wire n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134;
  wire n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144;
  wire n10145, n10146, n10147, n10148, n10151, n10152, n10153, n10154;
  wire n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162;
  wire n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170;
  wire n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180;
  wire n10181, n10182, n10183, n10184, n10187, n10188, n10189, n10190;
  wire n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198;
  wire n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206;
  wire n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214;
  wire n10215, n10216, n10217, n10218, n10219, n10222, n10223, n10224;
  wire n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232;
  wire n10233, n10236, n10237, n10238, n10239, n10240, n10241, n10242;
  wire n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250;
  wire n10251, n10252, n10253, n10254, n10255, n10258, n10259, n10260;
  wire n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268;
  wire n10269, n10272, n10273, n10274, n10275, n10276, n10277, n10278;
  wire n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286;
  wire n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294;
  wire n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302;
  wire n10303, n10304, n10305, n10306, n10307, n10308, n10311, n10312;
  wire n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320;
  wire n10321, n10322, n10325, n10326, n10327, n10328, n10329, n10330;
  wire n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338;
  wire n10339, n10340, n10341, n10342, n10343, n10344, n10347, n10348;
  wire n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356;
  wire n10357, n10358, n10361, n10362, n10363, n10364, n10365, n10366;
  wire n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374;
  wire n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382;
  wire n10383, n10384, n10385, n10386, n10387, n10388, n10391, n10392;
  wire n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400;
  wire n10401, n10402, n10405, n10406, n10407, n10408, n10409, n10410;
  wire n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418;
  wire n10419, n10420, n10421, n10422, n10423, n10424, n10427, n10428;
  wire n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436;
  wire n10437, n10438, n10441, n10442, n10443, n10444, n10445, n10446;
  wire n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454;
  wire n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462;
  wire n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470;
  wire n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478;
  wire n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486;
  wire n10487, n10488, n10491, n10492, n10493, n10494, n10495, n10496;
  wire n10497, n10498, n10499, n10500, n10501, n10502, n10505, n10506;
  wire n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514;
  wire n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522;
  wire n10523, n10524, n10527, n10528, n10529, n10530, n10531, n10532;
  wire n10533, n10534, n10535, n10536, n10537, n10538, n10541, n10542;
  wire n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550;
  wire n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558;
  wire n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566;
  wire n10567, n10568, n10571, n10572, n10573, n10574, n10575, n10576;
  wire n10577, n10578, n10579, n10580, n10581, n10582, n10585, n10586;
  wire n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594;
  wire n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602;
  wire n10603, n10604, n10607, n10608, n10609, n10610, n10611, n10612;
  wire n10613, n10614, n10615, n10616, n10617, n10618, n10621, n10622;
  wire n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630;
  wire n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638;
  wire n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646;
  wire n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654;
  wire n10655, n10656, n10659, n10660, n10661, n10662, n10663, n10664;
  wire n10665, n10666, n10667, n10668, n10669, n10670, n10673, n10674;
  wire n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682;
  wire n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690;
  wire n10691, n10692, n10695, n10696, n10697, n10698, n10699, n10700;
  wire n10701, n10702, n10703, n10704, n10705, n10706, n10709, n10710;
  wire n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718;
  wire n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726;
  wire n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734;
  wire n10735, n10736, n10739, n10740, n10741, n10742, n10743, n10744;
  wire n10745, n10746, n10747, n10748, n10749, n10750, n10753, n10754;
  wire n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762;
  wire n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770;
  wire n10771, n10772, n10775, n10776, n10777, n10778, n10779, n10780;
  wire n10781, n10782, n10783, n10784, n10785, n10786, n10789, n10790;
  wire n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798;
  wire n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806;
  wire n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814;
  wire n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822;
  wire n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830;
  wire n10831, n10832, n10835, n10836, n10837, n10838, n10839, n10840;
  wire n10841, n10842, n10843, n10844, n10845, n10846, n10849, n10850;
  wire n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858;
  wire n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866;
  wire n10867, n10868, n10871, n10872, n10873, n10874, n10875, n10876;
  wire n10877, n10878, n10879, n10880, n10881, n10882, n10885, n10886;
  wire n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894;
  wire n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902;
  wire n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910;
  wire n10911, n10912, n10915, n10916, n10917, n10918, n10919, n10920;
  wire n10921, n10922, n10923, n10924, n10925, n10926, n10929, n10930;
  wire n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938;
  wire n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946;
  wire n10947, n10948, n10951, n10952, n10953, n10954, n10955, n10956;
  wire n10957, n10958, n10959, n10960, n10961, n10962, n10965, n10966;
  wire n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974;
  wire n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982;
  wire n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990;
  wire n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998;
  wire n10999, n11000, n11003, n11004, n11005, n11006, n11007, n11008;
  wire n11009, n11010, n11011, n11012, n11013, n11014, n11017, n11018;
  wire n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026;
  wire n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034;
  wire n11035, n11036, n11039, n11040, n11041, n11042, n11043, n11044;
  wire n11045, n11046, n11047, n11048, n11049, n11050, n11053, n11054;
  wire n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062;
  wire n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070;
  wire n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078;
  wire n11079, n11080, n11083, n11084, n11085, n11086, n11087, n11088;
  wire n11089, n11090, n11091, n11092, n11093, n11094, n11097, n11098;
  wire n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106;
  wire n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114;
  wire n11115, n11116, n11119, n11120, n11121, n11122, n11123, n11124;
  wire n11125, n11126, n11127, n11128, n11129, n11130, n11133, n11134;
  wire n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142;
  wire n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150;
  wire n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158;
  wire n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166;
  wire n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174;
  wire n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182;
  wire n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190;
  wire n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200;
  wire n11201, n11202, n11203, n11204, n11207, n11208, n11209, n11210;
  wire n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218;
  wire n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226;
  wire n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236;
  wire n11237, n11238, n11239, n11240, n11243, n11244, n11245, n11246;
  wire n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254;
  wire n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262;
  wire n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270;
  wire n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280;
  wire n11281, n11282, n11283, n11284, n11287, n11288, n11289, n11290;
  wire n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298;
  wire n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306;
  wire n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316;
  wire n11317, n11318, n11319, n11320, n11323, n11324, n11325, n11326;
  wire n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334;
  wire n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342;
  wire n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350;
  wire n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358;
  wire n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368;
  wire n11369, n11370, n11371, n11372, n11375, n11376, n11377, n11378;
  wire n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386;
  wire n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394;
  wire n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404;
  wire n11405, n11406, n11407, n11408, n11411, n11412, n11413, n11414;
  wire n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422;
  wire n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430;
  wire n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438;
  wire n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448;
  wire n11449, n11450, n11451, n11452, n11455, n11456, n11457, n11458;
  wire n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466;
  wire n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474;
  wire n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484;
  wire n11485, n11486, n11487, n11488, n11491, n11492, n11493, n11494;
  wire n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502;
  wire n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510;
  wire n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518;
  wire n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526;
  wire n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534;
  wire n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544;
  wire n11545, n11546, n11547, n11548, n11551, n11552, n11553, n11554;
  wire n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562;
  wire n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570;
  wire n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580;
  wire n11581, n11582, n11583, n11584, n11587, n11588, n11589, n11590;
  wire n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598;
  wire n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606;
  wire n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614;
  wire n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624;
  wire n11625, n11626, n11627, n11628, n11631, n11632, n11633, n11634;
  wire n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642;
  wire n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650;
  wire n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660;
  wire n11661, n11662, n11663, n11664, n11667, n11668, n11669, n11670;
  wire n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678;
  wire n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686;
  wire n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694;
  wire n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702;
  wire n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712;
  wire n11713, n11714, n11715, n11716, n11719, n11720, n11721, n11722;
  wire n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730;
  wire n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738;
  wire n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748;
  wire n11749, n11750, n11751, n11752, n11755, n11756, n11757, n11758;
  wire n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766;
  wire n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774;
  wire n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782;
  wire n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792;
  wire n11793, n11794, n11795, n11796, n11799, n11800, n11801, n11802;
  wire n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810;
  wire n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818;
  wire n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828;
  wire n11829, n11830, n11831, n11832, n11835, n11836, n11837, n11838;
  wire n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846;
  wire n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854;
  wire n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862;
  wire n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870;
  wire n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878;
  wire n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886;
  wire n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11896;
  wire n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904;
  wire n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11914;
  wire n11915, n11916, n11917, n11920, n11921, n11922, n11923, n11924;
  wire n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932;
  wire n11933, n11934, n11935, n11938, n11939, n11940, n11941, n11942;
  wire n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950;
  wire n11951, n11954, n11955, n11956, n11957, n11958, n11959, n11960;
  wire n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968;
  wire n11969, n11972, n11973, n11974, n11975, n11978, n11979, n11980;
  wire n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988;
  wire n11989, n11990, n11991, n11992, n11993, n11996, n11997, n11998;
  wire n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006;
  wire n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014;
  wire n12015, n12016, n12017, n12018, n12019, n12022, n12023, n12024;
  wire n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032;
  wire n12033, n12034, n12035, n12036, n12037, n12040, n12041, n12042;
  wire n12043, n12046, n12047, n12048, n12049, n12050, n12051, n12052;
  wire n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060;
  wire n12061, n12064, n12065, n12066, n12067, n12068, n12069, n12070;
  wire n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12080;
  wire n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088;
  wire n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12098;
  wire n12099, n12100, n12101, n12104, n12105, n12106, n12107, n12108;
  wire n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116;
  wire n12117, n12118, n12119, n12122, n12123, n12124, n12125, n12126;
  wire n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134;
  wire n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142;
  wire n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150;
  wire n12151, n12152, n12153, n12154, n12155, n12158, n12159, n12160;
  wire n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168;
  wire n12169, n12170, n12171, n12172, n12173, n12176, n12177, n12178;
  wire n12179, n12182, n12183, n12184, n12185, n12186, n12187, n12188;
  wire n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196;
  wire n12197, n12200, n12201, n12202, n12203, n12204, n12205, n12206;
  wire n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12216;
  wire n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224;
  wire n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12234;
  wire n12235, n12236, n12237, n12240, n12241, n12242, n12243, n12244;
  wire n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252;
  wire n12253, n12254, n12255, n12258, n12259, n12260, n12261, n12262;
  wire n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270;
  wire n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278;
  wire n12279, n12280, n12281, n12284, n12285, n12286, n12287, n12288;
  wire n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296;
  wire n12297, n12298, n12299, n12302, n12303, n12304, n12305, n12308;
  wire n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316;
  wire n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12326;
  wire n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334;
  wire n12335, n12336, n12337, n12338, n12339, n12342, n12343, n12344;
  wire n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352;
  wire n12353, n12354, n12355, n12356, n12357, n12360, n12361, n12362;
  wire n12363, n12366, n12367, n12368, n12369, n12370, n12371, n12372;
  wire n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380;
  wire n12381, n12384, n12385, n12386, n12387, n12388, n12389, n12390;
  wire n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398;
  wire n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406;
  wire n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414;
  wire n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422;
  wire n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12432;
  wire n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440;
  wire n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12450;
  wire n12451, n12452, n12453, n12456, n12457, n12458, n12459, n12460;
  wire n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468;
  wire n12469, n12470, n12471, n12474, n12475, n12476, n12477, n12478;
  wire n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486;
  wire n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494;
  wire n12495, n12496, n12497, n12498, n12501, n12502, n12503, n12504;
  wire n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512;
  wire n12513, n12514, n12515, n12516, n12519, n12520, n12521, n12522;
  wire n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530;
  wire n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538;
  wire n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548;
  wire n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556;
  wire n12559, n12560, n12561, n12562, n12565, n12566, n12567, n12568;
  wire n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576;
  wire n12577, n12578, n12579, n12580, n12583, n12584, n12585, n12586;
  wire n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594;
  wire n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602;
  wire n12603, n12604, n12605, n12606, n12607, n12610, n12611, n12612;
  wire n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620;
  wire n12621, n12622, n12623, n12624, n12625, n12628, n12629, n12630;
  wire n12631, n12634, n12635, n12636, n12637, n12638, n12639, n12640;
  wire n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648;
  wire n12649, n12652, n12653, n12654, n12655, n12656, n12657, n12658;
  wire n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12668;
  wire n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676;
  wire n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12686;
  wire n12687, n12688, n12689, n12692, n12693, n12694, n12695, n12696;
  wire n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704;
  wire n12705, n12706, n12707, n12710, n12711, n12712, n12713, n12714;
  wire n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722;
  wire n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730;
  wire n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738;
  wire n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746;
  wire n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754;
  wire n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764;
  wire n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772;
  wire n12775, n12776, n12777, n12778, n12781, n12782, n12783, n12784;
  wire n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792;
  wire n12793, n12794, n12795, n12796, n12799, n12800, n12801, n12802;
  wire n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810;
  wire n12811, n12812, n12815, n12816, n12817, n12818, n12819, n12820;
  wire n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828;
  wire n12829, n12830, n12833, n12834, n12835, n12836, n12839, n12840;
  wire n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848;
  wire n12849, n12850, n12851, n12852, n12853, n12854, n12857, n12858;
  wire n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866;
  wire n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874;
  wire n12875, n12876, n12877, n12878, n12879, n12880, n12883, n12884;
  wire n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892;
  wire n12893, n12894, n12895, n12896, n12897, n12898, n12901, n12902;
  wire n12903, n12904, n12907, n12908, n12909, n12910, n12911, n12912;
  wire n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920;
  wire n12921, n12922, n12925, n12926, n12927, n12928, n12929, n12930;
  wire n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938;
  wire n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948;
  wire n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956;
  wire n12959, n12960, n12961, n12962, n12965, n12966, n12967, n12968;
  wire n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976;
  wire n12977, n12978, n12979, n12980, n12983, n12984, n12985, n12986;
  wire n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994;
  wire n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002;
  wire n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010;
  wire n13011, n13012, n13013, n13014, n13015, n13016, n13019, n13020;
  wire n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028;
  wire n13029, n13030, n13031, n13032, n13033, n13034, n13037, n13038;
  wire n13039, n13040, n13043, n13044, n13045, n13046, n13047, n13048;
  wire n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056;
  wire n13057, n13058, n13061, n13062, n13063, n13064, n13065, n13066;
  wire n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074;
  wire n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084;
  wire n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092;
  wire n13095, n13096, n13097, n13098, n13101, n13102, n13103, n13104;
  wire n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112;
  wire n13113, n13114, n13115, n13116, n13119, n13120, n13121, n13122;
  wire n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130;
  wire n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138;
  wire n13139, n13140, n13141, n13142, n13145, n13146, n13147, n13148;
  wire n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156;
  wire n13157, n13158, n13159, n13160, n13163, n13164, n13165, n13166;
  wire n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176;
  wire n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184;
  wire n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194;
  wire n13195, n13196, n13197, n13198, n13199, n13200, n13203, n13204;
  wire n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212;
  wire n13213, n13214, n13215, n13216, n13217, n13218, n13221, n13222;
  wire n13223, n13224, n13227, n13228, n13229, n13230, n13231, n13232;
  wire n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240;
  wire n13241, n13242, n13245, n13246, n13247, n13248, n13249, n13250;
  wire n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258;
  wire n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266;
  wire n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274;
  wire n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282;
  wire n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290;
  wire n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298;
  wire n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306;
  wire n13307, n13308, n13309, n13312, n13313, n13314, n13315, n13316;
  wire n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324;
  wire n13325, n13328, n13329, n13330, n13331, n13332, n13333, n13334;
  wire n13335, n13336, n13339, n13340, n13341, n13342, n13343, n13344;
  wire n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352;
  wire n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362;
  wire n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13372;
  wire n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380;
  wire n13381, n13382, n13383, n13384, n13385, n13388, n13389, n13390;
  wire n13391, n13394, n13395, n13396, n13397, n13398, n13399, n13400;
  wire n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13410;
  wire n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418;
  wire n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426;
  wire n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434;
  wire n13435, n13436, n13437, n13438, n13439, n13442, n13443, n13444;
  wire n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452;
  wire n13453, n13454, n13455, n13458, n13459, n13460, n13461, n13464;
  wire n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472;
  wire n13473, n13474, n13475, n13476, n13477, n13480, n13481, n13482;
  wire n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490;
  wire n13491, n13492, n13493, n13496, n13497, n13498, n13499, n13500;
  wire n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508;
  wire n13509, n13512, n13513, n13514, n13515, n13518, n13519, n13520;
  wire n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528;
  wire n13529, n13530, n13531, n13534, n13535, n13536, n13537, n13538;
  wire n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546;
  wire n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554;
  wire n13555, n13556, n13557, n13560, n13561, n13562, n13563, n13564;
  wire n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572;
  wire n13573, n13576, n13577, n13578, n13579, n13582, n13583, n13584;
  wire n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592;
  wire n13593, n13594, n13595, n13598, n13599, n13600, n13601, n13602;
  wire n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610;
  wire n13611, n13614, n13615, n13616, n13617, n13618, n13619, n13620;
  wire n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13630;
  wire n13631, n13632, n13633, n13636, n13637, n13638, n13639, n13640;
  wire n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648;
  wire n13649, n13652, n13653, n13654, n13655, n13656, n13657, n13658;
  wire n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666;
  wire n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674;
  wire n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682;
  wire n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690;
  wire n13691, n13694, n13695, n13696, n13697, n13698, n13699, n13700;
  wire n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13710;
  wire n13711, n13712, n13713, n13716, n13717, n13718, n13719, n13720;
  wire n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728;
  wire n13729, n13732, n13733, n13734, n13735, n13736, n13737, n13738;
  wire n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13748;
  wire n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756;
  wire n13757, n13758, n13759, n13760, n13761, n13764, n13765, n13766;
  wire n13767, n13770, n13771, n13772, n13773, n13774, n13775, n13776;
  wire n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13786;
  wire n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794;
  wire n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802;
  wire n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13812;
  wire n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820;
  wire n13821, n13822, n13823, n13824, n13825, n13828, n13829, n13830;
  wire n13831, n13834, n13835, n13836, n13837, n13838, n13839, n13840;
  wire n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13850;
  wire n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858;
  wire n13859, n13860, n13861, n13862, n13863, n13866, n13867, n13868;
  wire n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876;
  wire n13877, n13878, n13879, n13882, n13883, n13884, n13885, n13888;
  wire n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896;
  wire n13897, n13898, n13899, n13900, n13901, n13904, n13905, n13906;
  wire n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914;
  wire n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922;
  wire n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930;
  wire n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938;
  wire n13939, n13940, n13941, n13942, n13945, n13946, n13949, n13950;
  wire n13951, n13952, n13955, n13956, n13957, n13958, n13959, n13960;
  wire n13961, n13962, n13965, n13966, n13967, n13968, n13971, n13972;
  wire n13975, n13976, n13977, n13978, n13981, n13982, n13983, n13984;
  wire n13985, n13986, n13987, n13988, n13991, n13992, n13993, n13994;
  wire n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002;
  wire n14003, n14004, n14007, n14008, n14011, n14012, n14013, n14014;
  wire n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024;
  wire n14027, n14028, n14029, n14030, n14033, n14034, n14037, n14038;
  wire n14039, n14040, n14043, n14044, n14045, n14046, n14047, n14048;
  wire n14049, n14050, n14053, n14054, n14055, n14056, n14057, n14058;
  wire n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066;
  wire n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074;
  wire n14075, n14076, n14077, n14078, n14081, n14082, n14085, n14086;
  wire n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094;
  wire n14097, n14100, n14101, n14102, n14103, n14104, n14105, n14106;
  wire n14107, n14108, n14109, n14112, n14113, n14114, n14115, n14118;
  wire n14119, n14122, n14123, n14124, n14125, n14128, n14129, n14130;
  wire n14131, n14132, n14133, n14134, n14135, n14138, n14139, n14140;
  wire n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148;
  wire n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156;
  wire n14157, n14158, n14159, n14160, n14161, n14162, n14165, n14166;
  wire n14169, n14170, n14171, n14172, n14175, n14176, n14177, n14178;
  wire n14179, n14180, n14181, n14182, n14185, n14186, n14187, n14188;
  wire n14191, n14192, n14195, n14196, n14197, n14198, n14201, n14202;
  wire n14203, n14204, n14205, n14206, n14207, n14208, n14211, n14212;
  wire n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220;
  wire n14221, n14222, n14223, n14224, n14227, n14228, n14231, n14232;
  wire n14233, n14234, n14237, n14238, n14239, n14240, n14241, n14242;
  wire n14243, n14244, n14247, n14248, n14249, n14250, n14253, n14254;
  wire n14257, n14258, n14259, n14260, n14263, n14264, n14265, n14266;
  wire n14267, n14268, n14269, n14270, n14273, n14274, n14275, n14276;
  wire n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284;
  wire n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292;
  wire n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300;
  wire n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310;
  wire n14311, n14314, n14315, n14316, n14317, n14318, n14319, n14320;
  wire n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328;
  wire n14329, n14330, n14331, n14332, n14333, n14334, n14337, n14338;
  wire n14341, n14342, n14343, n14344, n14347, n14348, n14349, n14350;
  wire n14351, n14352, n14353, n14354, n14357, n14358, n14359, n14360;
  wire n14363, n14364, n14367, n14368, n14369, n14370, n14373, n14374;
  wire n14375, n14376, n14377, n14378, n14379, n14380, n14383, n14384;
  wire n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392;
  wire n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400;
  wire n14401, n14402, n14405, n14406, n14409, n14410, n14411, n14412;
  wire n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422;
  wire n14425, n14426, n14427, n14428, n14431, n14432, n14435, n14436;
  wire n14437, n14438, n14441, n14442, n14443, n14444, n14445, n14446;
  wire n14447, n14448, n14451, n14452, n14453, n14454, n14455, n14456;
  wire n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464;
  wire n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472;
  wire n14473, n14474, n14475, n14476, n14479, n14480, n14483, n14484;
  wire n14485, n14486, n14489, n14490, n14491, n14492, n14493, n14494;
  wire n14495, n14496, n14499, n14500, n14501, n14504, n14505, n14506;
  wire n14507, n14508, n14509, n14510, n14513, n14514, n14517, n14518;
  wire n14519, n14520, n14523, n14524, n14525, n14526, n14527, n14528;
  wire n14529, n14530, n14533, n14534, n14535, n14536, n14537, n14538;
  wire n14539, n14540, n14541, n14544, n14545, n14546, n14547, n14548;
  wire n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14558;
  wire n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566;
  wire n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574;
  wire n14575, n14578, n14579, n14580, n14581, n14582, n14583, n14584;
  wire n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592;
  wire n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600;
  wire n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608;
  wire n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616;
  wire n14617, n14618, n14619, n14620, n14622, n14623, n14624, n14625;
  wire n14626, n14627, n14628, n14629, n14630, n14632, n14633, n14634;
  wire n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642;
  wire n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650;
  wire n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658;
  wire n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666;
  wire n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674;
  wire n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682;
  wire n14683, n14684, n14685, n14686, n14692, n14695, n14696, n14697;
  wire n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705;
  wire n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713;
  wire n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721;
  wire n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729;
  wire n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737;
  wire n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745;
  wire n14746, n14747, n14748, n14749, n14750, n14753, n14754, n14755;
  wire n14756, n14757, n14758, n14759, n_3, n_4, n_5, n_6;
  wire n_8, n_9, n_10, n_13, n_14, n_15, n_16, n_18;
  wire n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_47, n_48, n_49, n_50, n_52, n_53;
  wire n_54, n_57, n_58, n_59, n_60, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_105;
  wire n_107, n_109, n_110, n_111, n_112, n_113, n_114, n_116;
  wire n_118, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_149, n_151, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_160, n_162, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_226, n_227, n_228, n_229, n_231;
  wire n_232, n_233, n_236, n_237, n_238, n_239, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_270, n_271, n_272, n_273, n_275, n_276, n_277;
  wire n_280, n_281, n_282, n_283, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_327, n_328, n_329, n_330;
  wire n_332, n_333, n_334, n_337, n_338, n_339, n_340, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_371, n_372, n_373, n_374, n_376, n_377;
  wire n_378, n_381, n_382, n_383, n_384, n_386, n_387, n_388;
  wire n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444;
  wire n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_465, n_467, n_469, n_470, n_471;
  wire n_472, n_473, n_474, n_476, n_478, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_509, n_511, n_513, n_514, n_515, n_516, n_517;
  wire n_518, n_520, n_522, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_557, n_559, n_561, n_562, n_563;
  wire n_564, n_565, n_566, n_568, n_570, n_572, n_573, n_574;
  wire n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_601, n_603, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_612, n_614, n_616, n_617, n_618, n_619, n_620;
  wire n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636;
  wire n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644;
  wire n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_653;
  wire n_655, n_657, n_658, n_659, n_660, n_661, n_662, n_664;
  wire n_666, n_668, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682;
  wire n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_694, n_695, n_697, n_699, n_701;
  wire n_702, n_703, n_704, n_705, n_706, n_708, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_745;
  wire n_747, n_749, n_750, n_751, n_752, n_753, n_754, n_756;
  wire n_758, n_760, n_761, n_762, n_763, n_764, n_765, n_766;
  wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
  wire n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782;
  wire n_783, n_784, n_785, n_786, n_787, n_789, n_791, n_793;
  wire n_794, n_795, n_796, n_797, n_798, n_800, n_802, n_804;
  wire n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812;
  wire n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820;
  wire n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836;
  wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868;
  wire n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884;
  wire n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892;
  wire n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900;
  wire n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_941, n_942, n_943, n_946, n_947, n_948, n_949, n_951;
  wire n_952, n_953, n_956, n_957, n_958, n_959, n_961, n_962;
  wire n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970;
  wire n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978;
  wire n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986;
  wire n_987, n_990, n_991, n_992, n_993, n_995, n_996, n_997;
  wire n_1000, n_1001, n_1002, n_1003, n_1005, n_1006, n_1007, n_1008;
  wire n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016;
  wire n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1042, n_1043, n_1044, n_1047, n_1048, n_1049, n_1050;
  wire n_1052, n_1053, n_1054, n_1057, n_1058, n_1059, n_1060, n_1062;
  wire n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070;
  wire n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078;
  wire n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086;
  wire n_1087, n_1088, n_1091, n_1092, n_1093, n_1094, n_1096, n_1097;
  wire n_1098, n_1101, n_1102, n_1103, n_1104, n_1106, n_1107, n_1108;
  wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116;
  wire n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124;
  wire n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132;
  wire n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140;
  wire n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148;
  wire n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156;
  wire n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164;
  wire n_1165, n_1166, n_1168, n_1170, n_1172, n_1173, n_1174, n_1175;
  wire n_1176, n_1177, n_1179, n_1181, n_1183, n_1184, n_1185, n_1186;
  wire n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194;
  wire n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202;
  wire n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210;
  wire n_1212, n_1214, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221;
  wire n_1223, n_1225, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1260, n_1262, n_1264, n_1265, n_1266, n_1267;
  wire n_1268, n_1269, n_1271, n_1273, n_1275, n_1276, n_1277, n_1278;
  wire n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286;
  wire n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294;
  wire n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302;
  wire n_1304, n_1306, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313;
  wire n_1315, n_1317, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332;
  wire n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340;
  wire n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348;
  wire n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356;
  wire n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364;
  wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372;
  wire n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380;
  wire n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388;
  wire n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396;
  wire n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404;
  wire n_1405, n_1406, n_1409, n_1410, n_1411, n_1412, n_1414, n_1415;
  wire n_1416, n_1419, n_1420, n_1421, n_1422, n_1424, n_1425, n_1426;
  wire n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434;
  wire n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442;
  wire n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450;
  wire n_1453, n_1454, n_1455, n_1456, n_1458, n_1459, n_1460, n_1463;
  wire n_1464, n_1465, n_1466, n_1468, n_1469, n_1470, n_1471, n_1472;
  wire n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480;
  wire n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488;
  wire n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496;
  wire n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504;
  wire n_1505, n_1506, n_1507, n_1508, n_1509, n_1511, n_1513, n_1515;
  wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1522, n_1524, n_1526;
  wire n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534;
  wire n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542;
  wire n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550;
  wire n_1551, n_1552, n_1553, n_1555, n_1557, n_1559, n_1560, n_1561;
  wire n_1562, n_1563, n_1564, n_1566, n_1568, n_1570, n_1571, n_1572;
  wire n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580;
  wire n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588;
  wire n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596;
  wire n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604;
  wire n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612;
  wire n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620;
  wire n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628;
  wire n_1629, n_1632, n_1633, n_1634, n_1635, n_1637, n_1638, n_1639;
  wire n_1642, n_1643, n_1644, n_1645, n_1647, n_1648, n_1649, n_1650;
  wire n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658;
  wire n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666;
  wire n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1676;
  wire n_1677, n_1678, n_1679, n_1681, n_1682, n_1683, n_1686, n_1687;
  wire n_1688, n_1689, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
  wire n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720;
  wire n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728;
  wire n_1729, n_1730, n_1733, n_1734, n_1735, n_1736, n_1738, n_1739;
  wire n_1740, n_1743, n_1744, n_1745, n_1746, n_1748, n_1749, n_1750;
  wire n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758;
  wire n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766;
  wire n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774;
  wire n_1777, n_1778, n_1779, n_1780, n_1782, n_1783, n_1784, n_1787;
  wire n_1788, n_1789, n_1790, n_1792, n_1793, n_1794, n_1795, n_1796;
  wire n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804;
  wire n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812;
  wire n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820;
  wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836;
  wire n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844;
  wire n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852;
  wire n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860;
  wire n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868;
  wire n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876;
  wire n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884;
  wire n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892;
  wire n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900;
  wire n_1901, n_1903, n_1905, n_1907, n_1908, n_1909, n_1910, n_1911;
  wire n_1912, n_1914, n_1916, n_1918, n_1919, n_1920, n_1921, n_1922;
  wire n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930;
  wire n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938;
  wire n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1947;
  wire n_1949, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1958;
  wire n_1960, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976;
  wire n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984;
  wire n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992;
  wire n_1993, n_1995, n_1997, n_1999, n_2000, n_2001, n_2002, n_2003;
  wire n_2004, n_2006, n_2008, n_2010, n_2011, n_2012, n_2013, n_2014;
  wire n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022;
  wire n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030;
  wire n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2039;
  wire n_2041, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2050;
  wire n_2052, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060;
  wire n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068;
  wire n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076;
  wire n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084;
  wire n_2085, n_2086, n_2087, n_2088, n_2089, n_2091, n_2093, n_2095;
  wire n_2096, n_2097, n_2098, n_2099, n_2100, n_2102, n_2104, n_2106;
  wire n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114;
  wire n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122;
  wire n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130;
  wire n_2131, n_2132, n_2133, n_2135, n_2137, n_2139, n_2140, n_2141;
  wire n_2142, n_2143, n_2144, n_2146, n_2148, n_2150, n_2151, n_2152;
  wire n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160;
  wire n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168;
  wire n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176;
  wire n_2177, n_2178, n_2179, n_2180, n_2181, n_2183, n_2185, n_2187;
  wire n_2188, n_2189, n_2190, n_2191, n_2192, n_2194, n_2196, n_2198;
  wire n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206;
  wire n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214;
  wire n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222;
  wire n_2223, n_2224, n_2225, n_2227, n_2229, n_2231, n_2232, n_2233;
  wire n_2234, n_2235, n_2236, n_2238, n_2240, n_2242, n_2243, n_2244;
  wire n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252;
  wire n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260;
  wire n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268;
  wire n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276;
  wire n_2277, n_2278, n_2279, n_2280, n_2281, n_2283, n_2285, n_2287;
  wire n_2288, n_2289, n_2290, n_2291, n_2292, n_2294, n_2296, n_2298;
  wire n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306;
  wire n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314;
  wire n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322;
  wire n_2323, n_2324, n_2325, n_2327, n_2329, n_2331, n_2332, n_2333;
  wire n_2334, n_2335, n_2336, n_2338, n_2340, n_2342, n_2343, n_2344;
  wire n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352;
  wire n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360;
  wire n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368;
  wire n_2369, n_2370, n_2371, n_2372, n_2373, n_2375, n_2377, n_2379;
  wire n_2380, n_2381, n_2382, n_2383, n_2384, n_2386, n_2388, n_2390;
  wire n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398;
  wire n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406;
  wire n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414;
  wire n_2415, n_2416, n_2417, n_2419, n_2421, n_2423, n_2424, n_2425;
  wire n_2426, n_2427, n_2428, n_2430, n_2432, n_2434, n_2435, n_2436;
  wire n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452;
  wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460;
  wire n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468;
  wire n_2469, n_2471, n_2473, n_2475, n_2476, n_2477, n_2478, n_2479;
  wire n_2480, n_2482, n_2484, n_2486, n_2487, n_2488, n_2489, n_2490;
  wire n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498;
  wire n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506;
  wire n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2515;
  wire n_2517, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2526;
  wire n_2528, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536;
  wire n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544;
  wire n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552;
  wire n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560;
  wire n_2561, n_2563, n_2565, n_2567, n_2568, n_2569, n_2570, n_2571;
  wire n_2572, n_2574, n_2576, n_2578, n_2579, n_2580, n_2581, n_2582;
  wire n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590;
  wire n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598;
  wire n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2607;
  wire n_2609, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2618;
  wire n_2620, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628;
  wire n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636;
  wire n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644;
  wire n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652;
  wire n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660;
  wire n_2661, n_2662, n_2663, n_2664, n_2665, n_2667, n_2669, n_2671;
  wire n_2672, n_2673, n_2674, n_2675, n_2676, n_2678, n_2680, n_2682;
  wire n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690;
  wire n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698;
  wire n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706;
  wire n_2707, n_2708, n_2709, n_2711, n_2713, n_2715, n_2716, n_2717;
  wire n_2718, n_2719, n_2720, n_2722, n_2724, n_2726, n_2727, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736;
  wire n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744;
  wire n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752;
  wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2759, n_2761, n_2763;
  wire n_2764, n_2765, n_2766, n_2767, n_2768, n_2770, n_2772, n_2774;
  wire n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782;
  wire n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790;
  wire n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798;
  wire n_2799, n_2800, n_2801, n_2803, n_2805, n_2807, n_2808, n_2809;
  wire n_2810, n_2811, n_2812, n_2814, n_2816, n_2818, n_2819, n_2820;
  wire n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828;
  wire n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836;
  wire n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844;
  wire n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852;
  wire n_2853, n_2855, n_2857, n_2859, n_2860, n_2861, n_2862, n_2863;
  wire n_2864, n_2866, n_2868, n_2870, n_2871, n_2872, n_2873, n_2874;
  wire n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882;
  wire n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890;
  wire n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2899;
  wire n_2901, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2910;
  wire n_2912, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920;
  wire n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928;
  wire n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936;
  wire n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944;
  wire n_2945, n_2947, n_2949, n_2951, n_2952, n_2953, n_2954, n_2955;
  wire n_2956, n_2958, n_2960, n_2962, n_2963, n_2964, n_2965, n_2966;
  wire n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974;
  wire n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982;
  wire n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2991;
  wire n_2993, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3002;
  wire n_3004, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012;
  wire n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020;
  wire n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028;
  wire n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036;
  wire n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044;
  wire n_3045, n_3047, n_3049, n_3051, n_3052, n_3053, n_3054, n_3055;
  wire n_3056, n_3058, n_3060, n_3062, n_3063, n_3064, n_3065, n_3066;
  wire n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074;
  wire n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082;
  wire n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3091;
  wire n_3093, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3102;
  wire n_3104, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112;
  wire n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120;
  wire n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128;
  wire n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136;
  wire n_3137, n_3139, n_3141, n_3143, n_3144, n_3145, n_3146, n_3147;
  wire n_3148, n_3150, n_3152, n_3154, n_3155, n_3156, n_3157, n_3158;
  wire n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166;
  wire n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174;
  wire n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3183;
  wire n_3185, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3194;
  wire n_3196, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204;
  wire n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212;
  wire n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220;
  wire n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228;
  wire n_3229, n_3230, n_3231, n_3232, n_3233, n_3235, n_3237, n_3239;
  wire n_3240, n_3241, n_3242, n_3243, n_3244, n_3246, n_3248, n_3250;
  wire n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258;
  wire n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266;
  wire n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274;
  wire n_3275, n_3276, n_3277, n_3279, n_3281, n_3283, n_3284, n_3285;
  wire n_3286, n_3287, n_3288, n_3290, n_3292, n_3294, n_3295, n_3296;
  wire n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304;
  wire n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312;
  wire n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320;
  wire n_3321, n_3322, n_3323, n_3324, n_3325, n_3327, n_3329, n_3331;
  wire n_3332, n_3333, n_3334, n_3335, n_3336, n_3338, n_3340, n_3342;
  wire n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350;
  wire n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358;
  wire n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366;
  wire n_3367, n_3368, n_3369, n_3371, n_3373, n_3375, n_3376, n_3377;
  wire n_3378, n_3379, n_3380, n_3382, n_3384, n_3386, n_3387, n_3388;
  wire n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396;
  wire n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404;
  wire n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, n_3412;
  wire n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, n_3420;
  wire n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428;
  wire n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436;
  wire n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444;
  wire n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452;
  wire n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460;
  wire n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468;
  wire n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476;
  wire n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484;
  wire n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492;
  wire n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500;
  wire n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508;
  wire n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516;
  wire n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524;
  wire n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532;
  wire n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540;
  wire n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548;
  wire n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556;
  wire n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564;
  wire n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572;
  wire n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580;
  wire n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588;
  wire n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596;
  wire n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604;
  wire n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612;
  wire n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620;
  wire n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628;
  wire n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636;
  wire n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644;
  wire n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652;
  wire n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660;
  wire n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668;
  wire n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676;
  wire n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684;
  wire n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692;
  wire n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700;
  wire n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708;
  wire n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716;
  wire n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724;
  wire n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732;
  wire n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740;
  wire n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748;
  wire n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756;
  wire n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764;
  wire n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772;
  wire n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780;
  wire n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788;
  wire n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796;
  wire n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804;
  wire n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812;
  wire n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820;
  wire n_3821, n_3822, n_3823, n_3826, n_3827, n_3828, n_3829, n_3831;
  wire n_3832, n_3833, n_3836, n_3837, n_3838, n_3839, n_3841, n_3842;
  wire n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850;
  wire n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858;
  wire n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866;
  wire n_3867, n_3870, n_3871, n_3872, n_3873, n_3875, n_3876, n_3877;
  wire n_3880, n_3881, n_3882, n_3883, n_3885, n_3886, n_3887, n_3888;
  wire n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896;
  wire n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904;
  wire n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912;
  wire n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920;
  wire n_3921, n_3922, n_3923, n_3924, n_3927, n_3928, n_3929, n_3930;
  wire n_3932, n_3933, n_3934, n_3937, n_3938, n_3939, n_3940, n_3942;
  wire n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950;
  wire n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958;
  wire n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966;
  wire n_3967, n_3968, n_3971, n_3972, n_3973, n_3974, n_3976, n_3977;
  wire n_3978, n_3981, n_3982, n_3983, n_3984, n_3986, n_3987, n_3988;
  wire n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996;
  wire n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004;
  wire n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012;
  wire n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020;
  wire n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028;
  wire n_4029, n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036;
  wire n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044;
  wire n_4045, n_4046, n_4048, n_4050, n_4052, n_4053, n_4054, n_4055;
  wire n_4056, n_4057, n_4059, n_4061, n_4063, n_4064, n_4065, n_4066;
  wire n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074;
  wire n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082;
  wire n_4083, n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090;
  wire n_4092, n_4094, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101;
  wire n_4103, n_4105, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112;
  wire n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120;
  wire n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128;
  wire n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136;
  wire n_4137, n_4138, n_4140, n_4142, n_4144, n_4145, n_4146, n_4147;
  wire n_4148, n_4149, n_4151, n_4153, n_4155, n_4156, n_4157, n_4158;
  wire n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166;
  wire n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174;
  wire n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182;
  wire n_4184, n_4186, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193;
  wire n_4195, n_4197, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204;
  wire n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212;
  wire n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220;
  wire n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, n_4228;
  wire n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236;
  wire n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244;
  wire n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252;
  wire n_4253, n_4254, n_4255, n_4256, n_4257, n_4258, n_4259, n_4260;
  wire n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, n_4268;
  wire n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276;
  wire n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284;
  wire n_4285, n_4286, n_4289, n_4290, n_4291, n_4292, n_4294, n_4295;
  wire n_4296, n_4299, n_4300, n_4301, n_4302, n_4304, n_4305, n_4306;
  wire n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313, n_4314;
  wire n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322;
  wire n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330;
  wire n_4333, n_4334, n_4335, n_4336, n_4338, n_4339, n_4340, n_4343;
  wire n_4344, n_4345, n_4346, n_4348, n_4349, n_4350, n_4351, n_4352;
  wire n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360;
  wire n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367, n_4368;
  wire n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375, n_4376;
  wire n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383, n_4384;
  wire n_4385, n_4386, n_4387, n_4390, n_4391, n_4392, n_4393, n_4395;
  wire n_4396, n_4397, n_4400, n_4401, n_4402, n_4403, n_4405, n_4406;
  wire n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413, n_4414;
  wire n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, n_4421, n_4422;
  wire n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430;
  wire n_4431, n_4434, n_4435, n_4436, n_4437, n_4439, n_4440, n_4441;
  wire n_4444, n_4445, n_4446, n_4447, n_4449, n_4450, n_4451, n_4452;
  wire n_4453, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460;
  wire n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4468;
  wire n_4469, n_4470, n_4471, n_4472, n_4473, n_4474, n_4475, n_4476;
  wire n_4477, n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484;
  wire n_4485, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492;
  wire n_4493, n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500;
  wire n_4501, n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508;
  wire n_4509, n_4511, n_4513, n_4515, n_4516, n_4517, n_4518, n_4519;
  wire n_4520, n_4522, n_4524, n_4526, n_4527, n_4528, n_4529, n_4530;
  wire n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, n_4537, n_4538;
  wire n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545, n_4546;
  wire n_4547, n_4548, n_4549, n_4550, n_4551, n_4552, n_4553, n_4556;
  wire n_4557, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4566;
  wire n_4568, n_4569, n_4570, n_4572, n_4573, n_4575, n_4576, n_4577;
  wire n_4578, n_4579, n_4580, n_4581, n_4582, n_4584, n_4586, n_4588;
  wire n_4589, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596;
  wire n_4597, n_4598, n_4599, n_4600, n_4601, n_4602, n_4603, n_4604;
  wire n_4605, n_4606, n_4607, n_4608, n_4609, n_4610, n_4611, n_4612;
  wire n_4613, n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620;
  wire n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628;
  wire n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636;
  wire n_4637, n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644;
  wire n_4645, n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652;
  wire n_4653, n_4654, n_4657, n_4658, n_4659, n_4660, n_4662, n_4663;
  wire n_4664, n_4667, n_4668, n_4669, n_4670, n_4672, n_4673, n_4674;
  wire n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681, n_4682;
  wire n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689, n_4690;
  wire n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697, n_4698;
  wire n_4701, n_4702, n_4703, n_4704, n_4706, n_4707, n_4708, n_4711;
  wire n_4712, n_4713, n_4714, n_4716, n_4717, n_4718, n_4719, n_4720;
  wire n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728;
  wire n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736;
  wire n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744;
  wire n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752;
  wire n_4753, n_4754, n_4755, n_4756, n_4757, n_4759, n_4761, n_4763;
  wire n_4764, n_4765, n_4766, n_4767, n_4768, n_4770, n_4772, n_4774;
  wire n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782;
  wire n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790;
  wire n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798;
  wire n_4799, n_4800, n_4801, n_4803, n_4805, n_4807, n_4808, n_4809;
  wire n_4810, n_4811, n_4812, n_4814, n_4816, n_4818, n_4819, n_4820;
  wire n_4821, n_4822, n_4823, n_4824, n_4825, n_4826, n_4827, n_4828;
  wire n_4829, n_4830, n_4831, n_4832, n_4833, n_4834, n_4835, n_4836;
  wire n_4837, n_4838, n_4839, n_4840, n_4841, n_4842, n_4843, n_4844;
  wire n_4845, n_4846, n_4847, n_4848, n_4849, n_4850, n_4851, n_4852;
  wire n_4853, n_4854, n_4855, n_4856, n_4857, n_4858, n_4859, n_4860;
  wire n_4861, n_4862, n_4863, n_4864, n_4865, n_4866, n_4867, n_4868;
  wire n_4869, n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876;
  wire n_4877, n_4880, n_4881, n_4882, n_4883, n_4885, n_4886, n_4887;
  wire n_4890, n_4891, n_4892, n_4893, n_4895, n_4896, n_4897, n_4898;
  wire n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, n_4906;
  wire n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914;
  wire n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4924;
  wire n_4925, n_4926, n_4927, n_4929, n_4930, n_4931, n_4934, n_4935;
  wire n_4936, n_4937, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944;
  wire n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952;
  wire n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960;
  wire n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968;
  wire n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976;
  wire n_4977, n_4978, n_4981, n_4982, n_4983, n_4984, n_4986, n_4987;
  wire n_4988, n_4991, n_4992, n_4993, n_4994, n_4996, n_4997, n_4998;
  wire n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, n_5005, n_5006;
  wire n_5007, n_5008, n_5009, n_5010, n_5011, n_5012, n_5013, n_5014;
  wire n_5015, n_5016, n_5017, n_5018, n_5019, n_5020, n_5021, n_5022;
  wire n_5025, n_5026, n_5027, n_5028, n_5030, n_5031, n_5032, n_5035;
  wire n_5036, n_5037, n_5038, n_5040, n_5041, n_5042, n_5043, n_5044;
  wire n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051, n_5052;
  wire n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059, n_5060;
  wire n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, n_5068;
  wire n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076;
  wire n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084;
  wire n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092;
  wire n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099, n_5100;
  wire n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108;
  wire n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116;
  wire n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124;
  wire n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132;
  wire n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, n_5140;
  wire n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147, n_5148;
  wire n_5149, n_5150, n_5151, n_5153, n_5155, n_5157, n_5158, n_5159;
  wire n_5160, n_5161, n_5162, n_5164, n_5166, n_5168, n_5169, n_5170;
  wire n_5171, n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178;
  wire n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186;
  wire n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194;
  wire n_5195, n_5197, n_5199, n_5201, n_5202, n_5203, n_5204, n_5205;
  wire n_5206, n_5208, n_5210, n_5212, n_5213, n_5214, n_5215, n_5216;
  wire n_5217, n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224;
  wire n_5225, n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232;
  wire n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240;
  wire n_5241, n_5242, n_5243, n_5245, n_5247, n_5249, n_5250, n_5251;
  wire n_5252, n_5253, n_5254, n_5256, n_5258, n_5260, n_5261, n_5262;
  wire n_5263, n_5264, n_5265, n_5266, n_5267, n_5268, n_5269, n_5270;
  wire n_5271, n_5272, n_5273, n_5274, n_5275, n_5276, n_5277, n_5278;
  wire n_5279, n_5280, n_5281, n_5282, n_5283, n_5284, n_5285, n_5286;
  wire n_5287, n_5289, n_5291, n_5293, n_5294, n_5295, n_5296, n_5297;
  wire n_5298, n_5300, n_5302, n_5304, n_5305, n_5306, n_5307, n_5308;
  wire n_5309, n_5310, n_5311, n_5312, n_5313, n_5314, n_5315, n_5316;
  wire n_5317, n_5318, n_5319, n_5320, n_5321, n_5322, n_5323, n_5324;
  wire n_5325, n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5332;
  wire n_5333, n_5334, n_5335, n_5336, n_5337, n_5338, n_5339, n_5341;
  wire n_5343, n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5352;
  wire n_5354, n_5356, n_5357, n_5358, n_5359, n_5360, n_5361, n_5362;
  wire n_5363, n_5364, n_5365, n_5366, n_5367, n_5368, n_5369, n_5370;
  wire n_5371, n_5372, n_5373, n_5374, n_5375, n_5376, n_5377, n_5378;
  wire n_5379, n_5380, n_5381, n_5382, n_5383, n_5385, n_5387, n_5389;
  wire n_5390, n_5391, n_5392, n_5393, n_5394, n_5396, n_5398, n_5400;
  wire n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408;
  wire n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416;
  wire n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424;
  wire n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5433;
  wire n_5435, n_5437, n_5438, n_5439, n_5440, n_5441, n_5442, n_5444;
  wire n_5446, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453, n_5454;
  wire n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462;
  wire n_5463, n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470;
  wire n_5471, n_5472, n_5473, n_5474, n_5475, n_5477, n_5479, n_5481;
  wire n_5482, n_5483, n_5484, n_5485, n_5486, n_5488, n_5490, n_5492;
  wire n_5493, n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, n_5500;
  wire n_5501, n_5502, n_5503, n_5504, n_5505, n_5506, n_5507, n_5508;
  wire n_5509, n_5510, n_5511, n_5512, n_5513, n_5514, n_5515, n_5516;
  wire n_5517, n_5518, n_5519, n_5520, n_5521, n_5522, n_5523, n_5524;
  wire n_5525, n_5526, n_5527, n_5528, n_5529, n_5530, n_5531, n_5533;
  wire n_5535, n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5544;
  wire n_5546, n_5548, n_5549, n_5550, n_5551, n_5552, n_5553, n_5554;
  wire n_5555, n_5556, n_5557, n_5558, n_5559, n_5560, n_5561, n_5562;
  wire n_5563, n_5564, n_5565, n_5566, n_5567, n_5568, n_5569, n_5570;
  wire n_5571, n_5572, n_5573, n_5574, n_5575, n_5577, n_5579, n_5581;
  wire n_5582, n_5583, n_5584, n_5585, n_5586, n_5588, n_5590, n_5592;
  wire n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600;
  wire n_5601, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608;
  wire n_5609, n_5610, n_5611, n_5612, n_5613, n_5614, n_5615, n_5616;
  wire n_5617, n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5625;
  wire n_5627, n_5629, n_5630, n_5631, n_5632, n_5633, n_5634, n_5636;
  wire n_5638, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645, n_5646;
  wire n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653, n_5654;
  wire n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661, n_5662;
  wire n_5663, n_5664, n_5665, n_5666, n_5667, n_5669, n_5671, n_5673;
  wire n_5674, n_5675, n_5676, n_5677, n_5678, n_5680, n_5682, n_5684;
  wire n_5685, n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692;
  wire n_5693, n_5694, n_5695, n_5696, n_5697, n_5698, n_5699, n_5700;
  wire n_5701, n_5702, n_5703, n_5704, n_5705, n_5706, n_5707, n_5708;
  wire n_5709, n_5710, n_5711, n_5712, n_5713, n_5714, n_5715, n_5716;
  wire n_5717, n_5718, n_5719, n_5721, n_5723, n_5725, n_5726, n_5727;
  wire n_5728, n_5729, n_5730, n_5732, n_5734, n_5736, n_5737, n_5738;
  wire n_5739, n_5740, n_5741, n_5742, n_5743, n_5744, n_5745, n_5746;
  wire n_5747, n_5748, n_5749, n_5750, n_5751, n_5752, n_5753, n_5754;
  wire n_5755, n_5756, n_5757, n_5758, n_5759, n_5760, n_5761, n_5762;
  wire n_5763, n_5765, n_5767, n_5769, n_5770, n_5771, n_5772, n_5773;
  wire n_5774, n_5776, n_5778, n_5780, n_5781, n_5782, n_5783, n_5784;
  wire n_5785, n_5786, n_5787, n_5788, n_5789, n_5790, n_5791, n_5792;
  wire n_5793, n_5794, n_5795, n_5796, n_5797, n_5798, n_5799, n_5800;
  wire n_5801, n_5802, n_5803, n_5804, n_5805, n_5806, n_5807, n_5808;
  wire n_5809, n_5810, n_5811, n_5813, n_5815, n_5817, n_5818, n_5819;
  wire n_5820, n_5821, n_5822, n_5824, n_5826, n_5828, n_5829, n_5830;
  wire n_5831, n_5832, n_5833, n_5834, n_5835, n_5836, n_5837, n_5838;
  wire n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845, n_5846;
  wire n_5847, n_5848, n_5849, n_5850, n_5851, n_5852, n_5853, n_5854;
  wire n_5855, n_5857, n_5859, n_5861, n_5862, n_5863, n_5864, n_5865;
  wire n_5866, n_5868, n_5870, n_5872, n_5873, n_5874, n_5875, n_5876;
  wire n_5877, n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884;
  wire n_5885, n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892;
  wire n_5893, n_5894, n_5895, n_5896, n_5897, n_5898, n_5899, n_5900;
  wire n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907, n_5908;
  wire n_5909, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915, n_5916;
  wire n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923, n_5924;
  wire n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932;
  wire n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940;
  wire n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947, n_5948;
  wire n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956;
  wire n_5957, n_5958, n_5959, n_5960, n_5961, n_5962, n_5963, n_5964;
  wire n_5965, n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972;
  wire n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5980;
  wire n_5981, n_5982, n_5983, n_5984, n_5985, n_5986, n_5987, n_5988;
  wire n_5989, n_5990, n_5991, n_5992, n_5993, n_5994, n_5995, n_5996;
  wire n_5997, n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004;
  wire n_6005, n_6006, n_6007, n_6008, n_6009, n_6010, n_6011, n_6012;
  wire n_6013, n_6014, n_6015, n_6016, n_6017, n_6018, n_6019, n_6020;
  wire n_6021, n_6022, n_6023, n_6024, n_6025, n_6026, n_6027, n_6028;
  wire n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035, n_6036;
  wire n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044;
  wire n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051, n_6052;
  wire n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059, n_6060;
  wire n_6061, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067, n_6068;
  wire n_6069, n_6070, n_6071, n_6072, n_6073, n_6074, n_6075, n_6076;
  wire n_6077, n_6078, n_6079, n_6080, n_6081, n_6082, n_6083, n_6084;
  wire n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091, n_6092;
  wire n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099, n_6100;
  wire n_6101, n_6102, n_6103, n_6104, n_6105, n_6106, n_6107, n_6108;
  wire n_6109, n_6110, n_6111, n_6114, n_6115, n_6116, n_6117, n_6119;
  wire n_6120, n_6121, n_6124, n_6125, n_6126, n_6127, n_6129, n_6130;
  wire n_6131, n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138;
  wire n_6139, n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6146;
  wire n_6147, n_6148, n_6149, n_6150, n_6151, n_6152, n_6153, n_6154;
  wire n_6155, n_6158, n_6159, n_6160, n_6161, n_6163, n_6164, n_6165;
  wire n_6168, n_6169, n_6170, n_6171, n_6173, n_6174, n_6175, n_6176;
  wire n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184;
  wire n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192;
  wire n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6200;
  wire n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207, n_6208;
  wire n_6209, n_6210, n_6211, n_6212, n_6215, n_6216, n_6217, n_6218;
  wire n_6220, n_6221, n_6222, n_6225, n_6226, n_6227, n_6228, n_6230;
  wire n_6231, n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238;
  wire n_6239, n_6240, n_6241, n_6242, n_6243, n_6244, n_6245, n_6246;
  wire n_6247, n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254;
  wire n_6255, n_6256, n_6259, n_6260, n_6261, n_6262, n_6264, n_6265;
  wire n_6266, n_6269, n_6270, n_6271, n_6272, n_6274, n_6275, n_6276;
  wire n_6277, n_6278, n_6279, n_6280, n_6281, n_6282, n_6283, n_6284;
  wire n_6285, n_6286, n_6287, n_6288, n_6289, n_6290, n_6291, n_6292;
  wire n_6293, n_6294, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300;
  wire n_6301, n_6302, n_6303, n_6304, n_6305, n_6306, n_6307, n_6308;
  wire n_6309, n_6310, n_6311, n_6312, n_6313, n_6314, n_6315, n_6316;
  wire n_6317, n_6318, n_6319, n_6320, n_6321, n_6322, n_6323, n_6324;
  wire n_6325, n_6326, n_6327, n_6328, n_6329, n_6330, n_6331, n_6332;
  wire n_6333, n_6334, n_6336, n_6338, n_6340, n_6341, n_6342, n_6343;
  wire n_6344, n_6345, n_6347, n_6349, n_6351, n_6352, n_6353, n_6354;
  wire n_6355, n_6356, n_6357, n_6358, n_6359, n_6360, n_6361, n_6362;
  wire n_6363, n_6364, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370;
  wire n_6371, n_6372, n_6373, n_6374, n_6375, n_6376, n_6377, n_6378;
  wire n_6380, n_6382, n_6384, n_6385, n_6386, n_6387, n_6388, n_6389;
  wire n_6391, n_6393, n_6395, n_6396, n_6397, n_6398, n_6399, n_6400;
  wire n_6401, n_6402, n_6403, n_6404, n_6405, n_6406, n_6407, n_6408;
  wire n_6409, n_6410, n_6411, n_6412, n_6413, n_6414, n_6415, n_6416;
  wire n_6417, n_6418, n_6419, n_6420, n_6421, n_6422, n_6423, n_6424;
  wire n_6425, n_6426, n_6428, n_6430, n_6432, n_6433, n_6434, n_6435;
  wire n_6436, n_6437, n_6439, n_6441, n_6443, n_6444, n_6445, n_6446;
  wire n_6447, n_6448, n_6449, n_6450, n_6451, n_6452, n_6453, n_6454;
  wire n_6455, n_6456, n_6457, n_6458, n_6459, n_6460, n_6461, n_6462;
  wire n_6463, n_6464, n_6465, n_6466, n_6467, n_6468, n_6469, n_6470;
  wire n_6472, n_6474, n_6476, n_6477, n_6478, n_6479, n_6480, n_6481;
  wire n_6483, n_6485, n_6487, n_6488, n_6489, n_6490, n_6491, n_6492;
  wire n_6493, n_6494, n_6495, n_6496, n_6497, n_6498, n_6499, n_6500;
  wire n_6501, n_6502, n_6503, n_6504, n_6505, n_6506, n_6507, n_6508;
  wire n_6509, n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6516;
  wire n_6517, n_6518, n_6519, n_6520, n_6521, n_6522, n_6523, n_6524;
  wire n_6525, n_6526, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532;
  wire n_6533, n_6534, n_6535, n_6536, n_6537, n_6538, n_6539, n_6540;
  wire n_6541, n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548;
  wire n_6549, n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556;
  wire n_6557, n_6558, n_6559, n_6560, n_6561, n_6562, n_6563, n_6564;
  wire n_6565, n_6566, n_6567, n_6568, n_6569, n_6570, n_6571, n_6572;
  wire n_6573, n_6574, n_6577, n_6578, n_6579, n_6580, n_6582, n_6583;
  wire n_6584, n_6587, n_6588, n_6589, n_6590, n_6592, n_6593, n_6594;
  wire n_6595, n_6596, n_6597, n_6598, n_6599, n_6600, n_6601, n_6602;
  wire n_6603, n_6604, n_6605, n_6606, n_6607, n_6608, n_6609, n_6610;
  wire n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617, n_6618;
  wire n_6621, n_6622, n_6623, n_6624, n_6626, n_6627, n_6628, n_6631;
  wire n_6632, n_6633, n_6634, n_6636, n_6637, n_6638, n_6639, n_6640;
  wire n_6641, n_6642, n_6643, n_6644, n_6645, n_6646, n_6647, n_6648;
  wire n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655, n_6656;
  wire n_6657, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663, n_6664;
  wire n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671, n_6672;
  wire n_6673, n_6674, n_6675, n_6676, n_6677, n_6679, n_6681, n_6683;
  wire n_6684, n_6685, n_6686, n_6687, n_6688, n_6690, n_6692, n_6694;
  wire n_6695, n_6696, n_6697, n_6698, n_6699, n_6700, n_6701, n_6702;
  wire n_6703, n_6704, n_6705, n_6706, n_6707, n_6708, n_6709, n_6710;
  wire n_6711, n_6712, n_6713, n_6714, n_6715, n_6716, n_6717, n_6718;
  wire n_6719, n_6720, n_6721, n_6723, n_6725, n_6727, n_6728, n_6729;
  wire n_6730, n_6731, n_6732, n_6734, n_6736, n_6738, n_6739, n_6740;
  wire n_6741, n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748;
  wire n_6749, n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756;
  wire n_6757, n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764;
  wire n_6765, n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772;
  wire n_6773, n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780;
  wire n_6781, n_6782, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788;
  wire n_6789, n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796;
  wire n_6797, n_6800, n_6801, n_6802, n_6803, n_6805, n_6806, n_6807;
  wire n_6810, n_6811, n_6812, n_6813, n_6815, n_6816, n_6817, n_6818;
  wire n_6819, n_6820, n_6821, n_6822, n_6823, n_6824, n_6825, n_6826;
  wire n_6827, n_6828, n_6829, n_6830, n_6831, n_6832, n_6833, n_6834;
  wire n_6835, n_6836, n_6837, n_6838, n_6839, n_6840, n_6841, n_6844;
  wire n_6845, n_6846, n_6847, n_6849, n_6850, n_6851, n_6854, n_6855;
  wire n_6856, n_6857, n_6859, n_6860, n_6861, n_6862, n_6863, n_6864;
  wire n_6865, n_6866, n_6867, n_6868, n_6869, n_6870, n_6871, n_6872;
  wire n_6873, n_6874, n_6875, n_6876, n_6877, n_6878, n_6879, n_6880;
  wire n_6881, n_6882, n_6883, n_6884, n_6885, n_6886, n_6887, n_6888;
  wire n_6889, n_6890, n_6891, n_6892, n_6893, n_6894, n_6895, n_6896;
  wire n_6897, n_6898, n_6901, n_6902, n_6903, n_6904, n_6906, n_6907;
  wire n_6908, n_6911, n_6912, n_6913, n_6914, n_6916, n_6917, n_6918;
  wire n_6919, n_6920, n_6921, n_6922, n_6923, n_6924, n_6925, n_6926;
  wire n_6927, n_6928, n_6929, n_6930, n_6931, n_6932, n_6933, n_6934;
  wire n_6935, n_6936, n_6937, n_6938, n_6939, n_6940, n_6941, n_6942;
  wire n_6945, n_6946, n_6947, n_6948, n_6950, n_6951, n_6952, n_6955;
  wire n_6956, n_6957, n_6958, n_6960, n_6961, n_6962, n_6963, n_6964;
  wire n_6965, n_6966, n_6967, n_6968, n_6969, n_6970, n_6971, n_6972;
  wire n_6973, n_6974, n_6975, n_6976, n_6977, n_6978, n_6979, n_6980;
  wire n_6981, n_6982, n_6983, n_6984, n_6985, n_6986, n_6987, n_6988;
  wire n_6989, n_6990, n_6991, n_6992, n_6993, n_6994, n_6995, n_6996;
  wire n_6997, n_6998, n_6999, n_7000, n_7001, n_7002, n_7003, n_7004;
  wire n_7005, n_7006, n_7007, n_7008, n_7009, n_7010, n_7011, n_7012;
  wire n_7013, n_7014, n_7015, n_7016, n_7017, n_7018, n_7019, n_7020;
  wire n_7021, n_7022, n_7023, n_7024, n_7025, n_7026, n_7027, n_7028;
  wire n_7029, n_7030, n_7031, n_7032, n_7033, n_7034, n_7035, n_7036;
  wire n_7037, n_7038, n_7039, n_7040, n_7041, n_7042, n_7043, n_7044;
  wire n_7045, n_7046, n_7047, n_7048, n_7049, n_7050, n_7051, n_7052;
  wire n_7053, n_7054, n_7056, n_7058, n_7060, n_7061, n_7062, n_7063;
  wire n_7064, n_7065, n_7067, n_7069, n_7071, n_7072, n_7073, n_7074;
  wire n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081, n_7082;
  wire n_7083, n_7084, n_7085, n_7086, n_7087, n_7088, n_7089, n_7090;
  wire n_7091, n_7092, n_7093, n_7094, n_7095, n_7096, n_7097, n_7098;
  wire n_7100, n_7102, n_7104, n_7105, n_7106, n_7107, n_7108, n_7109;
  wire n_7111, n_7113, n_7115, n_7116, n_7117, n_7118, n_7119, n_7120;
  wire n_7121, n_7122, n_7123, n_7124, n_7125, n_7126, n_7127, n_7128;
  wire n_7129, n_7130, n_7131, n_7132, n_7133, n_7134, n_7135, n_7136;
  wire n_7137, n_7138, n_7139, n_7140, n_7141, n_7142, n_7143, n_7144;
  wire n_7145, n_7146, n_7148, n_7150, n_7152, n_7153, n_7154, n_7155;
  wire n_7156, n_7157, n_7159, n_7161, n_7163, n_7164, n_7165, n_7166;
  wire n_7167, n_7168, n_7169, n_7170, n_7171, n_7172, n_7173, n_7174;
  wire n_7175, n_7176, n_7177, n_7178, n_7179, n_7180, n_7181, n_7182;
  wire n_7183, n_7184, n_7185, n_7186, n_7187, n_7188, n_7189, n_7190;
  wire n_7192, n_7194, n_7196, n_7197, n_7198, n_7199, n_7200, n_7201;
  wire n_7203, n_7205, n_7207, n_7208, n_7209, n_7210, n_7211, n_7212;
  wire n_7213, n_7214, n_7215, n_7216, n_7217, n_7218, n_7219, n_7220;
  wire n_7221, n_7222, n_7223, n_7224, n_7225, n_7226, n_7227, n_7228;
  wire n_7229, n_7230, n_7231, n_7232, n_7233, n_7234, n_7235, n_7236;
  wire n_7237, n_7238, n_7239, n_7240, n_7241, n_7242, n_7244, n_7246;
  wire n_7248, n_7249, n_7250, n_7251, n_7252, n_7253, n_7255, n_7257;
  wire n_7259, n_7260, n_7261, n_7262, n_7263, n_7264, n_7265, n_7266;
  wire n_7267, n_7268, n_7269, n_7270, n_7271, n_7272, n_7273, n_7274;
  wire n_7275, n_7276, n_7277, n_7278, n_7279, n_7280, n_7281, n_7282;
  wire n_7283, n_7284, n_7285, n_7286, n_7288, n_7290, n_7292, n_7293;
  wire n_7294, n_7295, n_7296, n_7297, n_7299, n_7301, n_7303, n_7304;
  wire n_7305, n_7306, n_7307, n_7308, n_7309, n_7310, n_7311, n_7312;
  wire n_7313, n_7314, n_7315, n_7316, n_7317, n_7318, n_7319, n_7320;
  wire n_7321, n_7322, n_7323, n_7324, n_7325, n_7326, n_7327, n_7328;
  wire n_7329, n_7330, n_7331, n_7332, n_7333, n_7334, n_7336, n_7338;
  wire n_7340, n_7341, n_7342, n_7343, n_7344, n_7345, n_7347, n_7349;
  wire n_7351, n_7352, n_7353, n_7354, n_7355, n_7356, n_7357, n_7358;
  wire n_7359, n_7360, n_7361, n_7362, n_7363, n_7364, n_7365, n_7366;
  wire n_7367, n_7368, n_7369, n_7370, n_7371, n_7372, n_7373, n_7374;
  wire n_7375, n_7376, n_7377, n_7378, n_7380, n_7382, n_7384, n_7385;
  wire n_7386, n_7387, n_7388, n_7389, n_7391, n_7393, n_7395, n_7396;
  wire n_7397, n_7398, n_7399, n_7400, n_7401, n_7402, n_7403, n_7404;
  wire n_7405, n_7406, n_7407, n_7408, n_7409, n_7410, n_7411, n_7412;
  wire n_7413, n_7414, n_7415, n_7416, n_7417, n_7418, n_7419, n_7420;
  wire n_7421, n_7422, n_7423, n_7424, n_7425, n_7426, n_7427, n_7428;
  wire n_7429, n_7430, n_7431, n_7432, n_7433, n_7434, n_7436, n_7438;
  wire n_7440, n_7441, n_7442, n_7443, n_7444, n_7445, n_7447, n_7449;
  wire n_7451, n_7452, n_7453, n_7454, n_7455, n_7456, n_7457, n_7458;
  wire n_7459, n_7460, n_7461, n_7462, n_7463, n_7464, n_7465, n_7466;
  wire n_7467, n_7468, n_7469, n_7470, n_7471, n_7472, n_7473, n_7474;
  wire n_7475, n_7476, n_7477, n_7478, n_7480, n_7482, n_7484, n_7485;
  wire n_7486, n_7487, n_7488, n_7489, n_7491, n_7493, n_7495, n_7496;
  wire n_7497, n_7498, n_7499, n_7500, n_7501, n_7502, n_7503, n_7504;
  wire n_7505, n_7506, n_7507, n_7508, n_7509, n_7510, n_7511, n_7512;
  wire n_7513, n_7514, n_7515, n_7516, n_7517, n_7518, n_7519, n_7520;
  wire n_7521, n_7522, n_7523, n_7524, n_7525, n_7526, n_7528, n_7530;
  wire n_7532, n_7533, n_7534, n_7535, n_7536, n_7537, n_7539, n_7541;
  wire n_7543, n_7544, n_7545, n_7546, n_7547, n_7548, n_7549, n_7550;
  wire n_7551, n_7552, n_7553, n_7554, n_7555, n_7556, n_7557, n_7558;
  wire n_7559, n_7560, n_7561, n_7562, n_7563, n_7564, n_7565, n_7566;
  wire n_7567, n_7568, n_7569, n_7570, n_7572, n_7574, n_7576, n_7577;
  wire n_7578, n_7579, n_7580, n_7581, n_7583, n_7585, n_7587, n_7588;
  wire n_7589, n_7590, n_7591, n_7592, n_7593, n_7594, n_7595, n_7596;
  wire n_7597, n_7598, n_7599, n_7600, n_7601, n_7602, n_7603, n_7604;
  wire n_7605, n_7606, n_7607, n_7608, n_7609, n_7610, n_7611, n_7612;
  wire n_7613, n_7614, n_7615, n_7616, n_7617, n_7618, n_7619, n_7620;
  wire n_7621, n_7622, n_7624, n_7626, n_7628, n_7629, n_7630, n_7631;
  wire n_7632, n_7633, n_7635, n_7637, n_7639, n_7640, n_7641, n_7642;
  wire n_7643, n_7644, n_7645, n_7646, n_7647, n_7648, n_7649, n_7650;
  wire n_7651, n_7652, n_7653, n_7654, n_7655, n_7656, n_7657, n_7658;
  wire n_7659, n_7660, n_7661, n_7662, n_7663, n_7664, n_7665, n_7666;
  wire n_7668, n_7670, n_7672, n_7673, n_7674, n_7675, n_7676, n_7677;
  wire n_7679, n_7681, n_7683, n_7684, n_7685, n_7686, n_7687, n_7688;
  wire n_7689, n_7690, n_7691, n_7692, n_7693, n_7694, n_7695, n_7696;
  wire n_7697, n_7698, n_7699, n_7700, n_7701, n_7702, n_7703, n_7704;
  wire n_7705, n_7706, n_7707, n_7708, n_7709, n_7710, n_7711, n_7712;
  wire n_7713, n_7714, n_7716, n_7718, n_7720, n_7721, n_7722, n_7723;
  wire n_7724, n_7725, n_7727, n_7729, n_7731, n_7732, n_7733, n_7734;
  wire n_7735, n_7736, n_7737, n_7738, n_7739, n_7740, n_7741, n_7742;
  wire n_7743, n_7744, n_7745, n_7746, n_7747, n_7748, n_7749, n_7750;
  wire n_7751, n_7752, n_7753, n_7754, n_7755, n_7756, n_7757, n_7758;
  wire n_7760, n_7762, n_7764, n_7765, n_7766, n_7767, n_7768, n_7769;
  wire n_7771, n_7773, n_7775, n_7776, n_7777, n_7778, n_7779, n_7780;
  wire n_7781, n_7782, n_7783, n_7784, n_7785, n_7786, n_7787, n_7788;
  wire n_7789, n_7790, n_7791, n_7792, n_7793, n_7794, n_7795, n_7796;
  wire n_7797, n_7798, n_7799, n_7800, n_7801, n_7802, n_7803, n_7804;
  wire n_7805, n_7806, n_7807, n_7808, n_7809, n_7810, n_7811, n_7812;
  wire n_7813, n_7814, n_7815, n_7816, n_7817, n_7818, n_7819, n_7820;
  wire n_7821, n_7822, n_7823, n_7824, n_7825, n_7826, n_7827, n_7828;
  wire n_7829, n_7830, n_7831, n_7832, n_7833, n_7834, n_7835, n_7836;
  wire n_7837, n_7838, n_7839, n_7840, n_7841, n_7842, n_7843, n_7844;
  wire n_7845, n_7846, n_7847, n_7848, n_7849, n_7850, n_7851, n_7852;
  wire n_7853, n_7854, n_7855, n_7856, n_7857, n_7858, n_7859, n_7860;
  wire n_7861, n_7862, n_7863, n_7864, n_7865, n_7866, n_7867, n_7868;
  wire n_7869, n_7870, n_7871, n_7872, n_7873, n_7874, n_7875, n_7876;
  wire n_7877, n_7878, n_7879, n_7880, n_7881, n_7882, n_7883, n_7884;
  wire n_7885, n_7886, n_7887, n_7888, n_7889, n_7890, n_7891, n_7892;
  wire n_7893, n_7894, n_7895, n_7896, n_7897, n_7898, n_7899, n_7900;
  wire n_7901, n_7902, n_7903, n_7904, n_7905, n_7906, n_7907, n_7908;
  wire n_7909, n_7910, n_7911, n_7912, n_7913, n_7914, n_7915, n_7916;
  wire n_7917, n_7918, n_7919, n_7920, n_7921, n_7922, n_7923, n_7924;
  wire n_7925, n_7926, n_7927, n_7928, n_7929, n_7930, n_7931, n_7932;
  wire n_7933, n_7934, n_7935, n_7936, n_7937, n_7938, n_7939, n_7940;
  wire n_7941, n_7942, n_7943, n_7944, n_7945, n_7946, n_7947, n_7948;
  wire n_7949, n_7950, n_7951, n_7952, n_7953, n_7954, n_7955, n_7956;
  wire n_7957, n_7958, n_7959, n_7960, n_7961, n_7962, n_7963, n_7964;
  wire n_7965, n_7966, n_7967, n_7968, n_7969, n_7970, n_7971, n_7972;
  wire n_7973, n_7974, n_7975, n_7976, n_7977, n_7978, n_7979, n_7980;
  wire n_7981, n_7982, n_7983, n_7984, n_7985, n_7986, n_7987, n_7988;
  wire n_7989, n_7990, n_7991, n_7992, n_7993, n_7994, n_7995, n_7996;
  wire n_7997, n_7998, n_7999, n_8000, n_8001, n_8002, n_8003, n_8004;
  wire n_8005, n_8006, n_8007, n_8008, n_8009, n_8010, n_8011, n_8012;
  wire n_8013, n_8014, n_8017, n_8018, n_8019, n_8020, n_8022, n_8023;
  wire n_8024, n_8027, n_8028, n_8029, n_8030, n_8032, n_8033, n_8034;
  wire n_8035, n_8036, n_8037, n_8038, n_8039, n_8040, n_8041, n_8042;
  wire n_8043, n_8044, n_8045, n_8046, n_8047, n_8048, n_8049, n_8050;
  wire n_8051, n_8052, n_8053, n_8054, n_8055, n_8056, n_8057, n_8058;
  wire n_8061, n_8062, n_8063, n_8064, n_8066, n_8067, n_8068, n_8071;
  wire n_8072, n_8073, n_8074, n_8076, n_8077, n_8078, n_8079, n_8080;
  wire n_8081, n_8082, n_8083, n_8084, n_8085, n_8086, n_8087, n_8088;
  wire n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095, n_8096;
  wire n_8097, n_8098, n_8099, n_8100, n_8101, n_8102, n_8103, n_8104;
  wire n_8105, n_8106, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112;
  wire n_8113, n_8114, n_8115, n_8116, n_8117, n_8119, n_8121, n_8123;
  wire n_8124, n_8125, n_8126, n_8127, n_8128, n_8130, n_8132, n_8134;
  wire n_8135, n_8136, n_8137, n_8138, n_8139, n_8140, n_8141, n_8142;
  wire n_8143, n_8144, n_8145, n_8146, n_8147, n_8148, n_8149, n_8150;
  wire n_8151, n_8152, n_8153, n_8154, n_8155, n_8156, n_8157, n_8158;
  wire n_8159, n_8160, n_8161, n_8163, n_8165, n_8167, n_8168, n_8169;
  wire n_8170, n_8171, n_8172, n_8174, n_8176, n_8178, n_8179, n_8180;
  wire n_8181, n_8182, n_8183, n_8184, n_8185, n_8186, n_8187, n_8188;
  wire n_8189, n_8190, n_8191, n_8192, n_8193, n_8194, n_8195, n_8196;
  wire n_8197, n_8198, n_8199, n_8200, n_8201, n_8202, n_8203, n_8204;
  wire n_8205, n_8206, n_8207, n_8208, n_8209, n_8210, n_8211, n_8212;
  wire n_8213, n_8214, n_8215, n_8216, n_8217, n_8218, n_8219, n_8220;
  wire n_8221, n_8222, n_8223, n_8224, n_8225, n_8226, n_8227, n_8228;
  wire n_8229, n_8230, n_8231, n_8232, n_8233, n_8234, n_8235, n_8236;
  wire n_8237, n_8240, n_8241, n_8242, n_8243, n_8245, n_8246, n_8247;
  wire n_8250, n_8251, n_8252, n_8253, n_8255, n_8256, n_8257, n_8258;
  wire n_8259, n_8260, n_8261, n_8262, n_8263, n_8264, n_8265, n_8266;
  wire n_8267, n_8268, n_8269, n_8270, n_8271, n_8272, n_8273, n_8274;
  wire n_8275, n_8276, n_8277, n_8278, n_8279, n_8280, n_8281, n_8284;
  wire n_8285, n_8286, n_8287, n_8289, n_8290, n_8291, n_8294, n_8295;
  wire n_8296, n_8297, n_8299, n_8300, n_8301, n_8302, n_8303, n_8304;
  wire n_8305, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311, n_8312;
  wire n_8313, n_8314, n_8315, n_8316, n_8317, n_8318, n_8319, n_8320;
  wire n_8321, n_8322, n_8323, n_8324, n_8325, n_8326, n_8327, n_8328;
  wire n_8329, n_8330, n_8331, n_8332, n_8333, n_8334, n_8335, n_8336;
  wire n_8337, n_8338, n_8341, n_8342, n_8343, n_8344, n_8346, n_8347;
  wire n_8348, n_8351, n_8352, n_8353, n_8354, n_8356, n_8357, n_8358;
  wire n_8359, n_8360, n_8361, n_8362, n_8363, n_8364, n_8365, n_8366;
  wire n_8367, n_8368, n_8369, n_8370, n_8371, n_8372, n_8373, n_8374;
  wire n_8375, n_8376, n_8377, n_8378, n_8379, n_8380, n_8381, n_8382;
  wire n_8385, n_8386, n_8387, n_8388, n_8390, n_8391, n_8392, n_8395;
  wire n_8396, n_8397, n_8398, n_8400, n_8401, n_8402, n_8403, n_8404;
  wire n_8405, n_8406, n_8407, n_8408, n_8409, n_8410, n_8411, n_8412;
  wire n_8413, n_8414, n_8415, n_8416, n_8417, n_8418, n_8419, n_8420;
  wire n_8421, n_8422, n_8423, n_8424, n_8425, n_8426, n_8427, n_8428;
  wire n_8429, n_8430, n_8431, n_8432, n_8433, n_8434, n_8435, n_8436;
  wire n_8437, n_8438, n_8439, n_8440, n_8441, n_8442, n_8443, n_8444;
  wire n_8445, n_8446, n_8447, n_8448, n_8449, n_8450, n_8451, n_8452;
  wire n_8453, n_8454, n_8455, n_8456, n_8457, n_8458, n_8459, n_8460;
  wire n_8461, n_8462, n_8463, n_8464, n_8465, n_8466, n_8467, n_8468;
  wire n_8469, n_8470, n_8471, n_8472, n_8473, n_8474, n_8475, n_8476;
  wire n_8477, n_8479, n_8481, n_8483, n_8484, n_8485, n_8486, n_8487;
  wire n_8488, n_8490, n_8492, n_8494, n_8495, n_8496, n_8497, n_8498;
  wire n_8499, n_8500, n_8501, n_8502, n_8503, n_8504, n_8505, n_8506;
  wire n_8507, n_8508, n_8509, n_8510, n_8511, n_8512, n_8513, n_8514;
  wire n_8515, n_8516, n_8517, n_8518, n_8519, n_8520, n_8521, n_8523;
  wire n_8525, n_8527, n_8528, n_8529, n_8530, n_8531, n_8532, n_8534;
  wire n_8536, n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544;
  wire n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552;
  wire n_8553, n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560;
  wire n_8561, n_8562, n_8563, n_8564, n_8565, n_8566, n_8567, n_8568;
  wire n_8569, n_8571, n_8573, n_8575, n_8576, n_8577, n_8578, n_8579;
  wire n_8580, n_8582, n_8584, n_8586, n_8587, n_8588, n_8589, n_8590;
  wire n_8591, n_8592, n_8593, n_8594, n_8595, n_8596, n_8597, n_8598;
  wire n_8599, n_8600, n_8601, n_8602, n_8603, n_8604, n_8605, n_8606;
  wire n_8607, n_8608, n_8609, n_8610, n_8611, n_8612, n_8613, n_8615;
  wire n_8617, n_8619, n_8620, n_8621, n_8622, n_8623, n_8624, n_8626;
  wire n_8628, n_8630, n_8631, n_8632, n_8633, n_8634, n_8635, n_8636;
  wire n_8637, n_8638, n_8639, n_8640, n_8641, n_8642, n_8643, n_8644;
  wire n_8645, n_8646, n_8647, n_8648, n_8649, n_8650, n_8651, n_8652;
  wire n_8653, n_8654, n_8655, n_8656, n_8657, n_8658, n_8659, n_8660;
  wire n_8661, n_8662, n_8663, n_8664, n_8665, n_8667, n_8669, n_8671;
  wire n_8672, n_8673, n_8674, n_8675, n_8676, n_8678, n_8680, n_8682;
  wire n_8683, n_8684, n_8685, n_8686, n_8687, n_8688, n_8689, n_8690;
  wire n_8691, n_8692, n_8693, n_8694, n_8695, n_8696, n_8697, n_8698;
  wire n_8699, n_8700, n_8701, n_8702, n_8703, n_8704, n_8705, n_8706;
  wire n_8707, n_8708, n_8709, n_8711, n_8713, n_8715, n_8716, n_8717;
  wire n_8718, n_8719, n_8720, n_8722, n_8724, n_8726, n_8727, n_8728;
  wire n_8729, n_8730, n_8731, n_8732, n_8733, n_8734, n_8735, n_8736;
  wire n_8737, n_8738, n_8739, n_8740, n_8741, n_8742, n_8743, n_8744;
  wire n_8745, n_8746, n_8747, n_8748, n_8749, n_8750, n_8751, n_8752;
  wire n_8753, n_8754, n_8755, n_8756, n_8757, n_8759, n_8761, n_8763;
  wire n_8764, n_8765, n_8766, n_8767, n_8768, n_8770, n_8772, n_8774;
  wire n_8775, n_8776, n_8777, n_8778, n_8779, n_8780, n_8781, n_8782;
  wire n_8783, n_8784, n_8785, n_8786, n_8787, n_8788, n_8789, n_8790;
  wire n_8791, n_8792, n_8793, n_8794, n_8795, n_8796, n_8797, n_8798;
  wire n_8799, n_8800, n_8801, n_8803, n_8805, n_8807, n_8808, n_8809;
  wire n_8810, n_8811, n_8812, n_8814, n_8816, n_8818, n_8819, n_8820;
  wire n_8821, n_8822, n_8823, n_8824, n_8825, n_8826, n_8827, n_8828;
  wire n_8829, n_8830, n_8831, n_8832, n_8833, n_8834, n_8835, n_8836;
  wire n_8837, n_8838, n_8839, n_8840, n_8841, n_8842, n_8843, n_8844;
  wire n_8845, n_8846, n_8847, n_8848, n_8849, n_8850, n_8851, n_8852;
  wire n_8853, n_8854, n_8855, n_8856, n_8857, n_8858, n_8859, n_8860;
  wire n_8861, n_8862, n_8863, n_8864, n_8865, n_8866, n_8867, n_8868;
  wire n_8869, n_8870, n_8871, n_8872, n_8873, n_8874, n_8875, n_8876;
  wire n_8877, n_8878, n_8879, n_8880, n_8881, n_8882, n_8883, n_8884;
  wire n_8885, n_8886, n_8887, n_8888, n_8889, n_8890, n_8891, n_8892;
  wire n_8893, n_8894, n_8895, n_8896, n_8897, n_8898, n_8899, n_8900;
  wire n_8901, n_8902, n_8903, n_8904, n_8905, n_8906, n_8907, n_8908;
  wire n_8909, n_8910, n_8911, n_8912, n_8913, n_8914, n_8915, n_8916;
  wire n_8917, n_8918, n_8919, n_8920, n_8921, n_8922, n_8923, n_8924;
  wire n_8925, n_8926, n_8927, n_8928, n_8929, n_8930, n_8931, n_8932;
  wire n_8933, n_8934, n_8935, n_8936, n_8937, n_8938, n_8939, n_8940;
  wire n_8941, n_8942, n_8943, n_8944, n_8945, n_8946, n_8947, n_8948;
  wire n_8949, n_8950, n_8951, n_8952, n_8953, n_8954, n_8955, n_8956;
  wire n_8957, n_8960, n_8961, n_8962, n_8963, n_8965, n_8966, n_8967;
  wire n_8970, n_8971, n_8972, n_8973, n_8975, n_8976, n_8977, n_8978;
  wire n_8979, n_8980, n_8981, n_8982, n_8983, n_8984, n_8985, n_8986;
  wire n_8987, n_8988, n_8989, n_8990, n_8991, n_8992, n_8993, n_8994;
  wire n_8995, n_8996, n_8997, n_8998, n_8999, n_9000, n_9001, n_9004;
  wire n_9005, n_9006, n_9007, n_9009, n_9010, n_9011, n_9014, n_9015;
  wire n_9016, n_9017, n_9019, n_9020, n_9021, n_9022, n_9023, n_9024;
  wire n_9025, n_9026, n_9027, n_9028, n_9029, n_9030, n_9031, n_9032;
  wire n_9033, n_9034, n_9035, n_9036, n_9037, n_9038, n_9039, n_9040;
  wire n_9041, n_9042, n_9043, n_9044, n_9045, n_9046, n_9047, n_9048;
  wire n_9049, n_9050, n_9051, n_9052, n_9053, n_9054, n_9055, n_9056;
  wire n_9057, n_9058, n_9061, n_9062, n_9063, n_9064, n_9066, n_9067;
  wire n_9068, n_9071, n_9072, n_9073, n_9074, n_9076, n_9077, n_9078;
  wire n_9079, n_9080, n_9081, n_9082, n_9083, n_9084, n_9085, n_9086;
  wire n_9087, n_9088, n_9089, n_9090, n_9091, n_9092, n_9093, n_9094;
  wire n_9095, n_9096, n_9097, n_9098, n_9099, n_9100, n_9101, n_9102;
  wire n_9105, n_9106, n_9107, n_9108, n_9110, n_9111, n_9112, n_9115;
  wire n_9116, n_9117, n_9118, n_9120, n_9121, n_9122, n_9123, n_9124;
  wire n_9125, n_9126, n_9127, n_9128, n_9129, n_9130, n_9131, n_9132;
  wire n_9133, n_9134, n_9135, n_9136, n_9137, n_9138, n_9139, n_9140;
  wire n_9141, n_9142, n_9143, n_9144, n_9145, n_9146, n_9147, n_9148;
  wire n_9149, n_9150, n_9151, n_9152, n_9153, n_9154, n_9155, n_9156;
  wire n_9157, n_9158, n_9159, n_9160, n_9161, n_9162, n_9163, n_9164;
  wire n_9165, n_9166, n_9167, n_9168, n_9169, n_9170, n_9171, n_9172;
  wire n_9173, n_9174, n_9175, n_9176, n_9177, n_9178, n_9179, n_9180;
  wire n_9182, n_9184, n_9186, n_9187, n_9188, n_9189, n_9190, n_9191;
  wire n_9193, n_9195, n_9197, n_9198, n_9199, n_9200, n_9201, n_9202;
  wire n_9203, n_9204, n_9205, n_9206, n_9207, n_9208, n_9209, n_9210;
  wire n_9211, n_9212, n_9213, n_9214, n_9215, n_9216, n_9217, n_9218;
  wire n_9219, n_9220, n_9221, n_9222, n_9223, n_9224, n_9226, n_9228;
  wire n_9230, n_9231, n_9232, n_9233, n_9234, n_9235, n_9237, n_9239;
  wire n_9241, n_9242, n_9243, n_9244, n_9245, n_9246, n_9247, n_9248;
  wire n_9249, n_9250, n_9251, n_9252, n_9253, n_9254, n_9255, n_9256;
  wire n_9257, n_9258, n_9259, n_9260, n_9261, n_9262, n_9263, n_9264;
  wire n_9265, n_9266, n_9267, n_9268, n_9269, n_9270, n_9271, n_9272;
  wire n_9274, n_9276, n_9278, n_9279, n_9280, n_9281, n_9282, n_9283;
  wire n_9285, n_9287, n_9289, n_9290, n_9291, n_9292, n_9293, n_9294;
  wire n_9295, n_9296, n_9297, n_9298, n_9299, n_9300, n_9301, n_9302;
  wire n_9303, n_9304, n_9305, n_9306, n_9307, n_9308, n_9309, n_9310;
  wire n_9311, n_9312, n_9313, n_9314, n_9315, n_9316, n_9318, n_9320;
  wire n_9322, n_9323, n_9324, n_9325, n_9326, n_9327, n_9329, n_9331;
  wire n_9333, n_9334, n_9335, n_9336, n_9337, n_9338, n_9339, n_9340;
  wire n_9341, n_9342, n_9343, n_9344, n_9345, n_9346, n_9347, n_9348;
  wire n_9349, n_9350, n_9351, n_9352, n_9353, n_9354, n_9355, n_9356;
  wire n_9357, n_9358, n_9359, n_9360, n_9361, n_9362, n_9363, n_9364;
  wire n_9365, n_9366, n_9367, n_9368, n_9369, n_9370, n_9371, n_9372;
  wire n_9373, n_9374, n_9375, n_9376, n_9377, n_9378, n_9379, n_9380;
  wire n_9381, n_9382, n_9383, n_9384, n_9385, n_9386, n_9387, n_9388;
  wire n_9389, n_9390, n_9391, n_9392, n_9393, n_9394, n_9395, n_9396;
  wire n_9397, n_9398, n_9399, n_9400, n_9401, n_9402, n_9403, n_9404;
  wire n_9405, n_9406, n_9407, n_9408, n_9409, n_9410, n_9411, n_9412;
  wire n_9413, n_9414, n_9415, n_9416, n_9417, n_9418, n_9419, n_9420;
  wire n_9423, n_9424, n_9425, n_9426, n_9428, n_9429, n_9430, n_9433;
  wire n_9434, n_9435, n_9436, n_9438, n_9439, n_9440, n_9441, n_9442;
  wire n_9443, n_9444, n_9445, n_9446, n_9447, n_9448, n_9449, n_9450;
  wire n_9451, n_9452, n_9453, n_9454, n_9455, n_9456, n_9457, n_9458;
  wire n_9459, n_9460, n_9461, n_9462, n_9463, n_9464, n_9467, n_9468;
  wire n_9469, n_9470, n_9472, n_9473, n_9474, n_9477, n_9478, n_9479;
  wire n_9480, n_9482, n_9483, n_9484, n_9485, n_9486, n_9487, n_9488;
  wire n_9489, n_9490, n_9491, n_9492, n_9493, n_9494, n_9495, n_9496;
  wire n_9497, n_9498, n_9499, n_9500, n_9501, n_9502, n_9503, n_9504;
  wire n_9505, n_9506, n_9507, n_9508, n_9509, n_9510, n_9511, n_9512;
  wire n_9513, n_9514, n_9515, n_9516, n_9517, n_9518, n_9519, n_9520;
  wire n_9521, n_9522, n_9523, n_9525, n_9527, n_9529, n_9530, n_9531;
  wire n_9532, n_9533, n_9534, n_9536, n_9538, n_9540, n_9541, n_9542;
  wire n_9543, n_9544, n_9545, n_9546, n_9547, n_9548, n_9549, n_9550;
  wire n_9551, n_9552, n_9553, n_9554, n_9555, n_9556, n_9557, n_9558;
  wire n_9559, n_9560, n_9561, n_9562, n_9563, n_9564, n_9565, n_9566;
  wire n_9567, n_9569, n_9571, n_9573, n_9574, n_9575, n_9576, n_9577;
  wire n_9578, n_9580, n_9582, n_9584, n_9585, n_9586, n_9587, n_9588;
  wire n_9589, n_9590, n_9591, n_9592, n_9593, n_9594, n_9595, n_9596;
  wire n_9597, n_9598, n_9599, n_9600, n_9601, n_9602, n_9603, n_9604;
  wire n_9605, n_9606, n_9607, n_9608, n_9609, n_9610, n_9611, n_9612;
  wire n_9613, n_9614, n_9615, n_9616, n_9617, n_9618, n_9619, n_9620;
  wire n_9621, n_9622, n_9623, n_9624, n_9625, n_9626, n_9627, n_9628;
  wire n_9629, n_9630, n_9631, n_9632, n_9633, n_9634, n_9635, n_9636;
  wire n_9637, n_9638, n_9639, n_9640, n_9641, n_9642, n_9643, n_9646;
  wire n_9647, n_9648, n_9649, n_9651, n_9652, n_9653, n_9656, n_9657;
  wire n_9658, n_9659, n_9661, n_9662, n_9663, n_9664, n_9665, n_9666;
  wire n_9667, n_9668, n_9669, n_9670, n_9671, n_9672, n_9673, n_9674;
  wire n_9675, n_9676, n_9677, n_9678, n_9679, n_9680, n_9681, n_9682;
  wire n_9683, n_9684, n_9685, n_9686, n_9687, n_9690, n_9691, n_9692;
  wire n_9693, n_9695, n_9696, n_9697, n_9700, n_9701, n_9702, n_9703;
  wire n_9705, n_9706, n_9707, n_9708, n_9709, n_9710, n_9711, n_9712;
  wire n_9713, n_9714, n_9715, n_9716, n_9717, n_9718, n_9719, n_9720;
  wire n_9721, n_9722, n_9723, n_9724, n_9725, n_9726, n_9727, n_9728;
  wire n_9729, n_9730, n_9731, n_9732, n_9733, n_9734, n_9735, n_9736;
  wire n_9737, n_9738, n_9739, n_9740, n_9741, n_9742, n_9743, n_9744;
  wire n_9747, n_9748, n_9749, n_9750, n_9752, n_9753, n_9754, n_9757;
  wire n_9758, n_9759, n_9760, n_9762, n_9763, n_9764, n_9765, n_9766;
  wire n_9767, n_9768, n_9769, n_9770, n_9771, n_9772, n_9773, n_9774;
  wire n_9775, n_9776, n_9777, n_9778, n_9779, n_9780, n_9781, n_9782;
  wire n_9783, n_9784, n_9785, n_9786, n_9787, n_9788, n_9791, n_9792;
  wire n_9793, n_9794, n_9796, n_9797, n_9798, n_9801, n_9802, n_9803;
  wire n_9804, n_9806, n_9807, n_9808, n_9809, n_9810, n_9811, n_9812;
  wire n_9813, n_9814, n_9815, n_9816, n_9817, n_9818, n_9819, n_9820;
  wire n_9821, n_9822, n_9823, n_9824, n_9825, n_9826, n_9827, n_9828;
  wire n_9829, n_9830, n_9831, n_9832, n_9833, n_9834, n_9835, n_9836;
  wire n_9837, n_9838, n_9839, n_9840, n_9841, n_9842, n_9843, n_9844;
  wire n_9845, n_9846, n_9847, n_9848, n_9849, n_9850, n_9851, n_9852;
  wire n_9853, n_9854, n_9855, n_9856, n_9857, n_9858, n_9859, n_9860;
  wire n_9861, n_9862, n_9863, n_9864, n_9865, n_9866, n_9867, n_9868;
  wire n_9869, n_9870, n_9871, n_9872, n_9873, n_9874, n_9875, n_9876;
  wire n_9877, n_9878, n_9879, n_9880, n_9881, n_9882, n_9883, n_9884;
  wire n_9885, n_9886, n_9887, n_9888, n_9889, n_9890, n_9891, n_9892;
  wire n_9893, n_9894, n_9895, n_9896, n_9897, n_9898, n_9899, n_9900;
  wire n_9901, n_9902, n_9903, n_9904, n_9905, n_9906, n_9907, n_9908;
  wire n_9909, n_9910, n_9911, n_9912, n_9913, n_9914, n_9915, n_9916;
  wire n_9917, n_9918, n_9919, n_9920, n_9921, n_9922, n_9923, n_9924;
  wire n_9925, n_9926, n_9927, n_9928, n_9929, n_9930, n_9931, n_9932;
  wire n_9933, n_9934, n_9935, n_9936, n_9937, n_9938, n_9939, n_9940;
  wire n_9941, n_9942, n_9943, n_9944, n_9945, n_9946, n_9947, n_9948;
  wire n_9949, n_9950, n_9951, n_9952, n_9953, n_9954, n_9955, n_9956;
  wire n_9957, n_9958, n_9959, n_9960, n_9961, n_9962, n_9963, n_9964;
  wire n_9965, n_9966, n_9967, n_9968, n_9969, n_9970, n_9971, n_9972;
  wire n_9973, n_9974, n_9975, n_9976, n_9977, n_9978, n_9979, n_9980;
  wire n_9981, n_9982, n_9983, n_9984, n_9985, n_9986, n_9987, n_9988;
  wire n_9989, n_9990, n_9991, n_9992, n_9993, n_9994, n_9995, n_9996;
  wire n_9997, n_9998, n_9999, n_10000, n_10001, n_10002, n_10003,
       n_10004;
  wire n_10005, n_10006, n_10007, n_10008, n_10009, n_10010, n_10011,
       n_10012;
  wire n_10013, n_10014, n_10015, n_10016, n_10017, n_10018, n_10019,
       n_10020;
  wire n_10021, n_10022, n_10023, n_10024, n_10025, n_10026, n_10027,
       n_10028;
  wire n_10029, n_10030, n_10031, n_10032, n_10033, n_10034, n_10035,
       n_10036;
  wire n_10037, n_10038, n_10039, n_10040, n_10041, n_10042, n_10043,
       n_10044;
  wire n_10045, n_10046, n_10047, n_10048, n_10049, n_10050, n_10051,
       n_10052;
  wire n_10053, n_10054, n_10055, n_10056, n_10057, n_10058, n_10059,
       n_10060;
  wire n_10061, n_10062, n_10063, n_10064, n_10065, n_10066, n_10067,
       n_10068;
  wire n_10069, n_10070, n_10071, n_10072, n_10073, n_10074, n_10075,
       n_10076;
  wire n_10077, n_10078, n_10079, n_10080, n_10081, n_10082, n_10083,
       n_10084;
  wire n_10085, n_10086, n_10087, n_10088, n_10089, n_10090, n_10091,
       n_10092;
  wire n_10093, n_10094, n_10095, n_10096, n_10097, n_10098, n_10099,
       n_10100;
  wire n_10101, n_10102, n_10103, n_10104, n_10105, n_10106, n_10107,
       n_10108;
  wire n_10109, n_10110, n_10111, n_10112, n_10113, n_10114, n_10115,
       n_10116;
  wire n_10117, n_10118, n_10119, n_10120, n_10121, n_10122, n_10123,
       n_10124;
  wire n_10125, n_10126, n_10127, n_10128, n_10129, n_10130, n_10131,
       n_10132;
  wire n_10133, n_10134, n_10135, n_10136, n_10137, n_10138, n_10139,
       n_10140;
  wire n_10141, n_10142, n_10143, n_10144, n_10145, n_10146, n_10147,
       n_10148;
  wire n_10149, n_10150, n_10151, n_10152, n_10153, n_10154, n_10155,
       n_10156;
  wire n_10157, n_10158, n_10159, n_10160, n_10161, n_10162, n_10163,
       n_10164;
  wire n_10165, n_10166, n_10167, n_10168, n_10169, n_10170, n_10171,
       n_10172;
  wire n_10173, n_10174, n_10175, n_10176, n_10177, n_10178, n_10179,
       n_10180;
  wire n_10181, n_10182, n_10183, n_10184, n_10185, n_10186, n_10187,
       n_10188;
  wire n_10189, n_10190, n_10191, n_10192, n_10193, n_10194, n_10195,
       n_10196;
  wire n_10197, n_10198, n_10199, n_10200, n_10201, n_10202, n_10203,
       n_10204;
  wire n_10205, n_10206, n_10207, n_10208, n_10209, n_10210, n_10211,
       n_10212;
  wire n_10213, n_10214, n_10215, n_10216, n_10217, n_10218, n_10219,
       n_10220;
  wire n_10221, n_10222, n_10223, n_10224, n_10225, n_10226, n_10227,
       n_10228;
  wire n_10229, n_10230, n_10231, n_10232, n_10233, n_10234, n_10235,
       n_10236;
  wire n_10237, n_10238, n_10239, n_10240, n_10241, n_10242, n_10243,
       n_10244;
  wire n_10245, n_10246, n_10247, n_10248, n_10249, n_10250, n_10251,
       n_10252;
  wire n_10253, n_10254, n_10255, n_10256, n_10257, n_10258, n_10259,
       n_10260;
  wire n_10261, n_10262, n_10263, n_10264, n_10265, n_10266, n_10267,
       n_10268;
  wire n_10269, n_10270, n_10271, n_10272, n_10273, n_10274, n_10275,
       n_10276;
  wire n_10277, n_10278, n_10279, n_10280, n_10281, n_10282, n_10283,
       n_10284;
  wire n_10285, n_10286, n_10287, n_10288, n_10289, n_10290, n_10291,
       n_10292;
  wire n_10293, n_10294, n_10295, n_10296, n_10297, n_10298, n_10299,
       n_10300;
  wire n_10301, n_10302, n_10303, n_10304, n_10305, n_10306, n_10307,
       n_10308;
  wire n_10309, n_10310, n_10311, n_10312, n_10313, n_10314, n_10315,
       n_10316;
  wire n_10317, n_10318, n_10319, n_10320, n_10321, n_10322, n_10323,
       n_10324;
  wire n_10325, n_10326, n_10327, n_10328, n_10329, n_10330, n_10331,
       n_10332;
  wire n_10333, n_10334, n_10335, n_10336, n_10337, n_10338, n_10339,
       n_10340;
  wire n_10341, n_10342, n_10343, n_10344, n_10345, n_10346, n_10347,
       n_10348;
  wire n_10349, n_10350, n_10351, n_10352, n_10353, n_10354, n_10355,
       n_10356;
  wire n_10357, n_10358, n_10359, n_10360, n_10361, n_10362, n_10363,
       n_10364;
  wire n_10365, n_10366, n_10367, n_10368, n_10369, n_10370, n_10371,
       n_10372;
  wire n_10373, n_10374, n_10375, n_10376, n_10377, n_10378, n_10379,
       n_10380;
  wire n_10381, n_10382, n_10383, n_10384, n_10385, n_10386, n_10387,
       n_10388;
  wire n_10389, n_10390, n_10391, n_10392, n_10393, n_10394, n_10395,
       n_10396;
  wire n_10397, n_10398, n_10399, n_10400, n_10401, n_10402, n_10403,
       n_10404;
  wire n_10405, n_10406, n_10407, n_10408, n_10409, n_10410, n_10411,
       n_10412;
  wire n_10413, n_10414, n_10415, n_10416, n_10417, n_10418, n_10419,
       n_10420;
  wire n_10421, n_10422, n_10423, n_10424, n_10425, n_10426, n_10427,
       n_10428;
  wire n_10429, n_10430, n_10431, n_10432, n_10433, n_10434, n_10435,
       n_10436;
  wire n_10437, n_10438, n_10439, n_10440, n_10441, n_10442, n_10443,
       n_10444;
  wire n_10445, n_10446, n_10447, n_10448, n_10449, n_10450, n_10451,
       n_10452;
  wire n_10453, n_10454, n_10455, n_10456, n_10457, n_10458, n_10459,
       n_10460;
  wire n_10461, n_10462, n_10463, n_10464, n_10465, n_10466, n_10467,
       n_10468;
  wire n_10469, n_10470, n_10471, n_10472, n_10473, n_10474, n_10475,
       n_10476;
  wire n_10477, n_10478, n_10479, n_10480, n_10481, n_10482, n_10483,
       n_10484;
  wire n_10485, n_10486, n_10487, n_10488, n_10489, n_10490, n_10491,
       n_10492;
  wire n_10493, n_10494, n_10495, n_10496, n_10497, n_10498, n_10499,
       n_10500;
  wire n_10501, n_10502, n_10503, n_10504, n_10505, n_10506, n_10507,
       n_10508;
  wire n_10509, n_10510, n_10511, n_10512, n_10513, n_10514, n_10515,
       n_10516;
  wire n_10517, n_10518, n_10519, n_10520, n_10521, n_10522, n_10523,
       n_10524;
  wire n_10525, n_10526, n_10527, n_10528, n_10529, n_10530, n_10531,
       n_10532;
  wire n_10533, n_10534, n_10535, n_10536, n_10537, n_10538, n_10539,
       n_10540;
  wire n_10541, n_10542, n_10543, n_10544, n_10545, n_10546, n_10547,
       n_10548;
  wire n_10549, n_10550, n_10551, n_10552, n_10553, n_10554, n_10555,
       n_10556;
  wire n_10557, n_10558, n_10559, n_10560, n_10561, n_10562, n_10563,
       n_10564;
  wire n_10565, n_10566, n_10567, n_10568, n_10569, n_10570, n_10571,
       n_10572;
  wire n_10573, n_10574, n_10575, n_10576, n_10577, n_10578, n_10579,
       n_10580;
  wire n_10581, n_10582, n_10583, n_10584, n_10585, n_10586, n_10587,
       n_10588;
  wire n_10589, n_10590, n_10591, n_10592, n_10593, n_10594, n_10595,
       n_10596;
  wire n_10597, n_10598, n_10599, n_10600, n_10601, n_10602, n_10603,
       n_10604;
  wire n_10605, n_10606, n_10607, n_10608, n_10609, n_10610, n_10611,
       n_10612;
  wire n_10613, n_10614, n_10615, n_10616, n_10617, n_10618, n_10619,
       n_10620;
  wire n_10621, n_10622, n_10623, n_10624, n_10625, n_10626, n_10627,
       n_10628;
  wire n_10629, n_10630, n_10631, n_10632, n_10633, n_10634, n_10635,
       n_10636;
  wire n_10637, n_10638, n_10639, n_10640, n_10641, n_10642, n_10643,
       n_10644;
  wire n_10645, n_10646, n_10647, n_10648, n_10649, n_10650, n_10651,
       n_10652;
  wire n_10653, n_10654, n_10655, n_10656, n_10657, n_10658, n_10659,
       n_10660;
  wire n_10661, n_10662, n_10663, n_10664, n_10665, n_10666, n_10667,
       n_10668;
  wire n_10669, n_10670, n_10671, n_10672, n_10673, n_10674, n_10675,
       n_10676;
  wire n_10677, n_10678, n_10679, n_10680, n_10681, n_10682, n_10683,
       n_10684;
  wire n_10685, n_10686, n_10687, n_10688, n_10689, n_10690, n_10691,
       n_10692;
  wire n_10693, n_10694, n_10695, n_10696, n_10697, n_10698, n_10699,
       n_10700;
  wire n_10701, n_10702, n_10703, n_10704, n_10705, n_10706, n_10707,
       n_10708;
  wire n_10709, n_10710, n_10711, n_10712, n_10713, n_10714, n_10715,
       n_10716;
  wire n_10717, n_10718, n_10719, n_10720, n_10721, n_10722, n_10723,
       n_10724;
  wire n_10725, n_10726, n_10727, n_10728, n_10729, n_10730, n_10731,
       n_10732;
  wire n_10733, n_10734, n_10735, n_10736, n_10737, n_10738, n_10739,
       n_10740;
  wire n_10741, n_10742, n_10743, n_10744, n_10745, n_10746, n_10747,
       n_10748;
  wire n_10749, n_10750, n_10751, n_10752, n_10753, n_10754, n_10755,
       n_10756;
  wire n_10757, n_10758, n_10759, n_10760, n_10761, n_10762, n_10763,
       n_10764;
  wire n_10765, n_10766, n_10767, n_10768, n_10769, n_10770, n_10771,
       n_10772;
  wire n_10773, n_10774, n_10775, n_10776, n_10777, n_10778, n_10779,
       n_10780;
  wire n_10781, n_10782, n_10783, n_10784, n_10785, n_10786, n_10787,
       n_10788;
  wire n_10789, n_10790, n_10791, n_10792, n_10793, n_10794, n_10795,
       n_10796;
  wire n_10797, n_10798, n_10799, n_10800, n_10801, n_10802, n_10803,
       n_10804;
  wire n_10805, n_10806, n_10807, n_10808, n_10809, n_10810, n_10811,
       n_10812;
  wire n_10813, n_10814, n_10815, n_10816, n_10817, n_10818, n_10819,
       n_10820;
  wire n_10821, n_10822, n_10823, n_10824, n_10825, n_10826, n_10827,
       n_10828;
  wire n_10829, n_10830, n_10831, n_10832, n_10833, n_10834, n_10835,
       n_10836;
  wire n_10837, n_10838, n_10839, n_10840, n_10841, n_10842, n_10843,
       n_10844;
  wire n_10845, n_10846, n_10847, n_10848, n_10849, n_10850, n_10851,
       n_10852;
  wire n_10853, n_10854, n_10855, n_10856, n_10857, n_10858, n_10859,
       n_10860;
  wire n_10861, n_10862, n_10863, n_10864, n_10865, n_10866, n_10867,
       n_10868;
  wire n_10869, n_10870, n_10871, n_10872, n_10873, n_10874, n_10875,
       n_10876;
  wire n_10877, n_10878, n_10879, n_10880, n_10881, n_10882, n_10883,
       n_10884;
  wire n_10885, n_10886, n_10887, n_10888, n_10889, n_10890, n_10891,
       n_10892;
  wire n_10893, n_10894, n_10895, n_10896, n_10897, n_10898, n_10899,
       n_10900;
  wire n_10901, n_10902, n_10903, n_10904, n_10905, n_10906, n_10907,
       n_10908;
  wire n_10909, n_10910, n_10911, n_10912, n_10913, n_10914, n_10915,
       n_10916;
  wire n_10917, n_10918, n_10919, n_10920, n_10921, n_10922, n_10923,
       n_10924;
  wire n_10925, n_10926, n_10927, n_10928, n_10929, n_10930, n_10931,
       n_10932;
  wire n_10933, n_10934, n_10935, n_10936, n_10937, n_10938, n_10939,
       n_10940;
  wire n_10941, n_10942, n_10943, n_10944, n_10945, n_10946, n_10947,
       n_10948;
  wire n_10949, n_10950, n_10951, n_10952, n_10953, n_10954, n_10955,
       n_10956;
  wire n_10957, n_10958, n_10959, n_10960, n_10961, n_10962, n_10963,
       n_10964;
  wire n_10965, n_10966, n_10967, n_10968, n_10969, n_10970, n_10971,
       n_10972;
  wire n_10973, n_10974, n_10975, n_10976, n_10977, n_10978, n_10979,
       n_10980;
  wire n_10981, n_10982, n_10983, n_10984, n_10985, n_10986, n_10987,
       n_10988;
  wire n_10989, n_10990, n_10991, n_10992, n_10993, n_10994, n_10995,
       n_10996;
  wire n_10997, n_10998, n_10999, n_11000, n_11001, n_11002, n_11003,
       n_11004;
  wire n_11005, n_11006, n_11007, n_11008, n_11009, n_11010, n_11011,
       n_11012;
  wire n_11013, n_11014, n_11015, n_11016, n_11017, n_11018, n_11019,
       n_11020;
  wire n_11021, n_11022, n_11023, n_11024, n_11025, n_11026, n_11027,
       n_11028;
  wire n_11029, n_11030, n_11031, n_11032, n_11033, n_11034, n_11035,
       n_11036;
  wire n_11037, n_11038, n_11039, n_11040, n_11041, n_11042, n_11043,
       n_11044;
  wire n_11045, n_11046, n_11047, n_11048, n_11049, n_11050, n_11051,
       n_11052;
  wire n_11053, n_11054, n_11055, n_11056, n_11057, n_11058, n_11059,
       n_11060;
  wire n_11061, n_11062, n_11063, n_11064, n_11065, n_11066, n_11067,
       n_11068;
  wire n_11069, n_11070, n_11071, n_11072, n_11073, n_11074, n_11075,
       n_11076;
  wire n_11077, n_11078, n_11079, n_11080, n_11081, n_11082, n_11083,
       n_11084;
  wire n_11085, n_11086, n_11087, n_11088, n_11089, n_11090, n_11091,
       n_11092;
  wire n_11093, n_11094, n_11095, n_11096, n_11097, n_11098, n_11099,
       n_11100;
  wire n_11101, n_11102, n_11103, n_11104, n_11105, n_11106, n_11107,
       n_11108;
  wire n_11109, n_11110, n_11111, n_11112, n_11113, n_11114, n_11115,
       n_11116;
  wire n_11117, n_11118, n_11119, n_11120, n_11121, n_11122, n_11123,
       n_11124;
  wire n_11125, n_11126, n_11127, n_11128, n_11129, n_11130, n_11131,
       n_11132;
  wire n_11133, n_11134, n_11135, n_11136, n_11137, n_11138, n_11139,
       n_11140;
  wire n_11141, n_11142, n_11143, n_11144, n_11145, n_11146, n_11147,
       n_11148;
  wire n_11149, n_11150, n_11151, n_11152, n_11153, n_11154, n_11155,
       n_11156;
  wire n_11157, n_11158, n_11159, n_11160, n_11161, n_11162, n_11163,
       n_11164;
  wire n_11165, n_11166, n_11167, n_11168, n_11169, n_11170, n_11171,
       n_11172;
  wire n_11173, n_11174, n_11175, n_11176, n_11177, n_11178, n_11179,
       n_11180;
  wire n_11181, n_11182, n_11183, n_11184, n_11185, n_11186, n_11187,
       n_11188;
  wire n_11189, n_11190, n_11191, n_11192, n_11193, n_11194, n_11195,
       n_11196;
  wire n_11197, n_11198, n_11199, n_11200, n_11201, n_11202, n_11203,
       n_11204;
  wire n_11205, n_11206, n_11207, n_11208, n_11209, n_11210, n_11211,
       n_11212;
  wire n_11213, n_11214, n_11215, n_11216, n_11217, n_11218, n_11219,
       n_11220;
  wire n_11221, n_11222, n_11223, n_11224, n_11225, n_11226, n_11227,
       n_11228;
  wire n_11229, n_11230, n_11231, n_11232, n_11233, n_11234, n_11235,
       n_11236;
  wire n_11237, n_11238, n_11239, n_11240, n_11241, n_11242, n_11243,
       n_11244;
  wire n_11245, n_11246, n_11247, n_11248, n_11249, n_11250, n_11251,
       n_11252;
  wire n_11253, n_11254, n_11255, n_11256, n_11257, n_11258, n_11259,
       n_11260;
  wire n_11261, n_11262, n_11263, n_11264, n_11265, n_11266, n_11267,
       n_11268;
  wire n_11269, n_11270, n_11271, n_11272, n_11273, n_11274, n_11275,
       n_11276;
  wire n_11277, n_11278, n_11279, n_11280, n_11281, n_11282, n_11283,
       n_11284;
  wire n_11285, n_11286, n_11287, n_11288, n_11289, n_11290, n_11291,
       n_11292;
  wire n_11293, n_11294, n_11295, n_11296, n_11297, n_11298, n_11299,
       n_11300;
  wire n_11301, n_11302, n_11303, n_11304, n_11305, n_11306, n_11307,
       n_11308;
  wire n_11309, n_11310, n_11311, n_11312, n_11313, n_11314, n_11315,
       n_11316;
  wire n_11317, n_11318, n_11319, n_11320, n_11321, n_11322, n_11323,
       n_11324;
  wire n_11325, n_11326, n_11327, n_11328, n_11329, n_11330, n_11331,
       n_11332;
  wire n_11333, n_11334, n_11335, n_11336, n_11337, n_11338, n_11339,
       n_11340;
  wire n_11341, n_11342, n_11343, n_11344, n_11345, n_11346, n_11347,
       n_11348;
  wire n_11349, n_11350, n_11351, n_11352, n_11353, n_11354, n_11355,
       n_11356;
  wire n_11357, n_11358, n_11359, n_11360, n_11361, n_11362, n_11363,
       n_11364;
  wire n_11365, n_11366, n_11367, n_11368, n_11369, n_11370, n_11371,
       n_11372;
  wire n_11373, n_11374, n_11375, n_11376, n_11377, n_11378, n_11379,
       n_11380;
  wire n_11381, n_11382, n_11383, n_11384, n_11385, n_11386, n_11387,
       n_11388;
  wire n_11389, n_11390, n_11391, n_11392, n_11393, n_11394, n_11395,
       n_11396;
  wire n_11397, n_11398, n_11399, n_11400, n_11401, n_11402, n_11403,
       n_11404;
  wire n_11405, n_11406, n_11407, n_11408, n_11409, n_11410, n_11411,
       n_11412;
  wire n_11413, n_11414, n_11415, n_11416, n_11417, n_11418, n_11419,
       n_11420;
  wire n_11421, n_11422, n_11423, n_11424, n_11425, n_11426, n_11427,
       n_11428;
  wire n_11429, n_11430, n_11431, n_11432, n_11433, n_11434, n_11435,
       n_11436;
  wire n_11437, n_11438, n_11439, n_11440, n_11441, n_11442, n_11443,
       n_11444;
  wire n_11445, n_11446, n_11447, n_11448, n_11449, n_11450, n_11451,
       n_11452;
  wire n_11453, n_11454, n_11455, n_11456, n_11457, n_11458, n_11459,
       n_11460;
  wire n_11461, n_11462, n_11463, n_11464, n_11465, n_11466, n_11467,
       n_11468;
  wire n_11469, n_11470, n_11471, n_11472, n_11473, n_11474, n_11475,
       n_11476;
  wire n_11477, n_11478, n_11479, n_11480, n_11481, n_11482, n_11483,
       n_11484;
  wire n_11485, n_11486, n_11487, n_11488, n_11489, n_11490, n_11491,
       n_11492;
  wire n_11493, n_11494, n_11495, n_11496, n_11497, n_11498, n_11499,
       n_11500;
  wire n_11501, n_11502, n_11503, n_11504, n_11505, n_11506, n_11507,
       n_11508;
  wire n_11509, n_11510, n_11511, n_11512, n_11513, n_11514, n_11515,
       n_11516;
  wire n_11517, n_11518, n_11519, n_11520, n_11521, n_11522, n_11523,
       n_11524;
  wire n_11525, n_11526, n_11527, n_11528, n_11529, n_11530, n_11531,
       n_11532;
  wire n_11533, n_11534, n_11535, n_11536, n_11537, n_11538, n_11539,
       n_11540;
  wire n_11541, n_11542, n_11543, n_11544, n_11545, n_11546, n_11547,
       n_11548;
  wire n_11549, n_11550, n_11551, n_11552, n_11553, n_11554, n_11555,
       n_11556;
  wire n_11557, n_11558, n_11559, n_11560, n_11561, n_11562, n_11563,
       n_11564;
  wire n_11565, n_11566, n_11567, n_11568, n_11569, n_11570, n_11571,
       n_11572;
  wire n_11573, n_11574, n_11575, n_11576, n_11577, n_11578, n_11579,
       n_11580;
  wire n_11581, n_11582, n_11583, n_11584, n_11585, n_11586, n_11587,
       n_11588;
  wire n_11589, n_11590, n_11591, n_11592, n_11593, n_11594, n_11595,
       n_11596;
  wire n_11597, n_11598, n_11599, n_11600, n_11601, n_11602, n_11603,
       n_11604;
  wire n_11605, n_11606, n_11607, n_11608, n_11609, n_11610, n_11611,
       n_11612;
  wire n_11613, n_11614, n_11615, n_11616, n_11617, n_11618, n_11619,
       n_11620;
  wire n_11621, n_11622, n_11623, n_11624, n_11625, n_11626, n_11627,
       n_11628;
  wire n_11629, n_11630, n_11631, n_11632, n_11633, n_11634, n_11635,
       n_11636;
  wire n_11637, n_11638, n_11639, n_11640, n_11641, n_11642, n_11643,
       n_11644;
  wire n_11645, n_11646, n_11647, n_11648, n_11649, n_11650, n_11651,
       n_11652;
  wire n_11653, n_11654, n_11655, n_11656, n_11657, n_11658, n_11659,
       n_11660;
  wire n_11661, n_11662, n_11663, n_11664, n_11665, n_11666, n_11667,
       n_11668;
  wire n_11669, n_11670, n_11671, n_11672, n_11673, n_11674, n_11675,
       n_11676;
  wire n_11677, n_11678, n_11679, n_11680, n_11681, n_11682, n_11683,
       n_11684;
  wire n_11685, n_11686, n_11687, n_11688, n_11689, n_11690, n_11691,
       n_11692;
  wire n_11693, n_11694, n_11695, n_11696, n_11697, n_11698, n_11699,
       n_11700;
  wire n_11701, n_11702, n_11703, n_11704, n_11705, n_11706, n_11707,
       n_11708;
  wire n_11709, n_11710, n_11711, n_11712, n_11713, n_11714, n_11715,
       n_11716;
  wire n_11717, n_11718, n_11719, n_11720, n_11721, n_11722, n_11723,
       n_11724;
  wire n_11725, n_11726, n_11727, n_11728, n_11729, n_11730, n_11731,
       n_11732;
  wire n_11733, n_11734, n_11735, n_11736, n_11737, n_11738, n_11739,
       n_11740;
  wire n_11741, n_11742, n_11743, n_11744, n_11745, n_11746, n_11747,
       n_11748;
  wire n_11749, n_11750, n_11751, n_11752, n_11753, n_11754, n_11755,
       n_11756;
  wire n_11757, n_11758, n_11759, n_11760, n_11761, n_11762, n_11763,
       n_11764;
  wire n_11765, n_11766, n_11767, n_11768, n_11769, n_11770, n_11771,
       n_11772;
  wire n_11773, n_11774, n_11775, n_11776, n_11777, n_11778, n_11779,
       n_11780;
  wire n_11781, n_11782, n_11783, n_11784, n_11785, n_11786, n_11787,
       n_11788;
  wire n_11789, n_11790, n_11791, n_11792, n_11793, n_11794, n_11795,
       n_11796;
  wire n_11797, n_11798, n_11799, n_11800, n_11801, n_11802, n_11803,
       n_11804;
  wire n_11805, n_11806, n_11807, n_11808, n_11809, n_11810, n_11811,
       n_11812;
  wire n_11813, n_11814, n_11815, n_11816, n_11817, n_11818, n_11819,
       n_11820;
  wire n_11821, n_11822, n_11823, n_11824, n_11825, n_11826, n_11827,
       n_11828;
  wire n_11829, n_11830, n_11831, n_11832, n_11833, n_11834, n_11835,
       n_11836;
  wire n_11837, n_11838, n_11839, n_11840, n_11841, n_11842, n_11843,
       n_11844;
  wire n_11845, n_11846, n_11847, n_11848, n_11849, n_11850, n_11851,
       n_11852;
  wire n_11853, n_11854, n_11855, n_11856, n_11857, n_11858, n_11859,
       n_11860;
  wire n_11861, n_11862, n_11863, n_11864, n_11865, n_11866, n_11867,
       n_11868;
  wire n_11869, n_11870, n_11871, n_11872, n_11873, n_11874, n_11875,
       n_11876;
  wire n_11877, n_11878, n_11879, n_11880, n_11881, n_11882, n_11883,
       n_11884;
  wire n_11885, n_11886, n_11887, n_11888, n_11889, n_11890, n_11891,
       n_11892;
  wire n_11893, n_11894, n_11895, n_11896, n_11897, n_11898, n_11899,
       n_11900;
  wire n_11901, n_11902, n_11903, n_11904, n_11905, n_11906, n_11907,
       n_11908;
  wire n_11909, n_11910, n_11911, n_11912, n_11913, n_11914, n_11915,
       n_11916;
  wire n_11917, n_11918, n_11919, n_11920, n_11921, n_11922, n_11923,
       n_11924;
  wire n_11925, n_11926, n_11927, n_11928, n_11929, n_11930, n_11931,
       n_11932;
  wire n_11933, n_11934, n_11935, n_11936, n_11937, n_11938, n_11939,
       n_11940;
  wire n_11941, n_11942, n_11943, n_11944, n_11945, n_11946, n_11947,
       n_11948;
  wire n_11949, n_11950, n_11951, n_11952, n_11953, n_11954, n_11955,
       n_11956;
  wire n_11957, n_11958, n_11959, n_11960, n_11961, n_11962, n_11963,
       n_11964;
  wire n_11965, n_11966, n_11967, n_11968, n_11969, n_11970, n_11971,
       n_11972;
  wire n_11973, n_11974, n_11975, n_11976, n_11977, n_11978, n_11979,
       n_11980;
  wire n_11981, n_11982, n_11983, n_11984, n_11985, n_11986, n_11987,
       n_11988;
  wire n_11989, n_11990, n_11991, n_11992, n_11993, n_11994, n_11995,
       n_11996;
  wire n_11997, n_11998, n_11999, n_12000, n_12001, n_12002, n_12003,
       n_12004;
  wire n_12005, n_12006, n_12007, n_12008, n_12009, n_12010, n_12011,
       n_12012;
  wire n_12013, n_12014, n_12015, n_12016, n_12017, n_12018, n_12019,
       n_12020;
  wire n_12021, n_12022, n_12023, n_12024, n_12025, n_12026, n_12027,
       n_12028;
  wire n_12029, n_12030, n_12031, n_12032, n_12033, n_12034, n_12035,
       n_12036;
  wire n_12037, n_12038, n_12039, n_12040, n_12041, n_12042, n_12043,
       n_12044;
  wire n_12045, n_12046, n_12047, n_12048, n_12049, n_12050, n_12051,
       n_12052;
  wire n_12053, n_12054, n_12055, n_12056, n_12057, n_12058, n_12059,
       n_12060;
  wire n_12061, n_12062, n_12063, n_12064, n_12065, n_12066, n_12067,
       n_12068;
  wire n_12069, n_12070, n_12071, n_12072, n_12073, n_12074, n_12075,
       n_12076;
  wire n_12077, n_12078, n_12079, n_12080, n_12081, n_12082, n_12083,
       n_12084;
  wire n_12085, n_12086, n_12087, n_12088, n_12089, n_12090, n_12091,
       n_12092;
  wire n_12093, n_12094, n_12095, n_12096, n_12097, n_12098, n_12099,
       n_12100;
  wire n_12101, n_12102, n_12103, n_12104, n_12105, n_12106, n_12107,
       n_12108;
  wire n_12109, n_12110, n_12111, n_12112, n_12113, n_12114, n_12115,
       n_12116;
  wire n_12117, n_12118, n_12119, n_12120, n_12121, n_12122, n_12123,
       n_12124;
  wire n_12125, n_12126, n_12127, n_12128, n_12129, n_12130, n_12131,
       n_12132;
  wire n_12133, n_12134, n_12135, n_12136, n_12137, n_12138, n_12139,
       n_12140;
  wire n_12141, n_12142, n_12143, n_12144, n_12145, n_12146, n_12147,
       n_12148;
  wire n_12149, n_12150, n_12151, n_12152, n_12153, n_12154, n_12155,
       n_12156;
  wire n_12157, n_12158, n_12159, n_12160, n_12161, n_12162, n_12163,
       n_12164;
  wire n_12165, n_12166, n_12167, n_12168, n_12169, n_12170, n_12171,
       n_12172;
  wire n_12173, n_12174, n_12175, n_12176, n_12177, n_12178, n_12179,
       n_12180;
  wire n_12181, n_12182, n_12183, n_12184, n_12185, n_12186, n_12187,
       n_12188;
  wire n_12189, n_12190, n_12191, n_12192, n_12193, n_12194, n_12195,
       n_12196;
  wire n_12197, n_12198, n_12199, n_12200, n_12201, n_12202, n_12203,
       n_12204;
  wire n_12205, n_12206, n_12207, n_12208, n_12209, n_12210, n_12211,
       n_12212;
  wire n_12213, n_12214, n_12215, n_12216, n_12217, n_12218, n_12219,
       n_12220;
  wire n_12221, n_12222, n_12223, n_12224, n_12225, n_12226, n_12227,
       n_12228;
  wire n_12229, n_12230, n_12231, n_12232, n_12233, n_12234, n_12235,
       n_12236;
  wire n_12237, n_12238, n_12239, n_12240, n_12241, n_12242, n_12243,
       n_12244;
  wire n_12245, n_12246, n_12247, n_12248, n_12249, n_12250, n_12251,
       n_12252;
  wire n_12253, n_12254, n_12255, n_12256, n_12257, n_12258, n_12259,
       n_12260;
  wire n_12261, n_12262, n_12263, n_12264, n_12265, n_12266, n_12267,
       n_12268;
  wire n_12269, n_12270, n_12271, n_12272, n_12273, n_12274, n_12275,
       n_12276;
  wire n_12277, n_12278, n_12279, n_12280, n_12281, n_12282, n_12283,
       n_12284;
  wire n_12285, n_12286, n_12287, n_12288, n_12289, n_12290, n_12291,
       n_12292;
  wire n_12293, n_12294, n_12295, n_12296, n_12297, n_12298, n_12299,
       n_12300;
  wire n_12301, n_12302, n_12303, n_12304, n_12305, n_12306, n_12307,
       n_12308;
  wire n_12309, n_12310, n_12311, n_12312, n_12313, n_12314, n_12315,
       n_12316;
  wire n_12317, n_12318, n_12319, n_12320, n_12321, n_12322, n_12323,
       n_12324;
  wire n_12325, n_12326, n_12327, n_12328, n_12329, n_12330, n_12331,
       n_12332;
  wire n_12333, n_12334, n_12335, n_12336, n_12337, n_12338, n_12339,
       n_12340;
  wire n_12341, n_12342, n_12343, n_12344, n_12345, n_12346, n_12347,
       n_12348;
  wire n_12349, n_12350, n_12351, n_12352, n_12353, n_12354, n_12355,
       n_12356;
  wire n_12357, n_12358, n_12359, n_12360, n_12361, n_12362, n_12363,
       n_12364;
  wire n_12365, n_12366, n_12367, n_12368, n_12369, n_12370, n_12371,
       n_12372;
  wire n_12373, n_12374, n_12375, n_12376, n_12377, n_12378, n_12379,
       n_12380;
  wire n_12381, n_12382, n_12383, n_12384, n_12385, n_12386, n_12387,
       n_12388;
  wire n_12389, n_12390, n_12391, n_12392, n_12393, n_12394, n_12395,
       n_12396;
  wire n_12397, n_12398, n_12399, n_12400, n_12401, n_12402, n_12403,
       n_12404;
  wire n_12405, n_12406, n_12407, n_12408, n_12409, n_12410, n_12411,
       n_12412;
  wire n_12413, n_12414, n_12415, n_12416, n_12417, n_12418, n_12419,
       n_12420;
  wire n_12421, n_12422, n_12423, n_12424, n_12425, n_12426, n_12427,
       n_12428;
  wire n_12429, n_12430, n_12431, n_12432, n_12433, n_12434, n_12435,
       n_12436;
  wire n_12437, n_12438, n_12439, n_12440, n_12441, n_12442, n_12443,
       n_12444;
  wire n_12445, n_12446, n_12447, n_12448, n_12449, n_12450, n_12451,
       n_12452;
  wire n_12453, n_12454, n_12455, n_12456, n_12457, n_12458, n_12459,
       n_12460;
  wire n_12461, n_12462, n_12463, n_12464, n_12465, n_12466, n_12467,
       n_12468;
  wire n_12469, n_12470, n_12471, n_12472, n_12473, n_12474, n_12475,
       n_12476;
  wire n_12477, n_12478, n_12479, n_12480, n_12481, n_12482, n_12483,
       n_12484;
  wire n_12485, n_12486, n_12487, n_12488, n_12489, n_12490, n_12491,
       n_12492;
  wire n_12493, n_12494, n_12495, n_12496, n_12497, n_12498, n_12499,
       n_12500;
  wire n_12501, n_12502, n_12503, n_12504, n_12505, n_12506, n_12507,
       n_12508;
  wire n_12509, n_12510, n_12511, n_12512, n_12513, n_12514, n_12515,
       n_12516;
  wire n_12517, n_12518, n_12519, n_12520, n_12521, n_12522, n_12523,
       n_12524;
  wire n_12525, n_12526, n_12527, n_12528, n_12529, n_12530, n_12531,
       n_12532;
  wire n_12533, n_12534, n_12535, n_12536, n_12537, n_12538, n_12539,
       n_12540;
  wire n_12541, n_12542, n_12543, n_12544, n_12545, n_12546, n_12547,
       n_12548;
  wire n_12549, n_12550, n_12551, n_12552, n_12553, n_12554, n_12555,
       n_12556;
  wire n_12557, n_12558, n_12559, n_12560, n_12561, n_12562, n_12563,
       n_12564;
  wire n_12565, n_12566, n_12567, n_12568, n_12569, n_12570, n_12571,
       n_12572;
  wire n_12573, n_12574, n_12575, n_12576, n_12577, n_12578, n_12579,
       n_12580;
  wire n_12581, n_12582, n_12583, n_12584, n_12585, n_12586, n_12587,
       n_12588;
  wire n_12589, n_12590, n_12591, n_12592, n_12593, n_12594, n_12595,
       n_12596;
  wire n_12597, n_12598, n_12599, n_12600, n_12601, n_12602, n_12603,
       n_12604;
  wire n_12605, n_12606, n_12607, n_12608, n_12609, n_12610, n_12611,
       n_12612;
  wire n_12613, n_12614, n_12615, n_12616, n_12617, n_12618, n_12619,
       n_12620;
  wire n_12621, n_12622, n_12623, n_12624, n_12625, n_12626, n_12627,
       n_12628;
  wire n_12629, n_12630, n_12631, n_12632, n_12633, n_12634, n_12635,
       n_12636;
  wire n_12637, n_12638, n_12639, n_12640, n_12641, n_12642, n_12643,
       n_12644;
  wire n_12645, n_12646, n_12647, n_12648, n_12649, n_12650, n_12651,
       n_12652;
  wire n_12653, n_12654, n_12655, n_12656, n_12657, n_12658, n_12659,
       n_12660;
  wire n_12661, n_12662, n_12663, n_12664, n_12665, n_12666, n_12667,
       n_12668;
  wire n_12669, n_12670, n_12671, n_12672, n_12673, n_12674, n_12675,
       n_12676;
  wire n_12677, n_12678, n_12679, n_12680, n_12681, n_12682, n_12683,
       n_12684;
  wire n_12685, n_12686, n_12687, n_12688, n_12689, n_12690, n_12691,
       n_12692;
  wire n_12693, n_12694, n_12695, n_12696, n_12697, n_12698, n_12699,
       n_12700;
  wire n_12701, n_12702, n_12703, n_12704, n_12705, n_12706, n_12707,
       n_12708;
  wire n_12709, n_12710, n_12711, n_12712, n_12713, n_12714, n_12715,
       n_12716;
  wire n_12717, n_12718, n_12719, n_12720, n_12721, n_12722, n_12723,
       n_12724;
  wire n_12725, n_12726, n_12727, n_12728, n_12729, n_12730, n_12731,
       n_12732;
  wire n_12733, n_12734, n_12735, n_12736, n_12737, n_12738, n_12739,
       n_12740;
  wire n_12741, n_12742, n_12743, n_12744, n_12745, n_12746, n_12747,
       n_12748;
  wire n_12749, n_12750, n_12751, n_12752, n_12753, n_12754, n_12755,
       n_12756;
  wire n_12757, n_12758, n_12759, n_12760, n_12761, n_12762, n_12763,
       n_12764;
  wire n_12765, n_12766, n_12767, n_12768, n_12769, n_12770, n_12771,
       n_12772;
  wire n_12773, n_12774, n_12775, n_12776, n_12777, n_12778, n_12779,
       n_12780;
  wire n_12781, n_12782, n_12783, n_12784, n_12785, n_12786, n_12787,
       n_12788;
  wire n_12789, n_12790, n_12791, n_12792, n_12793, n_12794, n_12795,
       n_12796;
  wire n_12797, n_12798, n_12799, n_12800, n_12801, n_12802, n_12803,
       n_12804;
  wire n_12805, n_12806, n_12807, n_12808, n_12809, n_12810, n_12811,
       n_12812;
  wire n_12813, n_12814, n_12815, n_12816, n_12817, n_12818, n_12819,
       n_12820;
  wire n_12821, n_12822, n_12823, n_12824, n_12825, n_12826, n_12827,
       n_12828;
  wire n_12829, n_12830, n_12831, n_12832, n_12833, n_12834, n_12835,
       n_12836;
  wire n_12837, n_12838, n_12839, n_12840, n_12841, n_12842, n_12843,
       n_12844;
  wire n_12845, n_12846, n_12847, n_12848, n_12849, n_12850, n_12851,
       n_12852;
  wire n_12853, n_12854, n_12855, n_12856, n_12857, n_12858, n_12859,
       n_12860;
  wire n_12861, n_12862, n_12863, n_12864, n_12865, n_12866, n_12867,
       n_12868;
  wire n_12869, n_12870, n_12871, n_12872, n_12873, n_12874, n_12875,
       n_12876;
  wire n_12877, n_12878, n_12879, n_12880, n_12881, n_12882, n_12883,
       n_12884;
  wire n_12885, n_12886, n_12887, n_12888, n_12889, n_12890, n_12891,
       n_12892;
  wire n_12893, n_12894, n_12895, n_12896, n_12897, n_12898, n_12899,
       n_12900;
  wire n_12901, n_12902, n_12903, n_12904, n_12905, n_12906, n_12907,
       n_12908;
  wire n_12909, n_12910, n_12911, n_12912, n_12913, n_12914, n_12915,
       n_12916;
  wire n_12917, n_12918, n_12919, n_12920, n_12921, n_12922, n_12923,
       n_12924;
  wire n_12925, n_12926, n_12927, n_12928, n_12929, n_12930, n_12931,
       n_12932;
  wire n_12933, n_12934, n_12935, n_12936, n_12937, n_12938, n_12939,
       n_12940;
  wire n_12941, n_12942, n_12943, n_12944, n_12945, n_12946, n_12947,
       n_12948;
  wire n_12949, n_12950, n_12951, n_12952, n_12953, n_12954, n_12955,
       n_12956;
  wire n_12957, n_12958, n_12959, n_12960, n_12961, n_12962, n_12963,
       n_12964;
  wire n_12965, n_12966, n_12967, n_12968, n_12969, n_12970, n_12971,
       n_12972;
  wire n_12973, n_12974, n_12975, n_12976, n_12977, n_12978, n_12979,
       n_12980;
  wire n_12981, n_12982, n_12983, n_12984, n_12985, n_12986, n_12987,
       n_12988;
  wire n_12989, n_12990, n_12991, n_12992, n_12993, n_12994, n_12995,
       n_12996;
  wire n_12997, n_12998, n_12999, n_13000, n_13001, n_13002, n_13003,
       n_13004;
  wire n_13005, n_13006, n_13007, n_13008, n_13009, n_13010, n_13011,
       n_13012;
  wire n_13013, n_13014, n_13015, n_13016, n_13017, n_13018, n_13019,
       n_13020;
  wire n_13021, n_13022, n_13023, n_13024, n_13025, n_13026, n_13027,
       n_13028;
  wire n_13029, n_13030, n_13031, n_13032, n_13033, n_13034, n_13035,
       n_13036;
  wire n_13037, n_13038, n_13039, n_13040, n_13041, n_13042, n_13043,
       n_13044;
  wire n_13045, n_13046, n_13047, n_13048, n_13049, n_13050, n_13051,
       n_13052;
  wire n_13053, n_13054, n_13055, n_13056, n_13057, n_13058, n_13059,
       n_13060;
  wire n_13061, n_13062, n_13063, n_13064, n_13065, n_13066, n_13067,
       n_13068;
  wire n_13069, n_13070, n_13071, n_13072, n_13073, n_13074, n_13075,
       n_13076;
  wire n_13077, n_13078, n_13079, n_13080, n_13081, n_13082, n_13083,
       n_13084;
  wire n_13085, n_13086, n_13087, n_13088, n_13089, n_13090, n_13091,
       n_13092;
  wire n_13093, n_13094, n_13095, n_13096, n_13097, n_13098, n_13099,
       n_13100;
  wire n_13101, n_13102, n_13103, n_13104, n_13105, n_13106, n_13107,
       n_13108;
  wire n_13109, n_13110, n_13111, n_13112, n_13113, n_13114, n_13115,
       n_13116;
  wire n_13117, n_13118, n_13119, n_13120, n_13121, n_13122, n_13123,
       n_13124;
  wire n_13125, n_13126, n_13127, n_13128, n_13129, n_13130, n_13131,
       n_13132;
  wire n_13133, n_13134, n_13135, n_13136, n_13137, n_13138, n_13139,
       n_13140;
  wire n_13141, n_13142, n_13143, n_13144, n_13145, n_13146, n_13147,
       n_13148;
  wire n_13149, n_13150, n_13151, n_13152, n_13153, n_13154, n_13155,
       n_13156;
  wire n_13157, n_13158, n_13159, n_13160, n_13161, n_13162, n_13163,
       n_13164;
  wire n_13165, n_13166, n_13167, n_13168, n_13169, n_13170, n_13171,
       n_13172;
  wire n_13173, n_13174, n_13175, n_13176, n_13177, n_13178, n_13179,
       n_13180;
  wire n_13181, n_13182, n_13183, n_13184, n_13185, n_13186, n_13187,
       n_13188;
  wire n_13189, n_13190, n_13191, n_13192, n_13193, n_13194, n_13195,
       n_13196;
  wire n_13197, n_13198, n_13199, n_13200, n_13201, n_13202, n_13203,
       n_13204;
  wire n_13205, n_13206, n_13207, n_13208, n_13209, n_13210, n_13211,
       n_13212;
  wire n_13213, n_13214, n_13215, n_13216, n_13217, n_13218, n_13219,
       n_13220;
  wire n_13221, n_13222, n_13223, n_13224, n_13225, n_13226, n_13227,
       n_13228;
  wire n_13229, n_13230, n_13231, n_13232, n_13233, n_13234, n_13235,
       n_13236;
  wire n_13237, n_13238, n_13239, n_13240, n_13241, n_13242, n_13243,
       n_13244;
  wire n_13245, n_13246, n_13247, n_13248, n_13249, n_13250, n_13251,
       n_13252;
  wire n_13253, n_13254, n_13255, n_13256, n_13257, n_13258, n_13259,
       n_13260;
  wire n_13261, n_13262, n_13263, n_13264, n_13265, n_13266, n_13267,
       n_13268;
  wire n_13269, n_13270, n_13271, n_13272, n_13273, n_13274, n_13275,
       n_13276;
  wire n_13277, n_13278, n_13279, n_13280, n_13281, n_13282, n_13283,
       n_13284;
  wire n_13285, n_13286, n_13287, n_13288, n_13289, n_13290, n_13291,
       n_13292;
  wire n_13293, n_13294, n_13295, n_13296, n_13297, n_13298, n_13299,
       n_13300;
  wire n_13301, n_13302, n_13303, n_13304, n_13305, n_13306, n_13307,
       n_13308;
  wire n_13309, n_13310, n_13311, n_13312, n_13313, n_13314, n_13315,
       n_13316;
  wire n_13317, n_13318, n_13319, n_13320, n_13321, n_13322, n_13323,
       n_13324;
  wire n_13325, n_13326, n_13327, n_13328, n_13329, n_13330, n_13331,
       n_13332;
  wire n_13333, n_13334, n_13335, n_13336, n_13337, n_13338, n_13339,
       n_13340;
  wire n_13341, n_13342, n_13343, n_13344, n_13345, n_13346, n_13347,
       n_13348;
  wire n_13349, n_13350, n_13351, n_13352, n_13353, n_13354, n_13355,
       n_13356;
  wire n_13357, n_13358, n_13359, n_13360, n_13361, n_13362, n_13363,
       n_13364;
  wire n_13365, n_13366, n_13367, n_13368, n_13369, n_13370, n_13371,
       n_13372;
  wire n_13373, n_13374, n_13375, n_13376, n_13377, n_13378, n_13379,
       n_13380;
  wire n_13381, n_13382, n_13383, n_13384, n_13385, n_13386, n_13387,
       n_13388;
  wire n_13389, n_13390, n_13391, n_13392, n_13393, n_13394, n_13395,
       n_13396;
  wire n_13397, n_13398, n_13399, n_13400, n_13401, n_13402, n_13403,
       n_13404;
  wire n_13405, n_13406, n_13407, n_13408, n_13409, n_13410, n_13411,
       n_13412;
  wire n_13413, n_13414, n_13415, n_13416, n_13417, n_13418, n_13419,
       n_13420;
  wire n_13421, n_13422, n_13423, n_13424, n_13425, n_13426, n_13427,
       n_13428;
  wire n_13429, n_13430, n_13431, n_13432, n_13433, n_13434, n_13435,
       n_13436;
  wire n_13437, n_13438, n_13439, n_13440, n_13441, n_13442, n_13443,
       n_13444;
  wire n_13445, n_13446, n_13447, n_13448, n_13449, n_13450, n_13451,
       n_13452;
  wire n_13453, n_13454, n_13455, n_13456, n_13457, n_13458, n_13459,
       n_13460;
  wire n_13461, n_13462, n_13463, n_13464, n_13465, n_13466, n_13467,
       n_13468;
  wire n_13469, n_13470, n_13471, n_13472, n_13473, n_13474, n_13475,
       n_13476;
  wire n_13477, n_13478, n_13479, n_13480, n_13481, n_13482, n_13483,
       n_13484;
  wire n_13485, n_13486, n_13487, n_13488, n_13489, n_13490, n_13491,
       n_13492;
  wire n_13493, n_13494, n_13495, n_13496, n_13497, n_13498, n_13499,
       n_13500;
  wire n_13501, n_13502, n_13503, n_13504, n_13505, n_13506, n_13507,
       n_13508;
  wire n_13509, n_13510, n_13511, n_13512, n_13513, n_13514, n_13515,
       n_13516;
  wire n_13517, n_13518, n_13519, n_13520, n_13521, n_13522, n_13523,
       n_13524;
  wire n_13525, n_13526, n_13527, n_13528, n_13529, n_13530, n_13531,
       n_13532;
  wire n_13533, n_13534, n_13535, n_13536, n_13537, n_13538, n_13539,
       n_13540;
  wire n_13541, n_13542, n_13543, n_13544, n_13545, n_13546, n_13547,
       n_13548;
  wire n_13549, n_13550, n_13551, n_13552, n_13553, n_13554, n_13555,
       n_13556;
  wire n_13557, n_13558, n_13559, n_13560, n_13561, n_13562, n_13563,
       n_13564;
  wire n_13565, n_13566, n_13567, n_13568, n_13569, n_13570, n_13571,
       n_13572;
  wire n_13573, n_13574, n_13575, n_13576, n_13577, n_13578, n_13579,
       n_13580;
  wire n_13581, n_13582, n_13583, n_13584, n_13585, n_13586, n_13587,
       n_13588;
  wire n_13589, n_13590, n_13591, n_13592, n_13593, n_13594, n_13595,
       n_13596;
  wire n_13597, n_13598, n_13599, n_13600, n_13601, n_13602, n_13603,
       n_13604;
  wire n_13605, n_13606, n_13607, n_13608, n_13609, n_13610, n_13611,
       n_13612;
  wire n_13613, n_13614, n_13615, n_13616, n_13617, n_13618, n_13619,
       n_13620;
  wire n_13621, n_13622, n_13623, n_13624, n_13625, n_13626, n_13627,
       n_13628;
  wire n_13629, n_13630, n_13631, n_13632, n_13633, n_13634, n_13635,
       n_13636;
  wire n_13637, n_13638, n_13639, n_13640, n_13641, n_13642, n_13643,
       n_13644;
  wire n_13645, n_13646, n_13647, n_13648, n_13649, n_13650, n_13651,
       n_13652;
  wire n_13653, n_13654, n_13655, n_13656, n_13657, n_13658, n_13659,
       n_13660;
  wire n_13661, n_13662, n_13663, n_13664, n_13665, n_13666, n_13667,
       n_13668;
  wire n_13669, n_13670, n_13671, n_13672, n_13673, n_13674, n_13675,
       n_13676;
  wire n_13677, n_13678, n_13679, n_13680, n_13681, n_13682, n_13683,
       n_13684;
  wire n_13685, n_13686, n_13687, n_13688, n_13689, n_13690, n_13691,
       n_13692;
  wire n_13693, n_13694, n_13695, n_13696, n_13697, n_13698, n_13699,
       n_13700;
  wire n_13701, n_13702, n_13703, n_13704, n_13705, n_13706, n_13707,
       n_13708;
  wire n_13709, n_13710, n_13711, n_13712, n_13713, n_13714, n_13715,
       n_13716;
  wire n_13717, n_13718, n_13719, n_13720, n_13721, n_13722, n_13723,
       n_13724;
  wire n_13725, n_13726, n_13727, n_13728, n_13729, n_13730, n_13731,
       n_13732;
  wire n_13733, n_13734, n_13735, n_13736, n_13737, n_13738, n_13739,
       n_13740;
  wire n_13741, n_13742, n_13743, n_13744, n_13745, n_13746, n_13747,
       n_13748;
  wire n_13749, n_13750, n_13751, n_13752, n_13753, n_13754, n_13755,
       n_13756;
  wire n_13757, n_13758, n_13759, n_13760, n_13761, n_13762, n_13763,
       n_13764;
  wire n_13765, n_13766, n_13767, n_13768, n_13769, n_13770, n_13771,
       n_13772;
  wire n_13773, n_13774, n_13775, n_13776, n_13777, n_13778, n_13779,
       n_13780;
  wire n_13781, n_13782, n_13783, n_13784, n_13785, n_13786, n_13787,
       n_13788;
  wire n_13789, n_13790, n_13791, n_13792, n_13793, n_13794, n_13795,
       n_13796;
  wire n_13797, n_13798, n_13799, n_13800, n_13801, n_13802, n_13803,
       n_13804;
  wire n_13805, n_13806, n_13807, n_13808, n_13809, n_13810, n_13811,
       n_13812;
  wire n_13813, n_13814, n_13815, n_13816, n_13817, n_13818, n_13819,
       n_13820;
  wire n_13821, n_13822, n_13823, n_13824, n_13825, n_13826, n_13827,
       n_13828;
  wire n_13829, n_13830, n_13831, n_13832, n_13833, n_13834, n_13835,
       n_13836;
  wire n_13837, n_13838, n_13839, n_13840, n_13841, n_13842, n_13843,
       n_13845;
  wire n_13846, n_13847, n_13848, n_13849, n_13850, n_13851, n_13852,
       n_13853;
  wire n_13854, n_13855, n_13856, n_13857, n_13858, n_13859, n_13860,
       n_13861;
  wire n_13862, n_13863, n_13864, n_13865, n_13866, n_13867, n_13868,
       n_13869;
  wire n_13870, n_13871, n_13872, n_13873, n_13874, n_13875, n_13876,
       n_13877;
  wire n_13878, n_13879, n_13880, n_13881, n_13882, n_13883, n_13884,
       n_13885;
  wire n_13886, n_13887, n_13888, n_13889, n_13890, n_13891, n_13892,
       n_13893;
  wire n_13894, n_13895, n_13896, n_13897, n_13898, n_13899, n_13900,
       n_13901;
  wire n_13902, n_13903, n_13905, n_13906, n_13907, n_13908, n_13909,
       n_13910;
  wire n_13911, n_13912, n_13913, n_13914, n_13915, n_13916, n_13917,
       n_13918;
  wire n_13919, n_13920, n_13921, n_13922, n_13923, n_13924, n_13925,
       n_13926;
  wire n_13927, n_13928, n_13929, n_13930, n_13931, n_13932, n_13933,
       n_13934;
  wire n_13935, n_13936, n_13937, n_13938, n_13939, n_13940, n_13941,
       n_13942;
  wire n_13943, n_13944, n_13945, n_13946, n_13947, n_13948, n_13949,
       n_13950;
  wire n_13951, n_13952, n_13953, n_13954, n_13955, n_13956, n_13957,
       n_13958;
  wire n_13959, n_13960, n_13961, n_13963, n_13964, n_13966, n_13967,
       n_13968;
  wire n_13969, n_13970, n_13971, n_13972, n_13973, n_13974, n_13975,
       n_13976;
  wire n_13977, n_13978, n_13979, n_13980, n_13981, n_13982, n_13983,
       n_13984;
  wire n_13985, n_13986, n_13987, n_13988, n_13989, n_13990, n_13991,
       n_13992;
  wire n_13993, n_13994, n_13995, n_13996, n_13997, n_13998, n_13999,
       n_14000;
  wire n_14001, n_14002, n_14003, n_14004, n_14005, n_14006, n_14007,
       n_14008;
  wire n_14009, n_14010, n_14011, n_14012, n_14013, n_14014, n_14015,
       n_14016;
  wire n_14017, n_14018, n_14019, n_14020, n_14021, n_14022, n_14023,
       n_14024;
  wire n_14025, n_14026, n_14027, n_14028, n_14029, n_14030, n_14031,
       n_14032;
  wire n_14033, n_14034, n_14035, n_14036, n_14037, n_14038, n_14039,
       n_14040;
  wire n_14041, n_14042, n_14043, n_14044, n_14045, n_14046, n_14047,
       n_14048;
  and g1 (n1003, \A[718] , \A[719] );
  not g2 (n_3, \A[719] );
  and g3 (n1004, \A[718] , n_3);
  not g4 (n_4, \A[718] );
  and g5 (n1005, n_4, \A[719] );
  not g6 (n_5, n1004);
  not g7 (n_6, n1005);
  and g8 (n1006, n_5, n_6);
  not g9 (n_8, n1006);
  and g10 (n1007, \A[720] , n_8);
  not g11 (n_9, n1003);
  not g12 (n_10, n1007);
  and g13 (n1008, n_9, n_10);
  and g14 (n1009, \A[715] , \A[716] );
  not g15 (n_13, \A[716] );
  and g16 (n1010, \A[715] , n_13);
  not g17 (n_14, \A[715] );
  and g18 (n1011, n_14, \A[716] );
  not g19 (n_15, n1010);
  not g20 (n_16, n1011);
  and g21 (n1012, n_15, n_16);
  not g22 (n_18, n1012);
  and g23 (n1013, \A[717] , n_18);
  not g24 (n_19, n1009);
  not g25 (n_20, n1013);
  and g26 (n1014, n_19, n_20);
  not g27 (n_21, n1014);
  and g28 (n1015, n1008, n_21);
  not g29 (n_22, n1008);
  and g30 (n1016, n_22, n1014);
  and g31 (n1017, \A[717] , n_15);
  and g32 (n1018, n_16, n1017);
  not g33 (n_23, \A[717] );
  and g34 (n1019, n_23, n_18);
  not g35 (n_24, n1018);
  not g36 (n_25, n1019);
  and g37 (n1020, n_24, n_25);
  and g38 (n1021, \A[720] , n_5);
  and g39 (n1022, n_6, n1021);
  not g40 (n_26, \A[720] );
  and g41 (n1023, n_26, n_8);
  not g42 (n_27, n1022);
  not g43 (n_28, n1023);
  and g44 (n1024, n_27, n_28);
  not g45 (n_29, n1020);
  not g46 (n_30, n1024);
  and g47 (n1025, n_29, n_30);
  not g48 (n_31, n1016);
  and g49 (n1026, n_31, n1025);
  not g50 (n_32, n1015);
  and g51 (n1027, n_32, n1026);
  and g52 (n1028, n_32, n_31);
  not g53 (n_33, n1025);
  not g54 (n_34, n1028);
  and g55 (n1029, n_33, n_34);
  not g56 (n_35, n1027);
  not g57 (n_36, n1029);
  and g58 (n1030, n_35, n_36);
  and g59 (n1031, n_29, n1024);
  and g60 (n1032, n1020, n_30);
  not g61 (n_37, n1031);
  not g62 (n_38, n1032);
  and g63 (n1033, n_37, n_38);
  and g64 (n1034, n1025, n_34);
  and g65 (n1035, n_22, n_21);
  not g66 (n_39, n1034);
  not g67 (n_40, n1035);
  and g68 (n1036, n_39, n_40);
  not g69 (n_41, n1033);
  not g70 (n_42, n1036);
  and g71 (n1037, n_41, n_42);
  not g72 (n_43, n1030);
  not g73 (n_44, n1037);
  and g74 (n1038, n_43, n_44);
  and g75 (n1039, n_43, n_42);
  and g76 (n1040, \A[724] , \A[725] );
  not g77 (n_47, \A[725] );
  and g78 (n1041, \A[724] , n_47);
  not g79 (n_48, \A[724] );
  and g80 (n1042, n_48, \A[725] );
  not g81 (n_49, n1041);
  not g82 (n_50, n1042);
  and g83 (n1043, n_49, n_50);
  not g84 (n_52, n1043);
  and g85 (n1044, \A[726] , n_52);
  not g86 (n_53, n1040);
  not g87 (n_54, n1044);
  and g88 (n1045, n_53, n_54);
  and g89 (n1046, \A[721] , \A[722] );
  not g90 (n_57, \A[722] );
  and g91 (n1047, \A[721] , n_57);
  not g92 (n_58, \A[721] );
  and g93 (n1048, n_58, \A[722] );
  not g94 (n_59, n1047);
  not g95 (n_60, n1048);
  and g96 (n1049, n_59, n_60);
  not g97 (n_62, n1049);
  and g98 (n1050, \A[723] , n_62);
  not g99 (n_63, n1046);
  not g100 (n_64, n1050);
  and g101 (n1051, n_63, n_64);
  not g102 (n_65, n1045);
  and g103 (n1052, n_65, n1051);
  not g104 (n_66, n1051);
  and g105 (n1053, n1045, n_66);
  not g106 (n_67, n1052);
  not g107 (n_68, n1053);
  and g108 (n1054, n_67, n_68);
  and g109 (n1055, \A[723] , n_59);
  and g110 (n1056, n_60, n1055);
  not g111 (n_69, \A[723] );
  and g112 (n1057, n_69, n_62);
  not g113 (n_70, n1056);
  not g114 (n_71, n1057);
  and g115 (n1058, n_70, n_71);
  and g116 (n1059, \A[726] , n_49);
  and g117 (n1060, n_50, n1059);
  not g118 (n_72, \A[726] );
  and g119 (n1061, n_72, n_52);
  not g120 (n_73, n1060);
  not g121 (n_74, n1061);
  and g122 (n1062, n_73, n_74);
  not g123 (n_75, n1058);
  not g124 (n_76, n1062);
  and g125 (n1063, n_75, n_76);
  not g126 (n_77, n1054);
  and g127 (n1064, n_77, n1063);
  and g128 (n1065, n_65, n_66);
  not g129 (n_78, n1064);
  not g130 (n_79, n1065);
  and g131 (n1066, n_78, n_79);
  and g132 (n1067, n_67, n1063);
  and g133 (n1068, n_68, n1067);
  not g134 (n_80, n1063);
  and g135 (n1069, n_77, n_80);
  not g136 (n_81, n1068);
  not g137 (n_82, n1069);
  and g138 (n1070, n_81, n_82);
  not g139 (n_83, n1066);
  not g140 (n_84, n1070);
  and g141 (n1071, n_83, n_84);
  and g142 (n1072, n_75, n1062);
  and g143 (n1073, n1058, n_76);
  not g144 (n_85, n1072);
  not g145 (n_86, n1073);
  and g146 (n1074, n_85, n_86);
  not g147 (n_87, n1074);
  and g148 (n1075, n_41, n_87);
  not g149 (n_88, n1071);
  and g150 (n1076, n_88, n1075);
  not g151 (n_89, n1039);
  and g152 (n1077, n_89, n1076);
  and g153 (n1078, n_83, n_87);
  not g154 (n_90, n1078);
  and g155 (n1079, n_84, n_90);
  not g156 (n_91, n1077);
  not g157 (n_92, n1079);
  and g158 (n1080, n_91, n_92);
  not g163 (n_93, n1080);
  not g164 (n_94, n1084);
  and g165 (n1085, n_93, n_94);
  not g166 (n_95, n1085);
  and g167 (n1086, n1038, n_95);
  and g168 (n1087, n_91, n1079);
  and g169 (n1088, n1077, n_92);
  not g170 (n_96, n1087);
  not g171 (n_97, n1088);
  and g172 (n1089, n_96, n_97);
  not g173 (n_98, n1038);
  not g174 (n_99, n1089);
  and g175 (n1090, n_98, n_99);
  and g176 (n1091, n_88, n_87);
  and g177 (n1092, n_41, n_89);
  not g178 (n_100, n1091);
  and g179 (n1093, n_100, n1092);
  not g180 (n_101, n1092);
  and g181 (n1094, n1091, n_101);
  not g182 (n_102, n1093);
  not g183 (n_103, n1094);
  and g184 (n1095, n_102, n_103);
  not g185 (n_105, \A[709] );
  and g186 (n1096, n_105, \A[710] );
  not g187 (n_107, \A[710] );
  and g188 (n1097, \A[709] , n_107);
  not g189 (n_109, n1097);
  and g190 (n1098, \A[711] , n_109);
  not g191 (n_110, n1096);
  and g192 (n1099, n_110, n1098);
  and g193 (n1100, n_110, n_109);
  not g194 (n_111, \A[711] );
  not g195 (n_112, n1100);
  and g196 (n1101, n_111, n_112);
  not g197 (n_113, n1099);
  not g198 (n_114, n1101);
  and g199 (n1102, n_113, n_114);
  not g200 (n_116, \A[712] );
  and g201 (n1103, n_116, \A[713] );
  not g202 (n_118, \A[713] );
  and g203 (n1104, \A[712] , n_118);
  not g204 (n_120, n1104);
  and g205 (n1105, \A[714] , n_120);
  not g206 (n_121, n1103);
  and g207 (n1106, n_121, n1105);
  and g208 (n1107, n_121, n_120);
  not g209 (n_122, \A[714] );
  not g210 (n_123, n1107);
  and g211 (n1108, n_122, n_123);
  not g212 (n_124, n1106);
  not g213 (n_125, n1108);
  and g214 (n1109, n_124, n_125);
  not g215 (n_126, n1102);
  and g216 (n1110, n_126, n1109);
  not g217 (n_127, n1109);
  and g218 (n1111, n1102, n_127);
  not g219 (n_128, n1110);
  not g220 (n_129, n1111);
  and g221 (n1112, n_128, n_129);
  and g222 (n1113, \A[712] , \A[713] );
  and g223 (n1114, \A[714] , n_123);
  not g224 (n_130, n1113);
  not g225 (n_131, n1114);
  and g226 (n1115, n_130, n_131);
  and g227 (n1116, \A[709] , \A[710] );
  and g228 (n1117, \A[711] , n_112);
  not g229 (n_132, n1116);
  not g230 (n_133, n1117);
  and g231 (n1118, n_132, n_133);
  not g232 (n_134, n1115);
  and g233 (n1119, n_134, n1118);
  not g234 (n_135, n1118);
  and g235 (n1120, n1115, n_135);
  not g236 (n_136, n1119);
  not g237 (n_137, n1120);
  and g238 (n1121, n_136, n_137);
  and g239 (n1122, n_126, n_127);
  not g240 (n_138, n1121);
  and g241 (n1123, n_138, n1122);
  and g242 (n1124, n_134, n_135);
  not g243 (n_139, n1123);
  not g244 (n_140, n1124);
  and g245 (n1125, n_139, n_140);
  and g246 (n1126, n_136, n1122);
  and g247 (n1127, n_137, n1126);
  not g248 (n_141, n1122);
  and g249 (n1128, n_138, n_141);
  not g250 (n_142, n1127);
  not g251 (n_143, n1128);
  and g252 (n1129, n_142, n_143);
  not g253 (n_144, n1125);
  not g254 (n_145, n1129);
  and g255 (n1130, n_144, n_145);
  not g256 (n_146, n1112);
  not g257 (n_147, n1130);
  and g258 (n1131, n_146, n_147);
  not g259 (n_149, \A[703] );
  and g260 (n1132, n_149, \A[704] );
  not g261 (n_151, \A[704] );
  and g262 (n1133, \A[703] , n_151);
  not g263 (n_153, n1133);
  and g264 (n1134, \A[705] , n_153);
  not g265 (n_154, n1132);
  and g266 (n1135, n_154, n1134);
  and g267 (n1136, n_154, n_153);
  not g268 (n_155, \A[705] );
  not g269 (n_156, n1136);
  and g270 (n1137, n_155, n_156);
  not g271 (n_157, n1135);
  not g272 (n_158, n1137);
  and g273 (n1138, n_157, n_158);
  not g274 (n_160, \A[706] );
  and g275 (n1139, n_160, \A[707] );
  not g276 (n_162, \A[707] );
  and g277 (n1140, \A[706] , n_162);
  not g278 (n_164, n1140);
  and g279 (n1141, \A[708] , n_164);
  not g280 (n_165, n1139);
  and g281 (n1142, n_165, n1141);
  and g282 (n1143, n_165, n_164);
  not g283 (n_166, \A[708] );
  not g284 (n_167, n1143);
  and g285 (n1144, n_166, n_167);
  not g286 (n_168, n1142);
  not g287 (n_169, n1144);
  and g288 (n1145, n_168, n_169);
  not g289 (n_170, n1138);
  and g290 (n1146, n_170, n1145);
  not g291 (n_171, n1145);
  and g292 (n1147, n1138, n_171);
  not g293 (n_172, n1146);
  not g294 (n_173, n1147);
  and g295 (n1148, n_172, n_173);
  and g296 (n1149, \A[706] , \A[707] );
  and g297 (n1150, \A[708] , n_167);
  not g298 (n_174, n1149);
  not g299 (n_175, n1150);
  and g300 (n1151, n_174, n_175);
  and g301 (n1152, \A[703] , \A[704] );
  and g302 (n1153, \A[705] , n_156);
  not g303 (n_176, n1152);
  not g304 (n_177, n1153);
  and g305 (n1154, n_176, n_177);
  not g306 (n_178, n1151);
  and g307 (n1155, n_178, n1154);
  not g308 (n_179, n1154);
  and g309 (n1156, n1151, n_179);
  not g310 (n_180, n1155);
  not g311 (n_181, n1156);
  and g312 (n1157, n_180, n_181);
  and g313 (n1158, n_170, n_171);
  not g314 (n_182, n1157);
  and g315 (n1159, n_182, n1158);
  and g316 (n1160, n_178, n_179);
  not g317 (n_183, n1159);
  not g318 (n_184, n1160);
  and g319 (n1161, n_183, n_184);
  and g320 (n1162, n_180, n1158);
  and g321 (n1163, n_181, n1162);
  not g322 (n_185, n1158);
  and g323 (n1164, n_182, n_185);
  not g324 (n_186, n1163);
  not g325 (n_187, n1164);
  and g326 (n1165, n_186, n_187);
  not g327 (n_188, n1161);
  not g328 (n_189, n1165);
  and g329 (n1166, n_188, n_189);
  not g330 (n_190, n1148);
  not g331 (n_191, n1166);
  and g332 (n1167, n_190, n_191);
  not g333 (n_192, n1131);
  and g334 (n1168, n_192, n1167);
  not g335 (n_193, n1167);
  and g336 (n1169, n1131, n_193);
  not g337 (n_194, n1168);
  not g338 (n_195, n1169);
  and g339 (n1170, n_194, n_195);
  not g340 (n_196, n1095);
  not g341 (n_197, n1170);
  and g342 (n1171, n_196, n_197);
  not g343 (n_198, n1090);
  and g344 (n1172, n_198, n1171);
  not g345 (n_199, n1086);
  and g346 (n1173, n_199, n1172);
  and g347 (n1174, n_199, n_198);
  not g348 (n_200, n1171);
  not g349 (n_201, n1174);
  and g350 (n1175, n_200, n_201);
  not g351 (n_202, n1173);
  not g352 (n_203, n1175);
  and g353 (n1176, n_202, n_203);
  and g354 (n1177, n_190, n_188);
  not g355 (n_204, n1177);
  and g356 (n1178, n_189, n_204);
  and g357 (n1179, n_146, n_190);
  and g358 (n1180, n_147, n1179);
  and g359 (n1181, n_191, n1180);
  and g360 (n1182, n_146, n_144);
  not g361 (n_205, n1182);
  and g362 (n1183, n_145, n_205);
  not g363 (n_206, n1181);
  and g364 (n1184, n_206, n1183);
  not g365 (n_207, n1183);
  and g366 (n1185, n1181, n_207);
  not g367 (n_208, n1184);
  not g368 (n_209, n1185);
  and g369 (n1186, n_208, n_209);
  not g370 (n_210, n1178);
  not g371 (n_211, n1186);
  and g372 (n1187, n_210, n_211);
  and g373 (n1188, n_206, n_207);
  not g378 (n_212, n1188);
  not g379 (n_213, n1192);
  and g380 (n1193, n_212, n_213);
  not g381 (n_214, n1193);
  and g382 (n1194, n1178, n_214);
  not g383 (n_215, n1187);
  not g384 (n_216, n1194);
  and g385 (n1195, n_215, n_216);
  not g386 (n_217, n1176);
  and g387 (n1196, n_217, n1195);
  and g388 (n1197, n_198, n_200);
  and g389 (n1198, n_199, n1197);
  and g390 (n1199, n1171, n_201);
  not g391 (n_218, n1198);
  not g392 (n_219, n1199);
  and g393 (n1200, n_218, n_219);
  not g394 (n_220, n1195);
  not g395 (n_221, n1200);
  and g396 (n1201, n_220, n_221);
  not g397 (n_222, n1196);
  not g398 (n_223, n1201);
  and g399 (n1202, n_222, n_223);
  and g400 (n1203, \A[730] , \A[731] );
  not g401 (n_226, \A[731] );
  and g402 (n1204, \A[730] , n_226);
  not g403 (n_227, \A[730] );
  and g404 (n1205, n_227, \A[731] );
  not g405 (n_228, n1204);
  not g406 (n_229, n1205);
  and g407 (n1206, n_228, n_229);
  not g408 (n_231, n1206);
  and g409 (n1207, \A[732] , n_231);
  not g410 (n_232, n1203);
  not g411 (n_233, n1207);
  and g412 (n1208, n_232, n_233);
  and g413 (n1209, \A[727] , \A[728] );
  not g414 (n_236, \A[728] );
  and g415 (n1210, \A[727] , n_236);
  not g416 (n_237, \A[727] );
  and g417 (n1211, n_237, \A[728] );
  not g418 (n_238, n1210);
  not g419 (n_239, n1211);
  and g420 (n1212, n_238, n_239);
  not g421 (n_241, n1212);
  and g422 (n1213, \A[729] , n_241);
  not g423 (n_242, n1209);
  not g424 (n_243, n1213);
  and g425 (n1214, n_242, n_243);
  not g426 (n_244, n1214);
  and g427 (n1215, n1208, n_244);
  not g428 (n_245, n1208);
  and g429 (n1216, n_245, n1214);
  and g430 (n1217, \A[729] , n_238);
  and g431 (n1218, n_239, n1217);
  not g432 (n_246, \A[729] );
  and g433 (n1219, n_246, n_241);
  not g434 (n_247, n1218);
  not g435 (n_248, n1219);
  and g436 (n1220, n_247, n_248);
  and g437 (n1221, \A[732] , n_228);
  and g438 (n1222, n_229, n1221);
  not g439 (n_249, \A[732] );
  and g440 (n1223, n_249, n_231);
  not g441 (n_250, n1222);
  not g442 (n_251, n1223);
  and g443 (n1224, n_250, n_251);
  not g444 (n_252, n1220);
  not g445 (n_253, n1224);
  and g446 (n1225, n_252, n_253);
  not g447 (n_254, n1216);
  and g448 (n1226, n_254, n1225);
  not g449 (n_255, n1215);
  and g450 (n1227, n_255, n1226);
  and g451 (n1228, n_255, n_254);
  not g452 (n_256, n1225);
  not g453 (n_257, n1228);
  and g454 (n1229, n_256, n_257);
  not g455 (n_258, n1227);
  not g456 (n_259, n1229);
  and g457 (n1230, n_258, n_259);
  and g458 (n1231, n_252, n1224);
  and g459 (n1232, n1220, n_253);
  not g460 (n_260, n1231);
  not g461 (n_261, n1232);
  and g462 (n1233, n_260, n_261);
  and g463 (n1234, n1225, n_257);
  and g464 (n1235, n_245, n_244);
  not g465 (n_262, n1234);
  not g466 (n_263, n1235);
  and g467 (n1236, n_262, n_263);
  not g468 (n_264, n1233);
  not g469 (n_265, n1236);
  and g470 (n1237, n_264, n_265);
  not g471 (n_266, n1230);
  not g472 (n_267, n1237);
  and g473 (n1238, n_266, n_267);
  and g474 (n1239, n_266, n_265);
  and g475 (n1240, \A[736] , \A[737] );
  not g476 (n_270, \A[737] );
  and g477 (n1241, \A[736] , n_270);
  not g478 (n_271, \A[736] );
  and g479 (n1242, n_271, \A[737] );
  not g480 (n_272, n1241);
  not g481 (n_273, n1242);
  and g482 (n1243, n_272, n_273);
  not g483 (n_275, n1243);
  and g484 (n1244, \A[738] , n_275);
  not g485 (n_276, n1240);
  not g486 (n_277, n1244);
  and g487 (n1245, n_276, n_277);
  and g488 (n1246, \A[733] , \A[734] );
  not g489 (n_280, \A[734] );
  and g490 (n1247, \A[733] , n_280);
  not g491 (n_281, \A[733] );
  and g492 (n1248, n_281, \A[734] );
  not g493 (n_282, n1247);
  not g494 (n_283, n1248);
  and g495 (n1249, n_282, n_283);
  not g496 (n_285, n1249);
  and g497 (n1250, \A[735] , n_285);
  not g498 (n_286, n1246);
  not g499 (n_287, n1250);
  and g500 (n1251, n_286, n_287);
  not g501 (n_288, n1245);
  and g502 (n1252, n_288, n1251);
  not g503 (n_289, n1251);
  and g504 (n1253, n1245, n_289);
  not g505 (n_290, n1252);
  not g506 (n_291, n1253);
  and g507 (n1254, n_290, n_291);
  and g508 (n1255, \A[735] , n_282);
  and g509 (n1256, n_283, n1255);
  not g510 (n_292, \A[735] );
  and g511 (n1257, n_292, n_285);
  not g512 (n_293, n1256);
  not g513 (n_294, n1257);
  and g514 (n1258, n_293, n_294);
  and g515 (n1259, \A[738] , n_272);
  and g516 (n1260, n_273, n1259);
  not g517 (n_295, \A[738] );
  and g518 (n1261, n_295, n_275);
  not g519 (n_296, n1260);
  not g520 (n_297, n1261);
  and g521 (n1262, n_296, n_297);
  not g522 (n_298, n1258);
  not g523 (n_299, n1262);
  and g524 (n1263, n_298, n_299);
  not g525 (n_300, n1254);
  and g526 (n1264, n_300, n1263);
  and g527 (n1265, n_288, n_289);
  not g528 (n_301, n1264);
  not g529 (n_302, n1265);
  and g530 (n1266, n_301, n_302);
  and g531 (n1267, n_290, n1263);
  and g532 (n1268, n_291, n1267);
  not g533 (n_303, n1263);
  and g534 (n1269, n_300, n_303);
  not g535 (n_304, n1268);
  not g536 (n_305, n1269);
  and g537 (n1270, n_304, n_305);
  not g538 (n_306, n1266);
  not g539 (n_307, n1270);
  and g540 (n1271, n_306, n_307);
  and g541 (n1272, n_298, n1262);
  and g542 (n1273, n1258, n_299);
  not g543 (n_308, n1272);
  not g544 (n_309, n1273);
  and g545 (n1274, n_308, n_309);
  not g546 (n_310, n1274);
  and g547 (n1275, n_264, n_310);
  not g548 (n_311, n1271);
  and g549 (n1276, n_311, n1275);
  not g550 (n_312, n1239);
  and g551 (n1277, n_312, n1276);
  and g552 (n1278, n_306, n_310);
  not g553 (n_313, n1278);
  and g554 (n1279, n_307, n_313);
  not g555 (n_314, n1277);
  and g556 (n1280, n_314, n1279);
  not g557 (n_315, n1279);
  and g558 (n1281, n1277, n_315);
  not g559 (n_316, n1280);
  not g560 (n_317, n1281);
  and g561 (n1282, n_316, n_317);
  not g562 (n_318, n1238);
  not g563 (n_319, n1282);
  and g564 (n1283, n_318, n_319);
  and g565 (n1284, n_314, n_315);
  not g570 (n_320, n1284);
  not g571 (n_321, n1288);
  and g572 (n1289, n_320, n_321);
  not g573 (n_322, n1289);
  and g574 (n1290, n1238, n_322);
  not g575 (n_323, n1283);
  not g576 (n_324, n1290);
  and g577 (n1291, n_323, n_324);
  and g578 (n1292, \A[742] , \A[743] );
  not g579 (n_327, \A[743] );
  and g580 (n1293, \A[742] , n_327);
  not g581 (n_328, \A[742] );
  and g582 (n1294, n_328, \A[743] );
  not g583 (n_329, n1293);
  not g584 (n_330, n1294);
  and g585 (n1295, n_329, n_330);
  not g586 (n_332, n1295);
  and g587 (n1296, \A[744] , n_332);
  not g588 (n_333, n1292);
  not g589 (n_334, n1296);
  and g590 (n1297, n_333, n_334);
  and g591 (n1298, \A[739] , \A[740] );
  not g592 (n_337, \A[740] );
  and g593 (n1299, \A[739] , n_337);
  not g594 (n_338, \A[739] );
  and g595 (n1300, n_338, \A[740] );
  not g596 (n_339, n1299);
  not g597 (n_340, n1300);
  and g598 (n1301, n_339, n_340);
  not g599 (n_342, n1301);
  and g600 (n1302, \A[741] , n_342);
  not g601 (n_343, n1298);
  not g602 (n_344, n1302);
  and g603 (n1303, n_343, n_344);
  not g604 (n_345, n1303);
  and g605 (n1304, n1297, n_345);
  not g606 (n_346, n1297);
  and g607 (n1305, n_346, n1303);
  and g608 (n1306, \A[741] , n_339);
  and g609 (n1307, n_340, n1306);
  not g610 (n_347, \A[741] );
  and g611 (n1308, n_347, n_342);
  not g612 (n_348, n1307);
  not g613 (n_349, n1308);
  and g614 (n1309, n_348, n_349);
  and g615 (n1310, \A[744] , n_329);
  and g616 (n1311, n_330, n1310);
  not g617 (n_350, \A[744] );
  and g618 (n1312, n_350, n_332);
  not g619 (n_351, n1311);
  not g620 (n_352, n1312);
  and g621 (n1313, n_351, n_352);
  not g622 (n_353, n1309);
  not g623 (n_354, n1313);
  and g624 (n1314, n_353, n_354);
  not g625 (n_355, n1305);
  and g626 (n1315, n_355, n1314);
  not g627 (n_356, n1304);
  and g628 (n1316, n_356, n1315);
  and g629 (n1317, n_356, n_355);
  not g630 (n_357, n1314);
  not g631 (n_358, n1317);
  and g632 (n1318, n_357, n_358);
  not g633 (n_359, n1316);
  not g634 (n_360, n1318);
  and g635 (n1319, n_359, n_360);
  and g636 (n1320, n_353, n1313);
  and g637 (n1321, n1309, n_354);
  not g638 (n_361, n1320);
  not g639 (n_362, n1321);
  and g640 (n1322, n_361, n_362);
  and g641 (n1323, n1314, n_358);
  and g642 (n1324, n_346, n_345);
  not g643 (n_363, n1323);
  not g644 (n_364, n1324);
  and g645 (n1325, n_363, n_364);
  not g646 (n_365, n1322);
  not g647 (n_366, n1325);
  and g648 (n1326, n_365, n_366);
  not g649 (n_367, n1319);
  not g650 (n_368, n1326);
  and g651 (n1327, n_367, n_368);
  and g652 (n1328, n_367, n_366);
  and g653 (n1329, \A[748] , \A[749] );
  not g654 (n_371, \A[749] );
  and g655 (n1330, \A[748] , n_371);
  not g656 (n_372, \A[748] );
  and g657 (n1331, n_372, \A[749] );
  not g658 (n_373, n1330);
  not g659 (n_374, n1331);
  and g660 (n1332, n_373, n_374);
  not g661 (n_376, n1332);
  and g662 (n1333, \A[750] , n_376);
  not g663 (n_377, n1329);
  not g664 (n_378, n1333);
  and g665 (n1334, n_377, n_378);
  and g666 (n1335, \A[745] , \A[746] );
  not g667 (n_381, \A[746] );
  and g668 (n1336, \A[745] , n_381);
  not g669 (n_382, \A[745] );
  and g670 (n1337, n_382, \A[746] );
  not g671 (n_383, n1336);
  not g672 (n_384, n1337);
  and g673 (n1338, n_383, n_384);
  not g674 (n_386, n1338);
  and g675 (n1339, \A[747] , n_386);
  not g676 (n_387, n1335);
  not g677 (n_388, n1339);
  and g678 (n1340, n_387, n_388);
  not g679 (n_389, n1334);
  and g680 (n1341, n_389, n1340);
  not g681 (n_390, n1340);
  and g682 (n1342, n1334, n_390);
  not g683 (n_391, n1341);
  not g684 (n_392, n1342);
  and g685 (n1343, n_391, n_392);
  and g686 (n1344, \A[747] , n_383);
  and g687 (n1345, n_384, n1344);
  not g688 (n_393, \A[747] );
  and g689 (n1346, n_393, n_386);
  not g690 (n_394, n1345);
  not g691 (n_395, n1346);
  and g692 (n1347, n_394, n_395);
  and g693 (n1348, \A[750] , n_373);
  and g694 (n1349, n_374, n1348);
  not g695 (n_396, \A[750] );
  and g696 (n1350, n_396, n_376);
  not g697 (n_397, n1349);
  not g698 (n_398, n1350);
  and g699 (n1351, n_397, n_398);
  not g700 (n_399, n1347);
  not g701 (n_400, n1351);
  and g702 (n1352, n_399, n_400);
  not g703 (n_401, n1343);
  and g704 (n1353, n_401, n1352);
  and g705 (n1354, n_389, n_390);
  not g706 (n_402, n1353);
  not g707 (n_403, n1354);
  and g708 (n1355, n_402, n_403);
  and g709 (n1356, n_391, n1352);
  and g710 (n1357, n_392, n1356);
  not g711 (n_404, n1352);
  and g712 (n1358, n_401, n_404);
  not g713 (n_405, n1357);
  not g714 (n_406, n1358);
  and g715 (n1359, n_405, n_406);
  not g716 (n_407, n1355);
  not g717 (n_408, n1359);
  and g718 (n1360, n_407, n_408);
  and g719 (n1361, n_399, n1351);
  and g720 (n1362, n1347, n_400);
  not g721 (n_409, n1361);
  not g722 (n_410, n1362);
  and g723 (n1363, n_409, n_410);
  not g724 (n_411, n1363);
  and g725 (n1364, n_365, n_411);
  not g726 (n_412, n1360);
  and g727 (n1365, n_412, n1364);
  not g728 (n_413, n1328);
  and g729 (n1366, n_413, n1365);
  and g730 (n1367, n_407, n_411);
  not g731 (n_414, n1367);
  and g732 (n1368, n_408, n_414);
  not g733 (n_415, n1366);
  not g734 (n_416, n1368);
  and g735 (n1369, n_415, n_416);
  not g740 (n_417, n1369);
  not g741 (n_418, n1373);
  and g742 (n1374, n_417, n_418);
  not g743 (n_419, n1374);
  and g744 (n1375, n1327, n_419);
  and g745 (n1376, n_415, n1368);
  and g746 (n1377, n1366, n_416);
  not g747 (n_420, n1376);
  not g748 (n_421, n1377);
  and g749 (n1378, n_420, n_421);
  not g750 (n_422, n1327);
  not g751 (n_423, n1378);
  and g752 (n1379, n_422, n_423);
  and g753 (n1380, n_412, n_411);
  and g754 (n1381, n_365, n_413);
  not g755 (n_424, n1380);
  and g756 (n1382, n_424, n1381);
  not g757 (n_425, n1381);
  and g758 (n1383, n1380, n_425);
  not g759 (n_426, n1382);
  not g760 (n_427, n1383);
  and g761 (n1384, n_426, n_427);
  and g762 (n1385, n_311, n_310);
  and g763 (n1386, n_264, n_312);
  not g764 (n_428, n1385);
  and g765 (n1387, n_428, n1386);
  not g766 (n_429, n1386);
  and g767 (n1388, n1385, n_429);
  not g768 (n_430, n1387);
  not g769 (n_431, n1388);
  and g770 (n1389, n_430, n_431);
  not g771 (n_432, n1384);
  not g772 (n_433, n1389);
  and g773 (n1390, n_432, n_433);
  not g774 (n_434, n1379);
  not g775 (n_435, n1390);
  and g776 (n1391, n_434, n_435);
  not g777 (n_436, n1375);
  and g778 (n1392, n_436, n1391);
  and g779 (n1393, n_436, n_434);
  not g780 (n_437, n1393);
  and g781 (n1394, n1390, n_437);
  not g782 (n_438, n1392);
  not g783 (n_439, n1394);
  and g784 (n1395, n_438, n_439);
  not g785 (n_440, n1291);
  not g786 (n_441, n1395);
  and g787 (n1396, n_440, n_441);
  and g788 (n1397, n_434, n1390);
  and g789 (n1398, n_436, n1397);
  and g790 (n1399, n_435, n_437);
  not g791 (n_442, n1398);
  not g792 (n_443, n1399);
  and g793 (n1400, n_442, n_443);
  not g794 (n_444, n1400);
  and g795 (n1401, n1291, n_444);
  and g796 (n1402, n_432, n1389);
  and g797 (n1403, n1384, n_433);
  not g798 (n_445, n1402);
  not g799 (n_446, n1403);
  and g800 (n1404, n_445, n_446);
  and g801 (n1405, n_196, n1170);
  and g802 (n1406, n1095, n_197);
  not g803 (n_447, n1405);
  not g804 (n_448, n1406);
  and g805 (n1407, n_447, n_448);
  not g806 (n_449, n1404);
  not g807 (n_450, n1407);
  and g808 (n1408, n_449, n_450);
  not g809 (n_451, n1401);
  not g810 (n_452, n1408);
  and g811 (n1409, n_451, n_452);
  not g812 (n_453, n1396);
  and g813 (n1410, n_453, n1409);
  and g814 (n1411, n_453, n_451);
  not g815 (n_454, n1411);
  and g816 (n1412, n1408, n_454);
  not g817 (n_455, n1410);
  not g818 (n_456, n1412);
  and g819 (n1413, n_455, n_456);
  not g820 (n_457, n1202);
  not g821 (n_458, n1413);
  and g822 (n1414, n_457, n_458);
  and g823 (n1415, n_451, n1408);
  and g824 (n1416, n_453, n1415);
  and g825 (n1417, n_452, n_454);
  not g826 (n_459, n1416);
  not g827 (n_460, n1417);
  and g828 (n1418, n_459, n_460);
  not g829 (n_461, n1418);
  and g830 (n1419, n1202, n_461);
  and g831 (n1420, n_449, n1407);
  and g832 (n1421, n1404, n_450);
  not g833 (n_462, n1420);
  not g834 (n_463, n1421);
  and g835 (n1422, n_462, n_463);
  not g836 (n_465, \A[697] );
  and g837 (n1423, n_465, \A[698] );
  not g838 (n_467, \A[698] );
  and g839 (n1424, \A[697] , n_467);
  not g840 (n_469, n1424);
  and g841 (n1425, \A[699] , n_469);
  not g842 (n_470, n1423);
  and g843 (n1426, n_470, n1425);
  and g844 (n1427, n_470, n_469);
  not g845 (n_471, \A[699] );
  not g846 (n_472, n1427);
  and g847 (n1428, n_471, n_472);
  not g848 (n_473, n1426);
  not g849 (n_474, n1428);
  and g850 (n1429, n_473, n_474);
  not g851 (n_476, \A[700] );
  and g852 (n1430, n_476, \A[701] );
  not g853 (n_478, \A[701] );
  and g854 (n1431, \A[700] , n_478);
  not g855 (n_480, n1431);
  and g856 (n1432, \A[702] , n_480);
  not g857 (n_481, n1430);
  and g858 (n1433, n_481, n1432);
  and g859 (n1434, n_481, n_480);
  not g860 (n_482, \A[702] );
  not g861 (n_483, n1434);
  and g862 (n1435, n_482, n_483);
  not g863 (n_484, n1433);
  not g864 (n_485, n1435);
  and g865 (n1436, n_484, n_485);
  not g866 (n_486, n1429);
  and g867 (n1437, n_486, n1436);
  not g868 (n_487, n1436);
  and g869 (n1438, n1429, n_487);
  not g870 (n_488, n1437);
  not g871 (n_489, n1438);
  and g872 (n1439, n_488, n_489);
  and g873 (n1440, \A[700] , \A[701] );
  and g874 (n1441, \A[702] , n_483);
  not g875 (n_490, n1440);
  not g876 (n_491, n1441);
  and g877 (n1442, n_490, n_491);
  and g878 (n1443, \A[697] , \A[698] );
  and g879 (n1444, \A[699] , n_472);
  not g880 (n_492, n1443);
  not g881 (n_493, n1444);
  and g882 (n1445, n_492, n_493);
  not g883 (n_494, n1442);
  and g884 (n1446, n_494, n1445);
  not g885 (n_495, n1445);
  and g886 (n1447, n1442, n_495);
  not g887 (n_496, n1446);
  not g888 (n_497, n1447);
  and g889 (n1448, n_496, n_497);
  and g890 (n1449, n_486, n_487);
  not g891 (n_498, n1448);
  and g892 (n1450, n_498, n1449);
  and g893 (n1451, n_494, n_495);
  not g894 (n_499, n1450);
  not g895 (n_500, n1451);
  and g896 (n1452, n_499, n_500);
  and g897 (n1453, n_496, n1449);
  and g898 (n1454, n_497, n1453);
  not g899 (n_501, n1449);
  and g900 (n1455, n_498, n_501);
  not g901 (n_502, n1454);
  not g902 (n_503, n1455);
  and g903 (n1456, n_502, n_503);
  not g904 (n_504, n1452);
  not g905 (n_505, n1456);
  and g906 (n1457, n_504, n_505);
  not g907 (n_506, n1439);
  not g908 (n_507, n1457);
  and g909 (n1458, n_506, n_507);
  not g910 (n_509, \A[691] );
  and g911 (n1459, n_509, \A[692] );
  not g912 (n_511, \A[692] );
  and g913 (n1460, \A[691] , n_511);
  not g914 (n_513, n1460);
  and g915 (n1461, \A[693] , n_513);
  not g916 (n_514, n1459);
  and g917 (n1462, n_514, n1461);
  and g918 (n1463, n_514, n_513);
  not g919 (n_515, \A[693] );
  not g920 (n_516, n1463);
  and g921 (n1464, n_515, n_516);
  not g922 (n_517, n1462);
  not g923 (n_518, n1464);
  and g924 (n1465, n_517, n_518);
  not g925 (n_520, \A[694] );
  and g926 (n1466, n_520, \A[695] );
  not g927 (n_522, \A[695] );
  and g928 (n1467, \A[694] , n_522);
  not g929 (n_524, n1467);
  and g930 (n1468, \A[696] , n_524);
  not g931 (n_525, n1466);
  and g932 (n1469, n_525, n1468);
  and g933 (n1470, n_525, n_524);
  not g934 (n_526, \A[696] );
  not g935 (n_527, n1470);
  and g936 (n1471, n_526, n_527);
  not g937 (n_528, n1469);
  not g938 (n_529, n1471);
  and g939 (n1472, n_528, n_529);
  not g940 (n_530, n1465);
  and g941 (n1473, n_530, n1472);
  not g942 (n_531, n1472);
  and g943 (n1474, n1465, n_531);
  not g944 (n_532, n1473);
  not g945 (n_533, n1474);
  and g946 (n1475, n_532, n_533);
  and g947 (n1476, \A[694] , \A[695] );
  and g948 (n1477, \A[696] , n_527);
  not g949 (n_534, n1476);
  not g950 (n_535, n1477);
  and g951 (n1478, n_534, n_535);
  and g952 (n1479, \A[691] , \A[692] );
  and g953 (n1480, \A[693] , n_516);
  not g954 (n_536, n1479);
  not g955 (n_537, n1480);
  and g956 (n1481, n_536, n_537);
  not g957 (n_538, n1478);
  and g958 (n1482, n_538, n1481);
  not g959 (n_539, n1481);
  and g960 (n1483, n1478, n_539);
  not g961 (n_540, n1482);
  not g962 (n_541, n1483);
  and g963 (n1484, n_540, n_541);
  and g964 (n1485, n_530, n_531);
  not g965 (n_542, n1484);
  and g966 (n1486, n_542, n1485);
  and g967 (n1487, n_538, n_539);
  not g968 (n_543, n1486);
  not g969 (n_544, n1487);
  and g970 (n1488, n_543, n_544);
  and g971 (n1489, n_540, n1485);
  and g972 (n1490, n_541, n1489);
  not g973 (n_545, n1485);
  and g974 (n1491, n_542, n_545);
  not g975 (n_546, n1490);
  not g976 (n_547, n1491);
  and g977 (n1492, n_546, n_547);
  not g978 (n_548, n1488);
  not g979 (n_549, n1492);
  and g980 (n1493, n_548, n_549);
  not g981 (n_550, n1475);
  not g982 (n_551, n1493);
  and g983 (n1494, n_550, n_551);
  not g984 (n_552, n1458);
  and g985 (n1495, n_552, n1494);
  not g986 (n_553, n1494);
  and g987 (n1496, n1458, n_553);
  not g988 (n_554, n1495);
  not g989 (n_555, n1496);
  and g990 (n1497, n_554, n_555);
  not g991 (n_557, \A[685] );
  and g992 (n1498, n_557, \A[686] );
  not g993 (n_559, \A[686] );
  and g994 (n1499, \A[685] , n_559);
  not g995 (n_561, n1499);
  and g996 (n1500, \A[687] , n_561);
  not g997 (n_562, n1498);
  and g998 (n1501, n_562, n1500);
  and g999 (n1502, n_562, n_561);
  not g1000 (n_563, \A[687] );
  not g1001 (n_564, n1502);
  and g1002 (n1503, n_563, n_564);
  not g1003 (n_565, n1501);
  not g1004 (n_566, n1503);
  and g1005 (n1504, n_565, n_566);
  not g1006 (n_568, \A[688] );
  and g1007 (n1505, n_568, \A[689] );
  not g1008 (n_570, \A[689] );
  and g1009 (n1506, \A[688] , n_570);
  not g1010 (n_572, n1506);
  and g1011 (n1507, \A[690] , n_572);
  not g1012 (n_573, n1505);
  and g1013 (n1508, n_573, n1507);
  and g1014 (n1509, n_573, n_572);
  not g1015 (n_574, \A[690] );
  not g1016 (n_575, n1509);
  and g1017 (n1510, n_574, n_575);
  not g1018 (n_576, n1508);
  not g1019 (n_577, n1510);
  and g1020 (n1511, n_576, n_577);
  not g1021 (n_578, n1504);
  and g1022 (n1512, n_578, n1511);
  not g1023 (n_579, n1511);
  and g1024 (n1513, n1504, n_579);
  not g1025 (n_580, n1512);
  not g1026 (n_581, n1513);
  and g1027 (n1514, n_580, n_581);
  and g1028 (n1515, \A[688] , \A[689] );
  and g1029 (n1516, \A[690] , n_575);
  not g1030 (n_582, n1515);
  not g1031 (n_583, n1516);
  and g1032 (n1517, n_582, n_583);
  and g1033 (n1518, \A[685] , \A[686] );
  and g1034 (n1519, \A[687] , n_564);
  not g1035 (n_584, n1518);
  not g1036 (n_585, n1519);
  and g1037 (n1520, n_584, n_585);
  not g1038 (n_586, n1517);
  and g1039 (n1521, n_586, n1520);
  not g1040 (n_587, n1520);
  and g1041 (n1522, n1517, n_587);
  not g1042 (n_588, n1521);
  not g1043 (n_589, n1522);
  and g1044 (n1523, n_588, n_589);
  and g1045 (n1524, n_578, n_579);
  not g1046 (n_590, n1523);
  and g1047 (n1525, n_590, n1524);
  and g1048 (n1526, n_586, n_587);
  not g1049 (n_591, n1525);
  not g1050 (n_592, n1526);
  and g1051 (n1527, n_591, n_592);
  and g1052 (n1528, n_588, n1524);
  and g1053 (n1529, n_589, n1528);
  not g1054 (n_593, n1524);
  and g1055 (n1530, n_590, n_593);
  not g1056 (n_594, n1529);
  not g1057 (n_595, n1530);
  and g1058 (n1531, n_594, n_595);
  not g1059 (n_596, n1527);
  not g1060 (n_597, n1531);
  and g1061 (n1532, n_596, n_597);
  not g1062 (n_598, n1514);
  not g1063 (n_599, n1532);
  and g1064 (n1533, n_598, n_599);
  not g1065 (n_601, \A[679] );
  and g1066 (n1534, n_601, \A[680] );
  not g1067 (n_603, \A[680] );
  and g1068 (n1535, \A[679] , n_603);
  not g1069 (n_605, n1535);
  and g1070 (n1536, \A[681] , n_605);
  not g1071 (n_606, n1534);
  and g1072 (n1537, n_606, n1536);
  and g1073 (n1538, n_606, n_605);
  not g1074 (n_607, \A[681] );
  not g1075 (n_608, n1538);
  and g1076 (n1539, n_607, n_608);
  not g1077 (n_609, n1537);
  not g1078 (n_610, n1539);
  and g1079 (n1540, n_609, n_610);
  not g1080 (n_612, \A[682] );
  and g1081 (n1541, n_612, \A[683] );
  not g1082 (n_614, \A[683] );
  and g1083 (n1542, \A[682] , n_614);
  not g1084 (n_616, n1542);
  and g1085 (n1543, \A[684] , n_616);
  not g1086 (n_617, n1541);
  and g1087 (n1544, n_617, n1543);
  and g1088 (n1545, n_617, n_616);
  not g1089 (n_618, \A[684] );
  not g1090 (n_619, n1545);
  and g1091 (n1546, n_618, n_619);
  not g1092 (n_620, n1544);
  not g1093 (n_621, n1546);
  and g1094 (n1547, n_620, n_621);
  not g1095 (n_622, n1540);
  and g1096 (n1548, n_622, n1547);
  not g1097 (n_623, n1547);
  and g1098 (n1549, n1540, n_623);
  not g1099 (n_624, n1548);
  not g1100 (n_625, n1549);
  and g1101 (n1550, n_624, n_625);
  and g1102 (n1551, \A[682] , \A[683] );
  and g1103 (n1552, \A[684] , n_619);
  not g1104 (n_626, n1551);
  not g1105 (n_627, n1552);
  and g1106 (n1553, n_626, n_627);
  and g1107 (n1554, \A[679] , \A[680] );
  and g1108 (n1555, \A[681] , n_608);
  not g1109 (n_628, n1554);
  not g1110 (n_629, n1555);
  and g1111 (n1556, n_628, n_629);
  not g1112 (n_630, n1553);
  and g1113 (n1557, n_630, n1556);
  not g1114 (n_631, n1556);
  and g1115 (n1558, n1553, n_631);
  not g1116 (n_632, n1557);
  not g1117 (n_633, n1558);
  and g1118 (n1559, n_632, n_633);
  and g1119 (n1560, n_622, n_623);
  not g1120 (n_634, n1559);
  and g1121 (n1561, n_634, n1560);
  and g1122 (n1562, n_630, n_631);
  not g1123 (n_635, n1561);
  not g1124 (n_636, n1562);
  and g1125 (n1563, n_635, n_636);
  and g1126 (n1564, n_632, n1560);
  and g1127 (n1565, n_633, n1564);
  not g1128 (n_637, n1560);
  and g1129 (n1566, n_634, n_637);
  not g1130 (n_638, n1565);
  not g1131 (n_639, n1566);
  and g1132 (n1567, n_638, n_639);
  not g1133 (n_640, n1563);
  not g1134 (n_641, n1567);
  and g1135 (n1568, n_640, n_641);
  not g1136 (n_642, n1550);
  not g1137 (n_643, n1568);
  and g1138 (n1569, n_642, n_643);
  not g1139 (n_644, n1533);
  and g1140 (n1570, n_644, n1569);
  not g1141 (n_645, n1569);
  and g1142 (n1571, n1533, n_645);
  not g1143 (n_646, n1570);
  not g1144 (n_647, n1571);
  and g1145 (n1572, n_646, n_647);
  not g1146 (n_648, n1497);
  and g1147 (n1573, n_648, n1572);
  not g1148 (n_649, n1572);
  and g1149 (n1574, n1497, n_649);
  not g1150 (n_650, n1573);
  not g1151 (n_651, n1574);
  and g1152 (n1575, n_650, n_651);
  not g1153 (n_653, \A[673] );
  and g1154 (n1576, n_653, \A[674] );
  not g1155 (n_655, \A[674] );
  and g1156 (n1577, \A[673] , n_655);
  not g1157 (n_657, n1577);
  and g1158 (n1578, \A[675] , n_657);
  not g1159 (n_658, n1576);
  and g1160 (n1579, n_658, n1578);
  and g1161 (n1580, n_658, n_657);
  not g1162 (n_659, \A[675] );
  not g1163 (n_660, n1580);
  and g1164 (n1581, n_659, n_660);
  not g1165 (n_661, n1579);
  not g1166 (n_662, n1581);
  and g1167 (n1582, n_661, n_662);
  not g1168 (n_664, \A[676] );
  and g1169 (n1583, n_664, \A[677] );
  not g1170 (n_666, \A[677] );
  and g1171 (n1584, \A[676] , n_666);
  not g1172 (n_668, n1584);
  and g1173 (n1585, \A[678] , n_668);
  not g1174 (n_669, n1583);
  and g1175 (n1586, n_669, n1585);
  and g1176 (n1587, n_669, n_668);
  not g1177 (n_670, \A[678] );
  not g1178 (n_671, n1587);
  and g1179 (n1588, n_670, n_671);
  not g1180 (n_672, n1586);
  not g1181 (n_673, n1588);
  and g1182 (n1589, n_672, n_673);
  not g1183 (n_674, n1582);
  and g1184 (n1590, n_674, n1589);
  not g1185 (n_675, n1589);
  and g1186 (n1591, n1582, n_675);
  not g1187 (n_676, n1590);
  not g1188 (n_677, n1591);
  and g1189 (n1592, n_676, n_677);
  and g1190 (n1593, \A[676] , \A[677] );
  and g1191 (n1594, \A[678] , n_671);
  not g1192 (n_678, n1593);
  not g1193 (n_679, n1594);
  and g1194 (n1595, n_678, n_679);
  and g1195 (n1596, \A[673] , \A[674] );
  and g1196 (n1597, \A[675] , n_660);
  not g1197 (n_680, n1596);
  not g1198 (n_681, n1597);
  and g1199 (n1598, n_680, n_681);
  not g1200 (n_682, n1595);
  and g1201 (n1599, n_682, n1598);
  not g1202 (n_683, n1598);
  and g1203 (n1600, n1595, n_683);
  not g1204 (n_684, n1599);
  not g1205 (n_685, n1600);
  and g1206 (n1601, n_684, n_685);
  and g1207 (n1602, n_674, n_675);
  not g1208 (n_686, n1601);
  and g1209 (n1603, n_686, n1602);
  and g1210 (n1604, n_682, n_683);
  not g1211 (n_687, n1603);
  not g1212 (n_688, n1604);
  and g1213 (n1605, n_687, n_688);
  and g1214 (n1606, n_684, n1602);
  and g1215 (n1607, n_685, n1606);
  not g1216 (n_689, n1602);
  and g1217 (n1608, n_686, n_689);
  not g1218 (n_690, n1607);
  not g1219 (n_691, n1608);
  and g1220 (n1609, n_690, n_691);
  not g1221 (n_692, n1605);
  not g1222 (n_693, n1609);
  and g1223 (n1610, n_692, n_693);
  not g1224 (n_694, n1592);
  not g1225 (n_695, n1610);
  and g1226 (n1611, n_694, n_695);
  not g1227 (n_697, \A[667] );
  and g1228 (n1612, n_697, \A[668] );
  not g1229 (n_699, \A[668] );
  and g1230 (n1613, \A[667] , n_699);
  not g1231 (n_701, n1613);
  and g1232 (n1614, \A[669] , n_701);
  not g1233 (n_702, n1612);
  and g1234 (n1615, n_702, n1614);
  and g1235 (n1616, n_702, n_701);
  not g1236 (n_703, \A[669] );
  not g1237 (n_704, n1616);
  and g1238 (n1617, n_703, n_704);
  not g1239 (n_705, n1615);
  not g1240 (n_706, n1617);
  and g1241 (n1618, n_705, n_706);
  not g1242 (n_708, \A[670] );
  and g1243 (n1619, n_708, \A[671] );
  not g1244 (n_710, \A[671] );
  and g1245 (n1620, \A[670] , n_710);
  not g1246 (n_712, n1620);
  and g1247 (n1621, \A[672] , n_712);
  not g1248 (n_713, n1619);
  and g1249 (n1622, n_713, n1621);
  and g1250 (n1623, n_713, n_712);
  not g1251 (n_714, \A[672] );
  not g1252 (n_715, n1623);
  and g1253 (n1624, n_714, n_715);
  not g1254 (n_716, n1622);
  not g1255 (n_717, n1624);
  and g1256 (n1625, n_716, n_717);
  not g1257 (n_718, n1618);
  and g1258 (n1626, n_718, n1625);
  not g1259 (n_719, n1625);
  and g1260 (n1627, n1618, n_719);
  not g1261 (n_720, n1626);
  not g1262 (n_721, n1627);
  and g1263 (n1628, n_720, n_721);
  and g1264 (n1629, \A[670] , \A[671] );
  and g1265 (n1630, \A[672] , n_715);
  not g1266 (n_722, n1629);
  not g1267 (n_723, n1630);
  and g1268 (n1631, n_722, n_723);
  and g1269 (n1632, \A[667] , \A[668] );
  and g1270 (n1633, \A[669] , n_704);
  not g1271 (n_724, n1632);
  not g1272 (n_725, n1633);
  and g1273 (n1634, n_724, n_725);
  not g1274 (n_726, n1631);
  and g1275 (n1635, n_726, n1634);
  not g1276 (n_727, n1634);
  and g1277 (n1636, n1631, n_727);
  not g1278 (n_728, n1635);
  not g1279 (n_729, n1636);
  and g1280 (n1637, n_728, n_729);
  and g1281 (n1638, n_718, n_719);
  not g1282 (n_730, n1637);
  and g1283 (n1639, n_730, n1638);
  and g1284 (n1640, n_726, n_727);
  not g1285 (n_731, n1639);
  not g1286 (n_732, n1640);
  and g1287 (n1641, n_731, n_732);
  and g1288 (n1642, n_728, n1638);
  and g1289 (n1643, n_729, n1642);
  not g1290 (n_733, n1638);
  and g1291 (n1644, n_730, n_733);
  not g1292 (n_734, n1643);
  not g1293 (n_735, n1644);
  and g1294 (n1645, n_734, n_735);
  not g1295 (n_736, n1641);
  not g1296 (n_737, n1645);
  and g1297 (n1646, n_736, n_737);
  not g1298 (n_738, n1628);
  not g1299 (n_739, n1646);
  and g1300 (n1647, n_738, n_739);
  not g1301 (n_740, n1611);
  and g1302 (n1648, n_740, n1647);
  not g1303 (n_741, n1647);
  and g1304 (n1649, n1611, n_741);
  not g1305 (n_742, n1648);
  not g1306 (n_743, n1649);
  and g1307 (n1650, n_742, n_743);
  not g1308 (n_745, \A[661] );
  and g1309 (n1651, n_745, \A[662] );
  not g1310 (n_747, \A[662] );
  and g1311 (n1652, \A[661] , n_747);
  not g1312 (n_749, n1652);
  and g1313 (n1653, \A[663] , n_749);
  not g1314 (n_750, n1651);
  and g1315 (n1654, n_750, n1653);
  and g1316 (n1655, n_750, n_749);
  not g1317 (n_751, \A[663] );
  not g1318 (n_752, n1655);
  and g1319 (n1656, n_751, n_752);
  not g1320 (n_753, n1654);
  not g1321 (n_754, n1656);
  and g1322 (n1657, n_753, n_754);
  not g1323 (n_756, \A[664] );
  and g1324 (n1658, n_756, \A[665] );
  not g1325 (n_758, \A[665] );
  and g1326 (n1659, \A[664] , n_758);
  not g1327 (n_760, n1659);
  and g1328 (n1660, \A[666] , n_760);
  not g1329 (n_761, n1658);
  and g1330 (n1661, n_761, n1660);
  and g1331 (n1662, n_761, n_760);
  not g1332 (n_762, \A[666] );
  not g1333 (n_763, n1662);
  and g1334 (n1663, n_762, n_763);
  not g1335 (n_764, n1661);
  not g1336 (n_765, n1663);
  and g1337 (n1664, n_764, n_765);
  not g1338 (n_766, n1657);
  and g1339 (n1665, n_766, n1664);
  not g1340 (n_767, n1664);
  and g1341 (n1666, n1657, n_767);
  not g1342 (n_768, n1665);
  not g1343 (n_769, n1666);
  and g1344 (n1667, n_768, n_769);
  and g1345 (n1668, \A[664] , \A[665] );
  and g1346 (n1669, \A[666] , n_763);
  not g1347 (n_770, n1668);
  not g1348 (n_771, n1669);
  and g1349 (n1670, n_770, n_771);
  and g1350 (n1671, \A[661] , \A[662] );
  and g1351 (n1672, \A[663] , n_752);
  not g1352 (n_772, n1671);
  not g1353 (n_773, n1672);
  and g1354 (n1673, n_772, n_773);
  not g1355 (n_774, n1670);
  and g1356 (n1674, n_774, n1673);
  not g1357 (n_775, n1673);
  and g1358 (n1675, n1670, n_775);
  not g1359 (n_776, n1674);
  not g1360 (n_777, n1675);
  and g1361 (n1676, n_776, n_777);
  and g1362 (n1677, n_766, n_767);
  not g1363 (n_778, n1676);
  and g1364 (n1678, n_778, n1677);
  and g1365 (n1679, n_774, n_775);
  not g1366 (n_779, n1678);
  not g1367 (n_780, n1679);
  and g1368 (n1680, n_779, n_780);
  and g1369 (n1681, n_776, n1677);
  and g1370 (n1682, n_777, n1681);
  not g1371 (n_781, n1677);
  and g1372 (n1683, n_778, n_781);
  not g1373 (n_782, n1682);
  not g1374 (n_783, n1683);
  and g1375 (n1684, n_782, n_783);
  not g1376 (n_784, n1680);
  not g1377 (n_785, n1684);
  and g1378 (n1685, n_784, n_785);
  not g1379 (n_786, n1667);
  not g1380 (n_787, n1685);
  and g1381 (n1686, n_786, n_787);
  not g1382 (n_789, \A[655] );
  and g1383 (n1687, n_789, \A[656] );
  not g1384 (n_791, \A[656] );
  and g1385 (n1688, \A[655] , n_791);
  not g1386 (n_793, n1688);
  and g1387 (n1689, \A[657] , n_793);
  not g1388 (n_794, n1687);
  and g1389 (n1690, n_794, n1689);
  and g1390 (n1691, n_794, n_793);
  not g1391 (n_795, \A[657] );
  not g1392 (n_796, n1691);
  and g1393 (n1692, n_795, n_796);
  not g1394 (n_797, n1690);
  not g1395 (n_798, n1692);
  and g1396 (n1693, n_797, n_798);
  not g1397 (n_800, \A[658] );
  and g1398 (n1694, n_800, \A[659] );
  not g1399 (n_802, \A[659] );
  and g1400 (n1695, \A[658] , n_802);
  not g1401 (n_804, n1695);
  and g1402 (n1696, \A[660] , n_804);
  not g1403 (n_805, n1694);
  and g1404 (n1697, n_805, n1696);
  and g1405 (n1698, n_805, n_804);
  not g1406 (n_806, \A[660] );
  not g1407 (n_807, n1698);
  and g1408 (n1699, n_806, n_807);
  not g1409 (n_808, n1697);
  not g1410 (n_809, n1699);
  and g1411 (n1700, n_808, n_809);
  not g1412 (n_810, n1693);
  and g1413 (n1701, n_810, n1700);
  not g1414 (n_811, n1700);
  and g1415 (n1702, n1693, n_811);
  not g1416 (n_812, n1701);
  not g1417 (n_813, n1702);
  and g1418 (n1703, n_812, n_813);
  and g1419 (n1704, \A[658] , \A[659] );
  and g1420 (n1705, \A[660] , n_807);
  not g1421 (n_814, n1704);
  not g1422 (n_815, n1705);
  and g1423 (n1706, n_814, n_815);
  and g1424 (n1707, \A[655] , \A[656] );
  and g1425 (n1708, \A[657] , n_796);
  not g1426 (n_816, n1707);
  not g1427 (n_817, n1708);
  and g1428 (n1709, n_816, n_817);
  not g1429 (n_818, n1706);
  and g1430 (n1710, n_818, n1709);
  not g1431 (n_819, n1709);
  and g1432 (n1711, n1706, n_819);
  not g1433 (n_820, n1710);
  not g1434 (n_821, n1711);
  and g1435 (n1712, n_820, n_821);
  and g1436 (n1713, n_810, n_811);
  not g1437 (n_822, n1712);
  and g1438 (n1714, n_822, n1713);
  and g1439 (n1715, n_818, n_819);
  not g1440 (n_823, n1714);
  not g1441 (n_824, n1715);
  and g1442 (n1716, n_823, n_824);
  and g1443 (n1717, n_820, n1713);
  and g1444 (n1718, n_821, n1717);
  not g1445 (n_825, n1713);
  and g1446 (n1719, n_822, n_825);
  not g1447 (n_826, n1718);
  not g1448 (n_827, n1719);
  and g1449 (n1720, n_826, n_827);
  not g1450 (n_828, n1716);
  not g1451 (n_829, n1720);
  and g1452 (n1721, n_828, n_829);
  not g1453 (n_830, n1703);
  not g1454 (n_831, n1721);
  and g1455 (n1722, n_830, n_831);
  not g1456 (n_832, n1686);
  and g1457 (n1723, n_832, n1722);
  not g1458 (n_833, n1722);
  and g1459 (n1724, n1686, n_833);
  not g1460 (n_834, n1723);
  not g1461 (n_835, n1724);
  and g1462 (n1725, n_834, n_835);
  not g1463 (n_836, n1650);
  and g1464 (n1726, n_836, n1725);
  not g1465 (n_837, n1725);
  and g1466 (n1727, n1650, n_837);
  not g1467 (n_838, n1726);
  not g1468 (n_839, n1727);
  and g1469 (n1728, n_838, n_839);
  not g1470 (n_840, n1575);
  and g1471 (n1729, n_840, n1728);
  not g1472 (n_841, n1728);
  and g1473 (n1730, n1575, n_841);
  not g1474 (n_842, n1729);
  not g1475 (n_843, n1730);
  and g1476 (n1731, n_842, n_843);
  not g1477 (n_844, n1422);
  not g1478 (n_845, n1731);
  and g1479 (n1732, n_844, n_845);
  not g1480 (n_846, n1419);
  and g1481 (n1733, n_846, n1732);
  not g1482 (n_847, n1414);
  and g1483 (n1734, n_847, n1733);
  and g1484 (n1735, n_847, n_846);
  not g1485 (n_848, n1732);
  not g1486 (n_849, n1735);
  and g1487 (n1736, n_848, n_849);
  not g1488 (n_850, n1734);
  not g1489 (n_851, n1736);
  and g1490 (n1737, n_850, n_851);
  and g1491 (n1738, n_642, n_640);
  not g1492 (n_852, n1738);
  and g1493 (n1739, n_641, n_852);
  and g1494 (n1740, n_598, n_642);
  and g1495 (n1741, n_599, n1740);
  and g1496 (n1742, n_643, n1741);
  and g1497 (n1743, n_598, n_596);
  not g1498 (n_853, n1743);
  and g1499 (n1744, n_597, n_853);
  not g1500 (n_854, n1742);
  and g1501 (n1745, n_854, n1744);
  not g1502 (n_855, n1744);
  and g1503 (n1746, n1742, n_855);
  not g1504 (n_856, n1745);
  not g1505 (n_857, n1746);
  and g1506 (n1747, n_856, n_857);
  not g1507 (n_858, n1739);
  not g1508 (n_859, n1747);
  and g1509 (n1748, n_858, n_859);
  and g1510 (n1749, n_854, n_855);
  not g1515 (n_860, n1749);
  not g1516 (n_861, n1753);
  and g1517 (n1754, n_860, n_861);
  not g1518 (n_862, n1754);
  and g1519 (n1755, n1739, n_862);
  not g1520 (n_863, n1748);
  not g1521 (n_864, n1755);
  and g1522 (n1756, n_863, n_864);
  and g1523 (n1757, n_550, n_548);
  not g1524 (n_865, n1757);
  and g1525 (n1758, n_549, n_865);
  and g1526 (n1759, n_506, n_550);
  and g1527 (n1760, n_507, n1759);
  and g1528 (n1761, n_551, n1760);
  and g1529 (n1762, n_506, n_504);
  not g1530 (n_866, n1762);
  and g1531 (n1763, n_505, n_866);
  not g1532 (n_867, n1761);
  not g1533 (n_868, n1763);
  and g1534 (n1764, n_867, n_868);
  not g1539 (n_869, n1764);
  not g1540 (n_870, n1768);
  and g1541 (n1769, n_869, n_870);
  not g1542 (n_871, n1769);
  and g1543 (n1770, n1758, n_871);
  and g1544 (n1771, n_867, n1763);
  and g1545 (n1772, n1761, n_868);
  not g1546 (n_872, n1771);
  not g1547 (n_873, n1772);
  and g1548 (n1773, n_872, n_873);
  not g1549 (n_874, n1758);
  not g1550 (n_875, n1773);
  and g1551 (n1774, n_874, n_875);
  and g1552 (n1775, n_648, n_649);
  not g1553 (n_876, n1774);
  not g1554 (n_877, n1775);
  and g1555 (n1776, n_876, n_877);
  not g1556 (n_878, n1770);
  and g1557 (n1777, n_878, n1776);
  and g1558 (n1778, n_878, n_876);
  not g1559 (n_879, n1778);
  and g1560 (n1779, n1775, n_879);
  not g1561 (n_880, n1777);
  not g1562 (n_881, n1779);
  and g1563 (n1780, n_880, n_881);
  not g1564 (n_882, n1756);
  not g1565 (n_883, n1780);
  and g1566 (n1781, n_882, n_883);
  and g1567 (n1782, n_876, n1775);
  and g1568 (n1783, n_878, n1782);
  and g1569 (n1784, n_877, n_879);
  not g1570 (n_884, n1783);
  not g1571 (n_885, n1784);
  and g1572 (n1785, n_884, n_885);
  not g1573 (n_886, n1785);
  and g1574 (n1786, n1756, n_886);
  and g1575 (n1787, n_840, n_841);
  not g1576 (n_887, n1786);
  and g1577 (n1788, n_887, n1787);
  not g1578 (n_888, n1781);
  and g1579 (n1789, n_888, n1788);
  and g1580 (n1790, n_888, n_887);
  not g1581 (n_889, n1787);
  not g1582 (n_890, n1790);
  and g1583 (n1791, n_889, n_890);
  not g1584 (n_891, n1789);
  not g1585 (n_892, n1791);
  and g1586 (n1792, n_891, n_892);
  and g1587 (n1793, n_738, n_736);
  not g1588 (n_893, n1793);
  and g1589 (n1794, n_737, n_893);
  and g1590 (n1795, n_694, n_738);
  and g1591 (n1796, n_695, n1795);
  and g1592 (n1797, n_739, n1796);
  and g1593 (n1798, n_694, n_692);
  not g1594 (n_894, n1798);
  and g1595 (n1799, n_693, n_894);
  not g1596 (n_895, n1797);
  not g1597 (n_896, n1799);
  and g1598 (n1800, n_895, n_896);
  not g1603 (n_897, n1800);
  not g1604 (n_898, n1804);
  and g1605 (n1805, n_897, n_898);
  not g1606 (n_899, n1805);
  and g1607 (n1806, n1794, n_899);
  and g1608 (n1807, n_895, n1799);
  and g1609 (n1808, n1797, n_896);
  not g1610 (n_900, n1807);
  not g1611 (n_901, n1808);
  and g1612 (n1809, n_900, n_901);
  not g1613 (n_902, n1794);
  not g1614 (n_903, n1809);
  and g1615 (n1810, n_902, n_903);
  and g1616 (n1811, n_836, n_837);
  not g1617 (n_904, n1810);
  and g1618 (n1812, n_904, n1811);
  not g1619 (n_905, n1806);
  and g1620 (n1813, n_905, n1812);
  and g1621 (n1814, n_905, n_904);
  not g1622 (n_906, n1811);
  not g1623 (n_907, n1814);
  and g1624 (n1815, n_906, n_907);
  not g1625 (n_908, n1813);
  not g1626 (n_909, n1815);
  and g1627 (n1816, n_908, n_909);
  and g1628 (n1817, n_830, n_828);
  not g1629 (n_910, n1817);
  and g1630 (n1818, n_829, n_910);
  and g1631 (n1819, n_786, n_830);
  and g1632 (n1820, n_787, n1819);
  and g1633 (n1821, n_831, n1820);
  and g1634 (n1822, n_786, n_784);
  not g1635 (n_911, n1822);
  and g1636 (n1823, n_785, n_911);
  not g1637 (n_912, n1821);
  and g1638 (n1824, n_912, n1823);
  not g1639 (n_913, n1823);
  and g1640 (n1825, n1821, n_913);
  not g1641 (n_914, n1824);
  not g1642 (n_915, n1825);
  and g1643 (n1826, n_914, n_915);
  not g1644 (n_916, n1818);
  not g1645 (n_917, n1826);
  and g1646 (n1827, n_916, n_917);
  and g1647 (n1828, n_912, n_913);
  not g1652 (n_918, n1828);
  not g1653 (n_919, n1832);
  and g1654 (n1833, n_918, n_919);
  not g1655 (n_920, n1833);
  and g1656 (n1834, n1818, n_920);
  not g1657 (n_921, n1827);
  not g1658 (n_922, n1834);
  and g1659 (n1835, n_921, n_922);
  not g1660 (n_923, n1816);
  and g1661 (n1836, n_923, n1835);
  and g1662 (n1837, n_904, n_906);
  and g1663 (n1838, n_905, n1837);
  and g1664 (n1839, n1811, n_907);
  not g1665 (n_924, n1838);
  not g1666 (n_925, n1839);
  and g1667 (n1840, n_924, n_925);
  not g1668 (n_926, n1835);
  not g1669 (n_927, n1840);
  and g1670 (n1841, n_926, n_927);
  not g1671 (n_928, n1836);
  not g1672 (n_929, n1841);
  and g1673 (n1842, n_928, n_929);
  not g1674 (n_930, n1792);
  and g1675 (n1843, n_930, n1842);
  and g1676 (n1844, n_887, n_889);
  and g1677 (n1845, n_888, n1844);
  and g1678 (n1846, n1787, n_890);
  not g1679 (n_931, n1845);
  not g1680 (n_932, n1846);
  and g1681 (n1847, n_931, n_932);
  not g1682 (n_933, n1842);
  not g1683 (n_934, n1847);
  and g1684 (n1848, n_933, n_934);
  not g1685 (n_935, n1843);
  not g1686 (n_936, n1848);
  and g1687 (n1849, n_935, n_936);
  not g1688 (n_937, n1737);
  and g1689 (n1850, n_937, n1849);
  and g1690 (n1851, n_846, n_848);
  and g1691 (n1852, n_847, n1851);
  and g1692 (n1853, n1732, n_849);
  not g1693 (n_938, n1852);
  not g1694 (n_939, n1853);
  and g1695 (n1854, n_938, n_939);
  not g1696 (n_940, n1849);
  not g1697 (n_941, n1854);
  and g1698 (n1855, n_940, n_941);
  not g1699 (n_942, n1850);
  not g1700 (n_943, n1855);
  and g1701 (n1856, n_942, n_943);
  and g1702 (n1857, \A[778] , \A[779] );
  not g1703 (n_946, \A[779] );
  and g1704 (n1858, \A[778] , n_946);
  not g1705 (n_947, \A[778] );
  and g1706 (n1859, n_947, \A[779] );
  not g1707 (n_948, n1858);
  not g1708 (n_949, n1859);
  and g1709 (n1860, n_948, n_949);
  not g1710 (n_951, n1860);
  and g1711 (n1861, \A[780] , n_951);
  not g1712 (n_952, n1857);
  not g1713 (n_953, n1861);
  and g1714 (n1862, n_952, n_953);
  and g1715 (n1863, \A[775] , \A[776] );
  not g1716 (n_956, \A[776] );
  and g1717 (n1864, \A[775] , n_956);
  not g1718 (n_957, \A[775] );
  and g1719 (n1865, n_957, \A[776] );
  not g1720 (n_958, n1864);
  not g1721 (n_959, n1865);
  and g1722 (n1866, n_958, n_959);
  not g1723 (n_961, n1866);
  and g1724 (n1867, \A[777] , n_961);
  not g1725 (n_962, n1863);
  not g1726 (n_963, n1867);
  and g1727 (n1868, n_962, n_963);
  not g1728 (n_964, n1868);
  and g1729 (n1869, n1862, n_964);
  not g1730 (n_965, n1862);
  and g1731 (n1870, n_965, n1868);
  and g1732 (n1871, \A[777] , n_958);
  and g1733 (n1872, n_959, n1871);
  not g1734 (n_966, \A[777] );
  and g1735 (n1873, n_966, n_961);
  not g1736 (n_967, n1872);
  not g1737 (n_968, n1873);
  and g1738 (n1874, n_967, n_968);
  and g1739 (n1875, \A[780] , n_948);
  and g1740 (n1876, n_949, n1875);
  not g1741 (n_969, \A[780] );
  and g1742 (n1877, n_969, n_951);
  not g1743 (n_970, n1876);
  not g1744 (n_971, n1877);
  and g1745 (n1878, n_970, n_971);
  not g1746 (n_972, n1874);
  not g1747 (n_973, n1878);
  and g1748 (n1879, n_972, n_973);
  not g1749 (n_974, n1870);
  and g1750 (n1880, n_974, n1879);
  not g1751 (n_975, n1869);
  and g1752 (n1881, n_975, n1880);
  and g1753 (n1882, n_975, n_974);
  not g1754 (n_976, n1879);
  not g1755 (n_977, n1882);
  and g1756 (n1883, n_976, n_977);
  not g1757 (n_978, n1881);
  not g1758 (n_979, n1883);
  and g1759 (n1884, n_978, n_979);
  and g1760 (n1885, n_972, n1878);
  and g1761 (n1886, n1874, n_973);
  not g1762 (n_980, n1885);
  not g1763 (n_981, n1886);
  and g1764 (n1887, n_980, n_981);
  and g1765 (n1888, n1879, n_977);
  and g1766 (n1889, n_965, n_964);
  not g1767 (n_982, n1888);
  not g1768 (n_983, n1889);
  and g1769 (n1890, n_982, n_983);
  not g1770 (n_984, n1887);
  not g1771 (n_985, n1890);
  and g1772 (n1891, n_984, n_985);
  not g1773 (n_986, n1884);
  not g1774 (n_987, n1891);
  and g1775 (n1892, n_986, n_987);
  and g1776 (n1893, n_986, n_985);
  and g1777 (n1894, \A[784] , \A[785] );
  not g1778 (n_990, \A[785] );
  and g1779 (n1895, \A[784] , n_990);
  not g1780 (n_991, \A[784] );
  and g1781 (n1896, n_991, \A[785] );
  not g1782 (n_992, n1895);
  not g1783 (n_993, n1896);
  and g1784 (n1897, n_992, n_993);
  not g1785 (n_995, n1897);
  and g1786 (n1898, \A[786] , n_995);
  not g1787 (n_996, n1894);
  not g1788 (n_997, n1898);
  and g1789 (n1899, n_996, n_997);
  and g1790 (n1900, \A[781] , \A[782] );
  not g1791 (n_1000, \A[782] );
  and g1792 (n1901, \A[781] , n_1000);
  not g1793 (n_1001, \A[781] );
  and g1794 (n1902, n_1001, \A[782] );
  not g1795 (n_1002, n1901);
  not g1796 (n_1003, n1902);
  and g1797 (n1903, n_1002, n_1003);
  not g1798 (n_1005, n1903);
  and g1799 (n1904, \A[783] , n_1005);
  not g1800 (n_1006, n1900);
  not g1801 (n_1007, n1904);
  and g1802 (n1905, n_1006, n_1007);
  not g1803 (n_1008, n1899);
  and g1804 (n1906, n_1008, n1905);
  not g1805 (n_1009, n1905);
  and g1806 (n1907, n1899, n_1009);
  not g1807 (n_1010, n1906);
  not g1808 (n_1011, n1907);
  and g1809 (n1908, n_1010, n_1011);
  and g1810 (n1909, \A[783] , n_1002);
  and g1811 (n1910, n_1003, n1909);
  not g1812 (n_1012, \A[783] );
  and g1813 (n1911, n_1012, n_1005);
  not g1814 (n_1013, n1910);
  not g1815 (n_1014, n1911);
  and g1816 (n1912, n_1013, n_1014);
  and g1817 (n1913, \A[786] , n_992);
  and g1818 (n1914, n_993, n1913);
  not g1819 (n_1015, \A[786] );
  and g1820 (n1915, n_1015, n_995);
  not g1821 (n_1016, n1914);
  not g1822 (n_1017, n1915);
  and g1823 (n1916, n_1016, n_1017);
  not g1824 (n_1018, n1912);
  not g1825 (n_1019, n1916);
  and g1826 (n1917, n_1018, n_1019);
  not g1827 (n_1020, n1908);
  and g1828 (n1918, n_1020, n1917);
  and g1829 (n1919, n_1008, n_1009);
  not g1830 (n_1021, n1918);
  not g1831 (n_1022, n1919);
  and g1832 (n1920, n_1021, n_1022);
  and g1833 (n1921, n_1010, n1917);
  and g1834 (n1922, n_1011, n1921);
  not g1835 (n_1023, n1917);
  and g1836 (n1923, n_1020, n_1023);
  not g1837 (n_1024, n1922);
  not g1838 (n_1025, n1923);
  and g1839 (n1924, n_1024, n_1025);
  not g1840 (n_1026, n1920);
  not g1841 (n_1027, n1924);
  and g1842 (n1925, n_1026, n_1027);
  and g1843 (n1926, n_1018, n1916);
  and g1844 (n1927, n1912, n_1019);
  not g1845 (n_1028, n1926);
  not g1846 (n_1029, n1927);
  and g1847 (n1928, n_1028, n_1029);
  not g1848 (n_1030, n1928);
  and g1849 (n1929, n_984, n_1030);
  not g1850 (n_1031, n1925);
  and g1851 (n1930, n_1031, n1929);
  not g1852 (n_1032, n1893);
  and g1853 (n1931, n_1032, n1930);
  and g1854 (n1932, n_1026, n_1030);
  not g1855 (n_1033, n1932);
  and g1856 (n1933, n_1027, n_1033);
  not g1857 (n_1034, n1931);
  and g1858 (n1934, n_1034, n1933);
  not g1859 (n_1035, n1933);
  and g1860 (n1935, n1931, n_1035);
  not g1861 (n_1036, n1934);
  not g1862 (n_1037, n1935);
  and g1863 (n1936, n_1036, n_1037);
  not g1864 (n_1038, n1892);
  not g1865 (n_1039, n1936);
  and g1866 (n1937, n_1038, n_1039);
  and g1867 (n1938, n_1034, n_1035);
  not g1872 (n_1040, n1938);
  not g1873 (n_1041, n1942);
  and g1874 (n1943, n_1040, n_1041);
  not g1875 (n_1042, n1943);
  and g1876 (n1944, n1892, n_1042);
  not g1877 (n_1043, n1937);
  not g1878 (n_1044, n1944);
  and g1879 (n1945, n_1043, n_1044);
  and g1880 (n1946, \A[790] , \A[791] );
  not g1881 (n_1047, \A[791] );
  and g1882 (n1947, \A[790] , n_1047);
  not g1883 (n_1048, \A[790] );
  and g1884 (n1948, n_1048, \A[791] );
  not g1885 (n_1049, n1947);
  not g1886 (n_1050, n1948);
  and g1887 (n1949, n_1049, n_1050);
  not g1888 (n_1052, n1949);
  and g1889 (n1950, \A[792] , n_1052);
  not g1890 (n_1053, n1946);
  not g1891 (n_1054, n1950);
  and g1892 (n1951, n_1053, n_1054);
  and g1893 (n1952, \A[787] , \A[788] );
  not g1894 (n_1057, \A[788] );
  and g1895 (n1953, \A[787] , n_1057);
  not g1896 (n_1058, \A[787] );
  and g1897 (n1954, n_1058, \A[788] );
  not g1898 (n_1059, n1953);
  not g1899 (n_1060, n1954);
  and g1900 (n1955, n_1059, n_1060);
  not g1901 (n_1062, n1955);
  and g1902 (n1956, \A[789] , n_1062);
  not g1903 (n_1063, n1952);
  not g1904 (n_1064, n1956);
  and g1905 (n1957, n_1063, n_1064);
  not g1906 (n_1065, n1957);
  and g1907 (n1958, n1951, n_1065);
  not g1908 (n_1066, n1951);
  and g1909 (n1959, n_1066, n1957);
  and g1910 (n1960, \A[789] , n_1059);
  and g1911 (n1961, n_1060, n1960);
  not g1912 (n_1067, \A[789] );
  and g1913 (n1962, n_1067, n_1062);
  not g1914 (n_1068, n1961);
  not g1915 (n_1069, n1962);
  and g1916 (n1963, n_1068, n_1069);
  and g1917 (n1964, \A[792] , n_1049);
  and g1918 (n1965, n_1050, n1964);
  not g1919 (n_1070, \A[792] );
  and g1920 (n1966, n_1070, n_1052);
  not g1921 (n_1071, n1965);
  not g1922 (n_1072, n1966);
  and g1923 (n1967, n_1071, n_1072);
  not g1924 (n_1073, n1963);
  not g1925 (n_1074, n1967);
  and g1926 (n1968, n_1073, n_1074);
  not g1927 (n_1075, n1959);
  and g1928 (n1969, n_1075, n1968);
  not g1929 (n_1076, n1958);
  and g1930 (n1970, n_1076, n1969);
  and g1931 (n1971, n_1076, n_1075);
  not g1932 (n_1077, n1968);
  not g1933 (n_1078, n1971);
  and g1934 (n1972, n_1077, n_1078);
  not g1935 (n_1079, n1970);
  not g1936 (n_1080, n1972);
  and g1937 (n1973, n_1079, n_1080);
  and g1938 (n1974, n_1073, n1967);
  and g1939 (n1975, n1963, n_1074);
  not g1940 (n_1081, n1974);
  not g1941 (n_1082, n1975);
  and g1942 (n1976, n_1081, n_1082);
  and g1943 (n1977, n1968, n_1078);
  and g1944 (n1978, n_1066, n_1065);
  not g1945 (n_1083, n1977);
  not g1946 (n_1084, n1978);
  and g1947 (n1979, n_1083, n_1084);
  not g1948 (n_1085, n1976);
  not g1949 (n_1086, n1979);
  and g1950 (n1980, n_1085, n_1086);
  not g1951 (n_1087, n1973);
  not g1952 (n_1088, n1980);
  and g1953 (n1981, n_1087, n_1088);
  and g1954 (n1982, n_1087, n_1086);
  and g1955 (n1983, \A[796] , \A[797] );
  not g1956 (n_1091, \A[797] );
  and g1957 (n1984, \A[796] , n_1091);
  not g1958 (n_1092, \A[796] );
  and g1959 (n1985, n_1092, \A[797] );
  not g1960 (n_1093, n1984);
  not g1961 (n_1094, n1985);
  and g1962 (n1986, n_1093, n_1094);
  not g1963 (n_1096, n1986);
  and g1964 (n1987, \A[798] , n_1096);
  not g1965 (n_1097, n1983);
  not g1966 (n_1098, n1987);
  and g1967 (n1988, n_1097, n_1098);
  and g1968 (n1989, \A[793] , \A[794] );
  not g1969 (n_1101, \A[794] );
  and g1970 (n1990, \A[793] , n_1101);
  not g1971 (n_1102, \A[793] );
  and g1972 (n1991, n_1102, \A[794] );
  not g1973 (n_1103, n1990);
  not g1974 (n_1104, n1991);
  and g1975 (n1992, n_1103, n_1104);
  not g1976 (n_1106, n1992);
  and g1977 (n1993, \A[795] , n_1106);
  not g1978 (n_1107, n1989);
  not g1979 (n_1108, n1993);
  and g1980 (n1994, n_1107, n_1108);
  not g1981 (n_1109, n1988);
  and g1982 (n1995, n_1109, n1994);
  not g1983 (n_1110, n1994);
  and g1984 (n1996, n1988, n_1110);
  not g1985 (n_1111, n1995);
  not g1986 (n_1112, n1996);
  and g1987 (n1997, n_1111, n_1112);
  and g1988 (n1998, \A[795] , n_1103);
  and g1989 (n1999, n_1104, n1998);
  not g1990 (n_1113, \A[795] );
  and g1991 (n2000, n_1113, n_1106);
  not g1992 (n_1114, n1999);
  not g1993 (n_1115, n2000);
  and g1994 (n2001, n_1114, n_1115);
  and g1995 (n2002, \A[798] , n_1093);
  and g1996 (n2003, n_1094, n2002);
  not g1997 (n_1116, \A[798] );
  and g1998 (n2004, n_1116, n_1096);
  not g1999 (n_1117, n2003);
  not g2000 (n_1118, n2004);
  and g2001 (n2005, n_1117, n_1118);
  not g2002 (n_1119, n2001);
  not g2003 (n_1120, n2005);
  and g2004 (n2006, n_1119, n_1120);
  not g2005 (n_1121, n1997);
  and g2006 (n2007, n_1121, n2006);
  and g2007 (n2008, n_1109, n_1110);
  not g2008 (n_1122, n2007);
  not g2009 (n_1123, n2008);
  and g2010 (n2009, n_1122, n_1123);
  and g2011 (n2010, n_1111, n2006);
  and g2012 (n2011, n_1112, n2010);
  not g2013 (n_1124, n2006);
  and g2014 (n2012, n_1121, n_1124);
  not g2015 (n_1125, n2011);
  not g2016 (n_1126, n2012);
  and g2017 (n2013, n_1125, n_1126);
  not g2018 (n_1127, n2009);
  not g2019 (n_1128, n2013);
  and g2020 (n2014, n_1127, n_1128);
  and g2021 (n2015, n_1119, n2005);
  and g2022 (n2016, n2001, n_1120);
  not g2023 (n_1129, n2015);
  not g2024 (n_1130, n2016);
  and g2025 (n2017, n_1129, n_1130);
  not g2026 (n_1131, n2017);
  and g2027 (n2018, n_1085, n_1131);
  not g2028 (n_1132, n2014);
  and g2029 (n2019, n_1132, n2018);
  not g2030 (n_1133, n1982);
  and g2031 (n2020, n_1133, n2019);
  and g2032 (n2021, n_1127, n_1131);
  not g2033 (n_1134, n2021);
  and g2034 (n2022, n_1128, n_1134);
  not g2035 (n_1135, n2020);
  not g2036 (n_1136, n2022);
  and g2037 (n2023, n_1135, n_1136);
  not g2042 (n_1137, n2023);
  not g2043 (n_1138, n2027);
  and g2044 (n2028, n_1137, n_1138);
  not g2045 (n_1139, n2028);
  and g2046 (n2029, n1981, n_1139);
  and g2047 (n2030, n_1135, n2022);
  and g2048 (n2031, n2020, n_1136);
  not g2049 (n_1140, n2030);
  not g2050 (n_1141, n2031);
  and g2051 (n2032, n_1140, n_1141);
  not g2052 (n_1142, n1981);
  not g2053 (n_1143, n2032);
  and g2054 (n2033, n_1142, n_1143);
  and g2055 (n2034, n_1132, n_1131);
  and g2056 (n2035, n_1085, n_1133);
  not g2057 (n_1144, n2034);
  and g2058 (n2036, n_1144, n2035);
  not g2059 (n_1145, n2035);
  and g2060 (n2037, n2034, n_1145);
  not g2061 (n_1146, n2036);
  not g2062 (n_1147, n2037);
  and g2063 (n2038, n_1146, n_1147);
  and g2064 (n2039, n_1031, n_1030);
  and g2065 (n2040, n_984, n_1032);
  not g2066 (n_1148, n2039);
  and g2067 (n2041, n_1148, n2040);
  not g2068 (n_1149, n2040);
  and g2069 (n2042, n2039, n_1149);
  not g2070 (n_1150, n2041);
  not g2071 (n_1151, n2042);
  and g2072 (n2043, n_1150, n_1151);
  not g2073 (n_1152, n2038);
  not g2074 (n_1153, n2043);
  and g2075 (n2044, n_1152, n_1153);
  not g2076 (n_1154, n2033);
  not g2077 (n_1155, n2044);
  and g2078 (n2045, n_1154, n_1155);
  not g2079 (n_1156, n2029);
  and g2080 (n2046, n_1156, n2045);
  and g2081 (n2047, n_1156, n_1154);
  not g2082 (n_1157, n2047);
  and g2083 (n2048, n2044, n_1157);
  not g2084 (n_1158, n2046);
  not g2085 (n_1159, n2048);
  and g2086 (n2049, n_1158, n_1159);
  not g2087 (n_1160, n1945);
  not g2088 (n_1161, n2049);
  and g2089 (n2050, n_1160, n_1161);
  and g2090 (n2051, n_1154, n2044);
  and g2091 (n2052, n_1156, n2051);
  and g2092 (n2053, n_1155, n_1157);
  not g2093 (n_1162, n2052);
  not g2094 (n_1163, n2053);
  and g2095 (n2054, n_1162, n_1163);
  not g2096 (n_1164, n2054);
  and g2097 (n2055, n1945, n_1164);
  and g2098 (n2056, n_1152, n2043);
  and g2099 (n2057, n2038, n_1153);
  not g2100 (n_1165, n2056);
  not g2101 (n_1166, n2057);
  and g2102 (n2058, n_1165, n_1166);
  not g2103 (n_1168, \A[769] );
  and g2104 (n2059, n_1168, \A[770] );
  not g2105 (n_1170, \A[770] );
  and g2106 (n2060, \A[769] , n_1170);
  not g2107 (n_1172, n2060);
  and g2108 (n2061, \A[771] , n_1172);
  not g2109 (n_1173, n2059);
  and g2110 (n2062, n_1173, n2061);
  and g2111 (n2063, n_1173, n_1172);
  not g2112 (n_1174, \A[771] );
  not g2113 (n_1175, n2063);
  and g2114 (n2064, n_1174, n_1175);
  not g2115 (n_1176, n2062);
  not g2116 (n_1177, n2064);
  and g2117 (n2065, n_1176, n_1177);
  not g2118 (n_1179, \A[772] );
  and g2119 (n2066, n_1179, \A[773] );
  not g2120 (n_1181, \A[773] );
  and g2121 (n2067, \A[772] , n_1181);
  not g2122 (n_1183, n2067);
  and g2123 (n2068, \A[774] , n_1183);
  not g2124 (n_1184, n2066);
  and g2125 (n2069, n_1184, n2068);
  and g2126 (n2070, n_1184, n_1183);
  not g2127 (n_1185, \A[774] );
  not g2128 (n_1186, n2070);
  and g2129 (n2071, n_1185, n_1186);
  not g2130 (n_1187, n2069);
  not g2131 (n_1188, n2071);
  and g2132 (n2072, n_1187, n_1188);
  not g2133 (n_1189, n2065);
  and g2134 (n2073, n_1189, n2072);
  not g2135 (n_1190, n2072);
  and g2136 (n2074, n2065, n_1190);
  not g2137 (n_1191, n2073);
  not g2138 (n_1192, n2074);
  and g2139 (n2075, n_1191, n_1192);
  and g2140 (n2076, \A[772] , \A[773] );
  and g2141 (n2077, \A[774] , n_1186);
  not g2142 (n_1193, n2076);
  not g2143 (n_1194, n2077);
  and g2144 (n2078, n_1193, n_1194);
  and g2145 (n2079, \A[769] , \A[770] );
  and g2146 (n2080, \A[771] , n_1175);
  not g2147 (n_1195, n2079);
  not g2148 (n_1196, n2080);
  and g2149 (n2081, n_1195, n_1196);
  not g2150 (n_1197, n2078);
  and g2151 (n2082, n_1197, n2081);
  not g2152 (n_1198, n2081);
  and g2153 (n2083, n2078, n_1198);
  not g2154 (n_1199, n2082);
  not g2155 (n_1200, n2083);
  and g2156 (n2084, n_1199, n_1200);
  and g2157 (n2085, n_1189, n_1190);
  not g2158 (n_1201, n2084);
  and g2159 (n2086, n_1201, n2085);
  and g2160 (n2087, n_1197, n_1198);
  not g2161 (n_1202, n2086);
  not g2162 (n_1203, n2087);
  and g2163 (n2088, n_1202, n_1203);
  and g2164 (n2089, n_1199, n2085);
  and g2165 (n2090, n_1200, n2089);
  not g2166 (n_1204, n2085);
  and g2167 (n2091, n_1201, n_1204);
  not g2168 (n_1205, n2090);
  not g2169 (n_1206, n2091);
  and g2170 (n2092, n_1205, n_1206);
  not g2171 (n_1207, n2088);
  not g2172 (n_1208, n2092);
  and g2173 (n2093, n_1207, n_1208);
  not g2174 (n_1209, n2075);
  not g2175 (n_1210, n2093);
  and g2176 (n2094, n_1209, n_1210);
  not g2177 (n_1212, \A[763] );
  and g2178 (n2095, n_1212, \A[764] );
  not g2179 (n_1214, \A[764] );
  and g2180 (n2096, \A[763] , n_1214);
  not g2181 (n_1216, n2096);
  and g2182 (n2097, \A[765] , n_1216);
  not g2183 (n_1217, n2095);
  and g2184 (n2098, n_1217, n2097);
  and g2185 (n2099, n_1217, n_1216);
  not g2186 (n_1218, \A[765] );
  not g2187 (n_1219, n2099);
  and g2188 (n2100, n_1218, n_1219);
  not g2189 (n_1220, n2098);
  not g2190 (n_1221, n2100);
  and g2191 (n2101, n_1220, n_1221);
  not g2192 (n_1223, \A[766] );
  and g2193 (n2102, n_1223, \A[767] );
  not g2194 (n_1225, \A[767] );
  and g2195 (n2103, \A[766] , n_1225);
  not g2196 (n_1227, n2103);
  and g2197 (n2104, \A[768] , n_1227);
  not g2198 (n_1228, n2102);
  and g2199 (n2105, n_1228, n2104);
  and g2200 (n2106, n_1228, n_1227);
  not g2201 (n_1229, \A[768] );
  not g2202 (n_1230, n2106);
  and g2203 (n2107, n_1229, n_1230);
  not g2204 (n_1231, n2105);
  not g2205 (n_1232, n2107);
  and g2206 (n2108, n_1231, n_1232);
  not g2207 (n_1233, n2101);
  and g2208 (n2109, n_1233, n2108);
  not g2209 (n_1234, n2108);
  and g2210 (n2110, n2101, n_1234);
  not g2211 (n_1235, n2109);
  not g2212 (n_1236, n2110);
  and g2213 (n2111, n_1235, n_1236);
  and g2214 (n2112, \A[766] , \A[767] );
  and g2215 (n2113, \A[768] , n_1230);
  not g2216 (n_1237, n2112);
  not g2217 (n_1238, n2113);
  and g2218 (n2114, n_1237, n_1238);
  and g2219 (n2115, \A[763] , \A[764] );
  and g2220 (n2116, \A[765] , n_1219);
  not g2221 (n_1239, n2115);
  not g2222 (n_1240, n2116);
  and g2223 (n2117, n_1239, n_1240);
  not g2224 (n_1241, n2114);
  and g2225 (n2118, n_1241, n2117);
  not g2226 (n_1242, n2117);
  and g2227 (n2119, n2114, n_1242);
  not g2228 (n_1243, n2118);
  not g2229 (n_1244, n2119);
  and g2230 (n2120, n_1243, n_1244);
  and g2231 (n2121, n_1233, n_1234);
  not g2232 (n_1245, n2120);
  and g2233 (n2122, n_1245, n2121);
  and g2234 (n2123, n_1241, n_1242);
  not g2235 (n_1246, n2122);
  not g2236 (n_1247, n2123);
  and g2237 (n2124, n_1246, n_1247);
  and g2238 (n2125, n_1243, n2121);
  and g2239 (n2126, n_1244, n2125);
  not g2240 (n_1248, n2121);
  and g2241 (n2127, n_1245, n_1248);
  not g2242 (n_1249, n2126);
  not g2243 (n_1250, n2127);
  and g2244 (n2128, n_1249, n_1250);
  not g2245 (n_1251, n2124);
  not g2246 (n_1252, n2128);
  and g2247 (n2129, n_1251, n_1252);
  not g2248 (n_1253, n2111);
  not g2249 (n_1254, n2129);
  and g2250 (n2130, n_1253, n_1254);
  not g2251 (n_1255, n2094);
  and g2252 (n2131, n_1255, n2130);
  not g2253 (n_1256, n2130);
  and g2254 (n2132, n2094, n_1256);
  not g2255 (n_1257, n2131);
  not g2256 (n_1258, n2132);
  and g2257 (n2133, n_1257, n_1258);
  not g2258 (n_1260, \A[757] );
  and g2259 (n2134, n_1260, \A[758] );
  not g2260 (n_1262, \A[758] );
  and g2261 (n2135, \A[757] , n_1262);
  not g2262 (n_1264, n2135);
  and g2263 (n2136, \A[759] , n_1264);
  not g2264 (n_1265, n2134);
  and g2265 (n2137, n_1265, n2136);
  and g2266 (n2138, n_1265, n_1264);
  not g2267 (n_1266, \A[759] );
  not g2268 (n_1267, n2138);
  and g2269 (n2139, n_1266, n_1267);
  not g2270 (n_1268, n2137);
  not g2271 (n_1269, n2139);
  and g2272 (n2140, n_1268, n_1269);
  not g2273 (n_1271, \A[760] );
  and g2274 (n2141, n_1271, \A[761] );
  not g2275 (n_1273, \A[761] );
  and g2276 (n2142, \A[760] , n_1273);
  not g2277 (n_1275, n2142);
  and g2278 (n2143, \A[762] , n_1275);
  not g2279 (n_1276, n2141);
  and g2280 (n2144, n_1276, n2143);
  and g2281 (n2145, n_1276, n_1275);
  not g2282 (n_1277, \A[762] );
  not g2283 (n_1278, n2145);
  and g2284 (n2146, n_1277, n_1278);
  not g2285 (n_1279, n2144);
  not g2286 (n_1280, n2146);
  and g2287 (n2147, n_1279, n_1280);
  not g2288 (n_1281, n2140);
  and g2289 (n2148, n_1281, n2147);
  not g2290 (n_1282, n2147);
  and g2291 (n2149, n2140, n_1282);
  not g2292 (n_1283, n2148);
  not g2293 (n_1284, n2149);
  and g2294 (n2150, n_1283, n_1284);
  and g2295 (n2151, \A[760] , \A[761] );
  and g2296 (n2152, \A[762] , n_1278);
  not g2297 (n_1285, n2151);
  not g2298 (n_1286, n2152);
  and g2299 (n2153, n_1285, n_1286);
  and g2300 (n2154, \A[757] , \A[758] );
  and g2301 (n2155, \A[759] , n_1267);
  not g2302 (n_1287, n2154);
  not g2303 (n_1288, n2155);
  and g2304 (n2156, n_1287, n_1288);
  not g2305 (n_1289, n2153);
  and g2306 (n2157, n_1289, n2156);
  not g2307 (n_1290, n2156);
  and g2308 (n2158, n2153, n_1290);
  not g2309 (n_1291, n2157);
  not g2310 (n_1292, n2158);
  and g2311 (n2159, n_1291, n_1292);
  and g2312 (n2160, n_1281, n_1282);
  not g2313 (n_1293, n2159);
  and g2314 (n2161, n_1293, n2160);
  and g2315 (n2162, n_1289, n_1290);
  not g2316 (n_1294, n2161);
  not g2317 (n_1295, n2162);
  and g2318 (n2163, n_1294, n_1295);
  and g2319 (n2164, n_1291, n2160);
  and g2320 (n2165, n_1292, n2164);
  not g2321 (n_1296, n2160);
  and g2322 (n2166, n_1293, n_1296);
  not g2323 (n_1297, n2165);
  not g2324 (n_1298, n2166);
  and g2325 (n2167, n_1297, n_1298);
  not g2326 (n_1299, n2163);
  not g2327 (n_1300, n2167);
  and g2328 (n2168, n_1299, n_1300);
  not g2329 (n_1301, n2150);
  not g2330 (n_1302, n2168);
  and g2331 (n2169, n_1301, n_1302);
  not g2332 (n_1304, \A[751] );
  and g2333 (n2170, n_1304, \A[752] );
  not g2334 (n_1306, \A[752] );
  and g2335 (n2171, \A[751] , n_1306);
  not g2336 (n_1308, n2171);
  and g2337 (n2172, \A[753] , n_1308);
  not g2338 (n_1309, n2170);
  and g2339 (n2173, n_1309, n2172);
  and g2340 (n2174, n_1309, n_1308);
  not g2341 (n_1310, \A[753] );
  not g2342 (n_1311, n2174);
  and g2343 (n2175, n_1310, n_1311);
  not g2344 (n_1312, n2173);
  not g2345 (n_1313, n2175);
  and g2346 (n2176, n_1312, n_1313);
  not g2347 (n_1315, \A[754] );
  and g2348 (n2177, n_1315, \A[755] );
  not g2349 (n_1317, \A[755] );
  and g2350 (n2178, \A[754] , n_1317);
  not g2351 (n_1319, n2178);
  and g2352 (n2179, \A[756] , n_1319);
  not g2353 (n_1320, n2177);
  and g2354 (n2180, n_1320, n2179);
  and g2355 (n2181, n_1320, n_1319);
  not g2356 (n_1321, \A[756] );
  not g2357 (n_1322, n2181);
  and g2358 (n2182, n_1321, n_1322);
  not g2359 (n_1323, n2180);
  not g2360 (n_1324, n2182);
  and g2361 (n2183, n_1323, n_1324);
  not g2362 (n_1325, n2176);
  and g2363 (n2184, n_1325, n2183);
  not g2364 (n_1326, n2183);
  and g2365 (n2185, n2176, n_1326);
  not g2366 (n_1327, n2184);
  not g2367 (n_1328, n2185);
  and g2368 (n2186, n_1327, n_1328);
  and g2369 (n2187, \A[754] , \A[755] );
  and g2370 (n2188, \A[756] , n_1322);
  not g2371 (n_1329, n2187);
  not g2372 (n_1330, n2188);
  and g2373 (n2189, n_1329, n_1330);
  and g2374 (n2190, \A[751] , \A[752] );
  and g2375 (n2191, \A[753] , n_1311);
  not g2376 (n_1331, n2190);
  not g2377 (n_1332, n2191);
  and g2378 (n2192, n_1331, n_1332);
  not g2379 (n_1333, n2189);
  and g2380 (n2193, n_1333, n2192);
  not g2381 (n_1334, n2192);
  and g2382 (n2194, n2189, n_1334);
  not g2383 (n_1335, n2193);
  not g2384 (n_1336, n2194);
  and g2385 (n2195, n_1335, n_1336);
  and g2386 (n2196, n_1325, n_1326);
  not g2387 (n_1337, n2195);
  and g2388 (n2197, n_1337, n2196);
  and g2389 (n2198, n_1333, n_1334);
  not g2390 (n_1338, n2197);
  not g2391 (n_1339, n2198);
  and g2392 (n2199, n_1338, n_1339);
  and g2393 (n2200, n_1335, n2196);
  and g2394 (n2201, n_1336, n2200);
  not g2395 (n_1340, n2196);
  and g2396 (n2202, n_1337, n_1340);
  not g2397 (n_1341, n2201);
  not g2398 (n_1342, n2202);
  and g2399 (n2203, n_1341, n_1342);
  not g2400 (n_1343, n2199);
  not g2401 (n_1344, n2203);
  and g2402 (n2204, n_1343, n_1344);
  not g2403 (n_1345, n2186);
  not g2404 (n_1346, n2204);
  and g2405 (n2205, n_1345, n_1346);
  not g2406 (n_1347, n2169);
  and g2407 (n2206, n_1347, n2205);
  not g2408 (n_1348, n2205);
  and g2409 (n2207, n2169, n_1348);
  not g2410 (n_1349, n2206);
  not g2411 (n_1350, n2207);
  and g2412 (n2208, n_1349, n_1350);
  not g2413 (n_1351, n2133);
  and g2414 (n2209, n_1351, n2208);
  not g2415 (n_1352, n2208);
  and g2416 (n2210, n2133, n_1352);
  not g2417 (n_1353, n2209);
  not g2418 (n_1354, n2210);
  and g2419 (n2211, n_1353, n_1354);
  not g2420 (n_1355, n2058);
  not g2421 (n_1356, n2211);
  and g2422 (n2212, n_1355, n_1356);
  not g2423 (n_1357, n2055);
  and g2424 (n2213, n_1357, n2212);
  not g2425 (n_1358, n2050);
  and g2426 (n2214, n_1358, n2213);
  and g2427 (n2215, n_1358, n_1357);
  not g2428 (n_1359, n2212);
  not g2429 (n_1360, n2215);
  and g2430 (n2216, n_1359, n_1360);
  not g2431 (n_1361, n2214);
  not g2432 (n_1362, n2216);
  and g2433 (n2217, n_1361, n_1362);
  and g2434 (n2218, n_1253, n_1251);
  not g2435 (n_1363, n2218);
  and g2436 (n2219, n_1252, n_1363);
  and g2437 (n2220, n_1209, n_1253);
  and g2438 (n2221, n_1210, n2220);
  and g2439 (n2222, n_1254, n2221);
  and g2440 (n2223, n_1209, n_1207);
  not g2441 (n_1364, n2223);
  and g2442 (n2224, n_1208, n_1364);
  not g2443 (n_1365, n2222);
  not g2444 (n_1366, n2224);
  and g2445 (n2225, n_1365, n_1366);
  not g2450 (n_1367, n2225);
  not g2451 (n_1368, n2229);
  and g2452 (n2230, n_1367, n_1368);
  not g2453 (n_1369, n2230);
  and g2454 (n2231, n2219, n_1369);
  and g2455 (n2232, n_1365, n2224);
  and g2456 (n2233, n2222, n_1366);
  not g2457 (n_1370, n2232);
  not g2458 (n_1371, n2233);
  and g2459 (n2234, n_1370, n_1371);
  not g2460 (n_1372, n2219);
  not g2461 (n_1373, n2234);
  and g2462 (n2235, n_1372, n_1373);
  and g2463 (n2236, n_1351, n_1352);
  not g2464 (n_1374, n2235);
  and g2465 (n2237, n_1374, n2236);
  not g2466 (n_1375, n2231);
  and g2467 (n2238, n_1375, n2237);
  and g2468 (n2239, n_1375, n_1374);
  not g2469 (n_1376, n2236);
  not g2470 (n_1377, n2239);
  and g2471 (n2240, n_1376, n_1377);
  not g2472 (n_1378, n2238);
  not g2473 (n_1379, n2240);
  and g2474 (n2241, n_1378, n_1379);
  and g2475 (n2242, n_1345, n_1343);
  not g2476 (n_1380, n2242);
  and g2477 (n2243, n_1344, n_1380);
  and g2478 (n2244, n_1301, n_1345);
  and g2479 (n2245, n_1302, n2244);
  and g2480 (n2246, n_1346, n2245);
  and g2481 (n2247, n_1301, n_1299);
  not g2482 (n_1381, n2247);
  and g2483 (n2248, n_1300, n_1381);
  not g2484 (n_1382, n2246);
  and g2485 (n2249, n_1382, n2248);
  not g2486 (n_1383, n2248);
  and g2487 (n2250, n2246, n_1383);
  not g2488 (n_1384, n2249);
  not g2489 (n_1385, n2250);
  and g2490 (n2251, n_1384, n_1385);
  not g2491 (n_1386, n2243);
  not g2492 (n_1387, n2251);
  and g2493 (n2252, n_1386, n_1387);
  and g2494 (n2253, n_1382, n_1383);
  not g2499 (n_1388, n2253);
  not g2500 (n_1389, n2257);
  and g2501 (n2258, n_1388, n_1389);
  not g2502 (n_1390, n2258);
  and g2503 (n2259, n2243, n_1390);
  not g2504 (n_1391, n2252);
  not g2505 (n_1392, n2259);
  and g2506 (n2260, n_1391, n_1392);
  not g2507 (n_1393, n2241);
  and g2508 (n2261, n_1393, n2260);
  and g2509 (n2262, n_1374, n_1376);
  and g2510 (n2263, n_1375, n2262);
  and g2511 (n2264, n2236, n_1377);
  not g2512 (n_1394, n2263);
  not g2513 (n_1395, n2264);
  and g2514 (n2265, n_1394, n_1395);
  not g2515 (n_1396, n2260);
  not g2516 (n_1397, n2265);
  and g2517 (n2266, n_1396, n_1397);
  not g2518 (n_1398, n2261);
  not g2519 (n_1399, n2266);
  and g2520 (n2267, n_1398, n_1399);
  not g2521 (n_1400, n2217);
  and g2522 (n2268, n_1400, n2267);
  and g2523 (n2269, n_1357, n_1359);
  and g2524 (n2270, n_1358, n2269);
  and g2525 (n2271, n2212, n_1360);
  not g2526 (n_1401, n2270);
  not g2527 (n_1402, n2271);
  and g2528 (n2272, n_1401, n_1402);
  not g2529 (n_1403, n2267);
  not g2530 (n_1404, n2272);
  and g2531 (n2273, n_1403, n_1404);
  not g2532 (n_1405, n2268);
  not g2533 (n_1406, n2273);
  and g2534 (n2274, n_1405, n_1406);
  and g2535 (n2275, \A[814] , \A[815] );
  not g2536 (n_1409, \A[815] );
  and g2537 (n2276, \A[814] , n_1409);
  not g2538 (n_1410, \A[814] );
  and g2539 (n2277, n_1410, \A[815] );
  not g2540 (n_1411, n2276);
  not g2541 (n_1412, n2277);
  and g2542 (n2278, n_1411, n_1412);
  not g2543 (n_1414, n2278);
  and g2544 (n2279, \A[816] , n_1414);
  not g2545 (n_1415, n2275);
  not g2546 (n_1416, n2279);
  and g2547 (n2280, n_1415, n_1416);
  and g2548 (n2281, \A[811] , \A[812] );
  not g2549 (n_1419, \A[812] );
  and g2550 (n2282, \A[811] , n_1419);
  not g2551 (n_1420, \A[811] );
  and g2552 (n2283, n_1420, \A[812] );
  not g2553 (n_1421, n2282);
  not g2554 (n_1422, n2283);
  and g2555 (n2284, n_1421, n_1422);
  not g2556 (n_1424, n2284);
  and g2557 (n2285, \A[813] , n_1424);
  not g2558 (n_1425, n2281);
  not g2559 (n_1426, n2285);
  and g2560 (n2286, n_1425, n_1426);
  not g2561 (n_1427, n2286);
  and g2562 (n2287, n2280, n_1427);
  not g2563 (n_1428, n2280);
  and g2564 (n2288, n_1428, n2286);
  and g2565 (n2289, \A[813] , n_1421);
  and g2566 (n2290, n_1422, n2289);
  not g2567 (n_1429, \A[813] );
  and g2568 (n2291, n_1429, n_1424);
  not g2569 (n_1430, n2290);
  not g2570 (n_1431, n2291);
  and g2571 (n2292, n_1430, n_1431);
  and g2572 (n2293, \A[816] , n_1411);
  and g2573 (n2294, n_1412, n2293);
  not g2574 (n_1432, \A[816] );
  and g2575 (n2295, n_1432, n_1414);
  not g2576 (n_1433, n2294);
  not g2577 (n_1434, n2295);
  and g2578 (n2296, n_1433, n_1434);
  not g2579 (n_1435, n2292);
  not g2580 (n_1436, n2296);
  and g2581 (n2297, n_1435, n_1436);
  not g2582 (n_1437, n2288);
  and g2583 (n2298, n_1437, n2297);
  not g2584 (n_1438, n2287);
  and g2585 (n2299, n_1438, n2298);
  and g2586 (n2300, n_1438, n_1437);
  not g2587 (n_1439, n2297);
  not g2588 (n_1440, n2300);
  and g2589 (n2301, n_1439, n_1440);
  not g2590 (n_1441, n2299);
  not g2591 (n_1442, n2301);
  and g2592 (n2302, n_1441, n_1442);
  and g2593 (n2303, n_1435, n2296);
  and g2594 (n2304, n2292, n_1436);
  not g2595 (n_1443, n2303);
  not g2596 (n_1444, n2304);
  and g2597 (n2305, n_1443, n_1444);
  and g2598 (n2306, n2297, n_1440);
  and g2599 (n2307, n_1428, n_1427);
  not g2600 (n_1445, n2306);
  not g2601 (n_1446, n2307);
  and g2602 (n2308, n_1445, n_1446);
  not g2603 (n_1447, n2305);
  not g2604 (n_1448, n2308);
  and g2605 (n2309, n_1447, n_1448);
  not g2606 (n_1449, n2302);
  not g2607 (n_1450, n2309);
  and g2608 (n2310, n_1449, n_1450);
  and g2609 (n2311, n_1449, n_1448);
  and g2610 (n2312, \A[820] , \A[821] );
  not g2611 (n_1453, \A[821] );
  and g2612 (n2313, \A[820] , n_1453);
  not g2613 (n_1454, \A[820] );
  and g2614 (n2314, n_1454, \A[821] );
  not g2615 (n_1455, n2313);
  not g2616 (n_1456, n2314);
  and g2617 (n2315, n_1455, n_1456);
  not g2618 (n_1458, n2315);
  and g2619 (n2316, \A[822] , n_1458);
  not g2620 (n_1459, n2312);
  not g2621 (n_1460, n2316);
  and g2622 (n2317, n_1459, n_1460);
  and g2623 (n2318, \A[817] , \A[818] );
  not g2624 (n_1463, \A[818] );
  and g2625 (n2319, \A[817] , n_1463);
  not g2626 (n_1464, \A[817] );
  and g2627 (n2320, n_1464, \A[818] );
  not g2628 (n_1465, n2319);
  not g2629 (n_1466, n2320);
  and g2630 (n2321, n_1465, n_1466);
  not g2631 (n_1468, n2321);
  and g2632 (n2322, \A[819] , n_1468);
  not g2633 (n_1469, n2318);
  not g2634 (n_1470, n2322);
  and g2635 (n2323, n_1469, n_1470);
  not g2636 (n_1471, n2317);
  and g2637 (n2324, n_1471, n2323);
  not g2638 (n_1472, n2323);
  and g2639 (n2325, n2317, n_1472);
  not g2640 (n_1473, n2324);
  not g2641 (n_1474, n2325);
  and g2642 (n2326, n_1473, n_1474);
  and g2643 (n2327, \A[819] , n_1465);
  and g2644 (n2328, n_1466, n2327);
  not g2645 (n_1475, \A[819] );
  and g2646 (n2329, n_1475, n_1468);
  not g2647 (n_1476, n2328);
  not g2648 (n_1477, n2329);
  and g2649 (n2330, n_1476, n_1477);
  and g2650 (n2331, \A[822] , n_1455);
  and g2651 (n2332, n_1456, n2331);
  not g2652 (n_1478, \A[822] );
  and g2653 (n2333, n_1478, n_1458);
  not g2654 (n_1479, n2332);
  not g2655 (n_1480, n2333);
  and g2656 (n2334, n_1479, n_1480);
  not g2657 (n_1481, n2330);
  not g2658 (n_1482, n2334);
  and g2659 (n2335, n_1481, n_1482);
  not g2660 (n_1483, n2326);
  and g2661 (n2336, n_1483, n2335);
  and g2662 (n2337, n_1471, n_1472);
  not g2663 (n_1484, n2336);
  not g2664 (n_1485, n2337);
  and g2665 (n2338, n_1484, n_1485);
  and g2666 (n2339, n_1473, n2335);
  and g2667 (n2340, n_1474, n2339);
  not g2668 (n_1486, n2335);
  and g2669 (n2341, n_1483, n_1486);
  not g2670 (n_1487, n2340);
  not g2671 (n_1488, n2341);
  and g2672 (n2342, n_1487, n_1488);
  not g2673 (n_1489, n2338);
  not g2674 (n_1490, n2342);
  and g2675 (n2343, n_1489, n_1490);
  and g2676 (n2344, n_1481, n2334);
  and g2677 (n2345, n2330, n_1482);
  not g2678 (n_1491, n2344);
  not g2679 (n_1492, n2345);
  and g2680 (n2346, n_1491, n_1492);
  not g2681 (n_1493, n2346);
  and g2682 (n2347, n_1447, n_1493);
  not g2683 (n_1494, n2343);
  and g2684 (n2348, n_1494, n2347);
  not g2685 (n_1495, n2311);
  and g2686 (n2349, n_1495, n2348);
  and g2687 (n2350, n_1489, n_1493);
  not g2688 (n_1496, n2350);
  and g2689 (n2351, n_1490, n_1496);
  not g2690 (n_1497, n2349);
  not g2691 (n_1498, n2351);
  and g2692 (n2352, n_1497, n_1498);
  not g2697 (n_1499, n2352);
  not g2698 (n_1500, n2356);
  and g2699 (n2357, n_1499, n_1500);
  not g2700 (n_1501, n2357);
  and g2701 (n2358, n2310, n_1501);
  and g2702 (n2359, n_1497, n2351);
  and g2703 (n2360, n2349, n_1498);
  not g2704 (n_1502, n2359);
  not g2705 (n_1503, n2360);
  and g2706 (n2361, n_1502, n_1503);
  not g2707 (n_1504, n2310);
  not g2708 (n_1505, n2361);
  and g2709 (n2362, n_1504, n_1505);
  and g2710 (n2363, n_1494, n_1493);
  and g2711 (n2364, n_1447, n_1495);
  not g2712 (n_1506, n2363);
  and g2713 (n2365, n_1506, n2364);
  not g2714 (n_1507, n2364);
  and g2715 (n2366, n2363, n_1507);
  not g2716 (n_1508, n2365);
  not g2717 (n_1509, n2366);
  and g2718 (n2367, n_1508, n_1509);
  not g2719 (n_1511, \A[805] );
  and g2720 (n2368, n_1511, \A[806] );
  not g2721 (n_1513, \A[806] );
  and g2722 (n2369, \A[805] , n_1513);
  not g2723 (n_1515, n2369);
  and g2724 (n2370, \A[807] , n_1515);
  not g2725 (n_1516, n2368);
  and g2726 (n2371, n_1516, n2370);
  and g2727 (n2372, n_1516, n_1515);
  not g2728 (n_1517, \A[807] );
  not g2729 (n_1518, n2372);
  and g2730 (n2373, n_1517, n_1518);
  not g2731 (n_1519, n2371);
  not g2732 (n_1520, n2373);
  and g2733 (n2374, n_1519, n_1520);
  not g2734 (n_1522, \A[808] );
  and g2735 (n2375, n_1522, \A[809] );
  not g2736 (n_1524, \A[809] );
  and g2737 (n2376, \A[808] , n_1524);
  not g2738 (n_1526, n2376);
  and g2739 (n2377, \A[810] , n_1526);
  not g2740 (n_1527, n2375);
  and g2741 (n2378, n_1527, n2377);
  and g2742 (n2379, n_1527, n_1526);
  not g2743 (n_1528, \A[810] );
  not g2744 (n_1529, n2379);
  and g2745 (n2380, n_1528, n_1529);
  not g2746 (n_1530, n2378);
  not g2747 (n_1531, n2380);
  and g2748 (n2381, n_1530, n_1531);
  not g2749 (n_1532, n2374);
  and g2750 (n2382, n_1532, n2381);
  not g2751 (n_1533, n2381);
  and g2752 (n2383, n2374, n_1533);
  not g2753 (n_1534, n2382);
  not g2754 (n_1535, n2383);
  and g2755 (n2384, n_1534, n_1535);
  and g2756 (n2385, \A[808] , \A[809] );
  and g2757 (n2386, \A[810] , n_1529);
  not g2758 (n_1536, n2385);
  not g2759 (n_1537, n2386);
  and g2760 (n2387, n_1536, n_1537);
  and g2761 (n2388, \A[805] , \A[806] );
  and g2762 (n2389, \A[807] , n_1518);
  not g2763 (n_1538, n2388);
  not g2764 (n_1539, n2389);
  and g2765 (n2390, n_1538, n_1539);
  not g2766 (n_1540, n2387);
  and g2767 (n2391, n_1540, n2390);
  not g2768 (n_1541, n2390);
  and g2769 (n2392, n2387, n_1541);
  not g2770 (n_1542, n2391);
  not g2771 (n_1543, n2392);
  and g2772 (n2393, n_1542, n_1543);
  and g2773 (n2394, n_1532, n_1533);
  not g2774 (n_1544, n2393);
  and g2775 (n2395, n_1544, n2394);
  and g2776 (n2396, n_1540, n_1541);
  not g2777 (n_1545, n2395);
  not g2778 (n_1546, n2396);
  and g2779 (n2397, n_1545, n_1546);
  and g2780 (n2398, n_1542, n2394);
  and g2781 (n2399, n_1543, n2398);
  not g2782 (n_1547, n2394);
  and g2783 (n2400, n_1544, n_1547);
  not g2784 (n_1548, n2399);
  not g2785 (n_1549, n2400);
  and g2786 (n2401, n_1548, n_1549);
  not g2787 (n_1550, n2397);
  not g2788 (n_1551, n2401);
  and g2789 (n2402, n_1550, n_1551);
  not g2790 (n_1552, n2384);
  not g2791 (n_1553, n2402);
  and g2792 (n2403, n_1552, n_1553);
  not g2793 (n_1555, \A[799] );
  and g2794 (n2404, n_1555, \A[800] );
  not g2795 (n_1557, \A[800] );
  and g2796 (n2405, \A[799] , n_1557);
  not g2797 (n_1559, n2405);
  and g2798 (n2406, \A[801] , n_1559);
  not g2799 (n_1560, n2404);
  and g2800 (n2407, n_1560, n2406);
  and g2801 (n2408, n_1560, n_1559);
  not g2802 (n_1561, \A[801] );
  not g2803 (n_1562, n2408);
  and g2804 (n2409, n_1561, n_1562);
  not g2805 (n_1563, n2407);
  not g2806 (n_1564, n2409);
  and g2807 (n2410, n_1563, n_1564);
  not g2808 (n_1566, \A[802] );
  and g2809 (n2411, n_1566, \A[803] );
  not g2810 (n_1568, \A[803] );
  and g2811 (n2412, \A[802] , n_1568);
  not g2812 (n_1570, n2412);
  and g2813 (n2413, \A[804] , n_1570);
  not g2814 (n_1571, n2411);
  and g2815 (n2414, n_1571, n2413);
  and g2816 (n2415, n_1571, n_1570);
  not g2817 (n_1572, \A[804] );
  not g2818 (n_1573, n2415);
  and g2819 (n2416, n_1572, n_1573);
  not g2820 (n_1574, n2414);
  not g2821 (n_1575, n2416);
  and g2822 (n2417, n_1574, n_1575);
  not g2823 (n_1576, n2410);
  and g2824 (n2418, n_1576, n2417);
  not g2825 (n_1577, n2417);
  and g2826 (n2419, n2410, n_1577);
  not g2827 (n_1578, n2418);
  not g2828 (n_1579, n2419);
  and g2829 (n2420, n_1578, n_1579);
  and g2830 (n2421, \A[802] , \A[803] );
  and g2831 (n2422, \A[804] , n_1573);
  not g2832 (n_1580, n2421);
  not g2833 (n_1581, n2422);
  and g2834 (n2423, n_1580, n_1581);
  and g2835 (n2424, \A[799] , \A[800] );
  and g2836 (n2425, \A[801] , n_1562);
  not g2837 (n_1582, n2424);
  not g2838 (n_1583, n2425);
  and g2839 (n2426, n_1582, n_1583);
  not g2840 (n_1584, n2423);
  and g2841 (n2427, n_1584, n2426);
  not g2842 (n_1585, n2426);
  and g2843 (n2428, n2423, n_1585);
  not g2844 (n_1586, n2427);
  not g2845 (n_1587, n2428);
  and g2846 (n2429, n_1586, n_1587);
  and g2847 (n2430, n_1576, n_1577);
  not g2848 (n_1588, n2429);
  and g2849 (n2431, n_1588, n2430);
  and g2850 (n2432, n_1584, n_1585);
  not g2851 (n_1589, n2431);
  not g2852 (n_1590, n2432);
  and g2853 (n2433, n_1589, n_1590);
  and g2854 (n2434, n_1586, n2430);
  and g2855 (n2435, n_1587, n2434);
  not g2856 (n_1591, n2430);
  and g2857 (n2436, n_1588, n_1591);
  not g2858 (n_1592, n2435);
  not g2859 (n_1593, n2436);
  and g2860 (n2437, n_1592, n_1593);
  not g2861 (n_1594, n2433);
  not g2862 (n_1595, n2437);
  and g2863 (n2438, n_1594, n_1595);
  not g2864 (n_1596, n2420);
  not g2865 (n_1597, n2438);
  and g2866 (n2439, n_1596, n_1597);
  not g2867 (n_1598, n2403);
  and g2868 (n2440, n_1598, n2439);
  not g2869 (n_1599, n2439);
  and g2870 (n2441, n2403, n_1599);
  not g2871 (n_1600, n2440);
  not g2872 (n_1601, n2441);
  and g2873 (n2442, n_1600, n_1601);
  not g2874 (n_1602, n2367);
  not g2875 (n_1603, n2442);
  and g2876 (n2443, n_1602, n_1603);
  not g2877 (n_1604, n2362);
  and g2878 (n2444, n_1604, n2443);
  not g2879 (n_1605, n2358);
  and g2880 (n2445, n_1605, n2444);
  and g2881 (n2446, n_1605, n_1604);
  not g2882 (n_1606, n2443);
  not g2883 (n_1607, n2446);
  and g2884 (n2447, n_1606, n_1607);
  not g2885 (n_1608, n2445);
  not g2886 (n_1609, n2447);
  and g2887 (n2448, n_1608, n_1609);
  and g2888 (n2449, n_1596, n_1594);
  not g2889 (n_1610, n2449);
  and g2890 (n2450, n_1595, n_1610);
  and g2891 (n2451, n_1552, n_1596);
  and g2892 (n2452, n_1553, n2451);
  and g2893 (n2453, n_1597, n2452);
  and g2894 (n2454, n_1552, n_1550);
  not g2895 (n_1611, n2454);
  and g2896 (n2455, n_1551, n_1611);
  not g2897 (n_1612, n2453);
  and g2898 (n2456, n_1612, n2455);
  not g2899 (n_1613, n2455);
  and g2900 (n2457, n2453, n_1613);
  not g2901 (n_1614, n2456);
  not g2902 (n_1615, n2457);
  and g2903 (n2458, n_1614, n_1615);
  not g2904 (n_1616, n2450);
  not g2905 (n_1617, n2458);
  and g2906 (n2459, n_1616, n_1617);
  and g2907 (n2460, n_1612, n_1613);
  not g2912 (n_1618, n2460);
  not g2913 (n_1619, n2464);
  and g2914 (n2465, n_1618, n_1619);
  not g2915 (n_1620, n2465);
  and g2916 (n2466, n2450, n_1620);
  not g2917 (n_1621, n2459);
  not g2918 (n_1622, n2466);
  and g2919 (n2467, n_1621, n_1622);
  not g2920 (n_1623, n2448);
  and g2921 (n2468, n_1623, n2467);
  and g2922 (n2469, n_1604, n_1606);
  and g2923 (n2470, n_1605, n2469);
  and g2924 (n2471, n2443, n_1607);
  not g2925 (n_1624, n2470);
  not g2926 (n_1625, n2471);
  and g2927 (n2472, n_1624, n_1625);
  not g2928 (n_1626, n2467);
  not g2929 (n_1627, n2472);
  and g2930 (n2473, n_1626, n_1627);
  not g2931 (n_1628, n2468);
  not g2932 (n_1629, n2473);
  and g2933 (n2474, n_1628, n_1629);
  and g2934 (n2475, \A[826] , \A[827] );
  not g2935 (n_1632, \A[827] );
  and g2936 (n2476, \A[826] , n_1632);
  not g2937 (n_1633, \A[826] );
  and g2938 (n2477, n_1633, \A[827] );
  not g2939 (n_1634, n2476);
  not g2940 (n_1635, n2477);
  and g2941 (n2478, n_1634, n_1635);
  not g2942 (n_1637, n2478);
  and g2943 (n2479, \A[828] , n_1637);
  not g2944 (n_1638, n2475);
  not g2945 (n_1639, n2479);
  and g2946 (n2480, n_1638, n_1639);
  and g2947 (n2481, \A[823] , \A[824] );
  not g2948 (n_1642, \A[824] );
  and g2949 (n2482, \A[823] , n_1642);
  not g2950 (n_1643, \A[823] );
  and g2951 (n2483, n_1643, \A[824] );
  not g2952 (n_1644, n2482);
  not g2953 (n_1645, n2483);
  and g2954 (n2484, n_1644, n_1645);
  not g2955 (n_1647, n2484);
  and g2956 (n2485, \A[825] , n_1647);
  not g2957 (n_1648, n2481);
  not g2958 (n_1649, n2485);
  and g2959 (n2486, n_1648, n_1649);
  not g2960 (n_1650, n2486);
  and g2961 (n2487, n2480, n_1650);
  not g2962 (n_1651, n2480);
  and g2963 (n2488, n_1651, n2486);
  and g2964 (n2489, \A[825] , n_1644);
  and g2965 (n2490, n_1645, n2489);
  not g2966 (n_1652, \A[825] );
  and g2967 (n2491, n_1652, n_1647);
  not g2968 (n_1653, n2490);
  not g2969 (n_1654, n2491);
  and g2970 (n2492, n_1653, n_1654);
  and g2971 (n2493, \A[828] , n_1634);
  and g2972 (n2494, n_1635, n2493);
  not g2973 (n_1655, \A[828] );
  and g2974 (n2495, n_1655, n_1637);
  not g2975 (n_1656, n2494);
  not g2976 (n_1657, n2495);
  and g2977 (n2496, n_1656, n_1657);
  not g2978 (n_1658, n2492);
  not g2979 (n_1659, n2496);
  and g2980 (n2497, n_1658, n_1659);
  not g2981 (n_1660, n2488);
  and g2982 (n2498, n_1660, n2497);
  not g2983 (n_1661, n2487);
  and g2984 (n2499, n_1661, n2498);
  and g2985 (n2500, n_1661, n_1660);
  not g2986 (n_1662, n2497);
  not g2987 (n_1663, n2500);
  and g2988 (n2501, n_1662, n_1663);
  not g2989 (n_1664, n2499);
  not g2990 (n_1665, n2501);
  and g2991 (n2502, n_1664, n_1665);
  and g2992 (n2503, n_1658, n2496);
  and g2993 (n2504, n2492, n_1659);
  not g2994 (n_1666, n2503);
  not g2995 (n_1667, n2504);
  and g2996 (n2505, n_1666, n_1667);
  and g2997 (n2506, n2497, n_1663);
  and g2998 (n2507, n_1651, n_1650);
  not g2999 (n_1668, n2506);
  not g3000 (n_1669, n2507);
  and g3001 (n2508, n_1668, n_1669);
  not g3002 (n_1670, n2505);
  not g3003 (n_1671, n2508);
  and g3004 (n2509, n_1670, n_1671);
  not g3005 (n_1672, n2502);
  not g3006 (n_1673, n2509);
  and g3007 (n2510, n_1672, n_1673);
  and g3008 (n2511, n_1672, n_1671);
  and g3009 (n2512, \A[832] , \A[833] );
  not g3010 (n_1676, \A[833] );
  and g3011 (n2513, \A[832] , n_1676);
  not g3012 (n_1677, \A[832] );
  and g3013 (n2514, n_1677, \A[833] );
  not g3014 (n_1678, n2513);
  not g3015 (n_1679, n2514);
  and g3016 (n2515, n_1678, n_1679);
  not g3017 (n_1681, n2515);
  and g3018 (n2516, \A[834] , n_1681);
  not g3019 (n_1682, n2512);
  not g3020 (n_1683, n2516);
  and g3021 (n2517, n_1682, n_1683);
  and g3022 (n2518, \A[829] , \A[830] );
  not g3023 (n_1686, \A[830] );
  and g3024 (n2519, \A[829] , n_1686);
  not g3025 (n_1687, \A[829] );
  and g3026 (n2520, n_1687, \A[830] );
  not g3027 (n_1688, n2519);
  not g3028 (n_1689, n2520);
  and g3029 (n2521, n_1688, n_1689);
  not g3030 (n_1691, n2521);
  and g3031 (n2522, \A[831] , n_1691);
  not g3032 (n_1692, n2518);
  not g3033 (n_1693, n2522);
  and g3034 (n2523, n_1692, n_1693);
  not g3035 (n_1694, n2517);
  and g3036 (n2524, n_1694, n2523);
  not g3037 (n_1695, n2523);
  and g3038 (n2525, n2517, n_1695);
  not g3039 (n_1696, n2524);
  not g3040 (n_1697, n2525);
  and g3041 (n2526, n_1696, n_1697);
  and g3042 (n2527, \A[831] , n_1688);
  and g3043 (n2528, n_1689, n2527);
  not g3044 (n_1698, \A[831] );
  and g3045 (n2529, n_1698, n_1691);
  not g3046 (n_1699, n2528);
  not g3047 (n_1700, n2529);
  and g3048 (n2530, n_1699, n_1700);
  and g3049 (n2531, \A[834] , n_1678);
  and g3050 (n2532, n_1679, n2531);
  not g3051 (n_1701, \A[834] );
  and g3052 (n2533, n_1701, n_1681);
  not g3053 (n_1702, n2532);
  not g3054 (n_1703, n2533);
  and g3055 (n2534, n_1702, n_1703);
  not g3056 (n_1704, n2530);
  not g3057 (n_1705, n2534);
  and g3058 (n2535, n_1704, n_1705);
  not g3059 (n_1706, n2526);
  and g3060 (n2536, n_1706, n2535);
  and g3061 (n2537, n_1694, n_1695);
  not g3062 (n_1707, n2536);
  not g3063 (n_1708, n2537);
  and g3064 (n2538, n_1707, n_1708);
  and g3065 (n2539, n_1696, n2535);
  and g3066 (n2540, n_1697, n2539);
  not g3067 (n_1709, n2535);
  and g3068 (n2541, n_1706, n_1709);
  not g3069 (n_1710, n2540);
  not g3070 (n_1711, n2541);
  and g3071 (n2542, n_1710, n_1711);
  not g3072 (n_1712, n2538);
  not g3073 (n_1713, n2542);
  and g3074 (n2543, n_1712, n_1713);
  and g3075 (n2544, n_1704, n2534);
  and g3076 (n2545, n2530, n_1705);
  not g3077 (n_1714, n2544);
  not g3078 (n_1715, n2545);
  and g3079 (n2546, n_1714, n_1715);
  not g3080 (n_1716, n2546);
  and g3081 (n2547, n_1670, n_1716);
  not g3082 (n_1717, n2543);
  and g3083 (n2548, n_1717, n2547);
  not g3084 (n_1718, n2511);
  and g3085 (n2549, n_1718, n2548);
  and g3086 (n2550, n_1712, n_1716);
  not g3087 (n_1719, n2550);
  and g3088 (n2551, n_1713, n_1719);
  not g3089 (n_1720, n2549);
  and g3090 (n2552, n_1720, n2551);
  not g3091 (n_1721, n2551);
  and g3092 (n2553, n2549, n_1721);
  not g3093 (n_1722, n2552);
  not g3094 (n_1723, n2553);
  and g3095 (n2554, n_1722, n_1723);
  not g3096 (n_1724, n2510);
  not g3097 (n_1725, n2554);
  and g3098 (n2555, n_1724, n_1725);
  and g3099 (n2556, n_1720, n_1721);
  not g3104 (n_1726, n2556);
  not g3105 (n_1727, n2560);
  and g3106 (n2561, n_1726, n_1727);
  not g3107 (n_1728, n2561);
  and g3108 (n2562, n2510, n_1728);
  not g3109 (n_1729, n2555);
  not g3110 (n_1730, n2562);
  and g3111 (n2563, n_1729, n_1730);
  and g3112 (n2564, \A[838] , \A[839] );
  not g3113 (n_1733, \A[839] );
  and g3114 (n2565, \A[838] , n_1733);
  not g3115 (n_1734, \A[838] );
  and g3116 (n2566, n_1734, \A[839] );
  not g3117 (n_1735, n2565);
  not g3118 (n_1736, n2566);
  and g3119 (n2567, n_1735, n_1736);
  not g3120 (n_1738, n2567);
  and g3121 (n2568, \A[840] , n_1738);
  not g3122 (n_1739, n2564);
  not g3123 (n_1740, n2568);
  and g3124 (n2569, n_1739, n_1740);
  and g3125 (n2570, \A[835] , \A[836] );
  not g3126 (n_1743, \A[836] );
  and g3127 (n2571, \A[835] , n_1743);
  not g3128 (n_1744, \A[835] );
  and g3129 (n2572, n_1744, \A[836] );
  not g3130 (n_1745, n2571);
  not g3131 (n_1746, n2572);
  and g3132 (n2573, n_1745, n_1746);
  not g3133 (n_1748, n2573);
  and g3134 (n2574, \A[837] , n_1748);
  not g3135 (n_1749, n2570);
  not g3136 (n_1750, n2574);
  and g3137 (n2575, n_1749, n_1750);
  not g3138 (n_1751, n2575);
  and g3139 (n2576, n2569, n_1751);
  not g3140 (n_1752, n2569);
  and g3141 (n2577, n_1752, n2575);
  and g3142 (n2578, \A[837] , n_1745);
  and g3143 (n2579, n_1746, n2578);
  not g3144 (n_1753, \A[837] );
  and g3145 (n2580, n_1753, n_1748);
  not g3146 (n_1754, n2579);
  not g3147 (n_1755, n2580);
  and g3148 (n2581, n_1754, n_1755);
  and g3149 (n2582, \A[840] , n_1735);
  and g3150 (n2583, n_1736, n2582);
  not g3151 (n_1756, \A[840] );
  and g3152 (n2584, n_1756, n_1738);
  not g3153 (n_1757, n2583);
  not g3154 (n_1758, n2584);
  and g3155 (n2585, n_1757, n_1758);
  not g3156 (n_1759, n2581);
  not g3157 (n_1760, n2585);
  and g3158 (n2586, n_1759, n_1760);
  not g3159 (n_1761, n2577);
  and g3160 (n2587, n_1761, n2586);
  not g3161 (n_1762, n2576);
  and g3162 (n2588, n_1762, n2587);
  and g3163 (n2589, n_1762, n_1761);
  not g3164 (n_1763, n2586);
  not g3165 (n_1764, n2589);
  and g3166 (n2590, n_1763, n_1764);
  not g3167 (n_1765, n2588);
  not g3168 (n_1766, n2590);
  and g3169 (n2591, n_1765, n_1766);
  and g3170 (n2592, n_1759, n2585);
  and g3171 (n2593, n2581, n_1760);
  not g3172 (n_1767, n2592);
  not g3173 (n_1768, n2593);
  and g3174 (n2594, n_1767, n_1768);
  and g3175 (n2595, n2586, n_1764);
  and g3176 (n2596, n_1752, n_1751);
  not g3177 (n_1769, n2595);
  not g3178 (n_1770, n2596);
  and g3179 (n2597, n_1769, n_1770);
  not g3180 (n_1771, n2594);
  not g3181 (n_1772, n2597);
  and g3182 (n2598, n_1771, n_1772);
  not g3183 (n_1773, n2591);
  not g3184 (n_1774, n2598);
  and g3185 (n2599, n_1773, n_1774);
  and g3186 (n2600, n_1773, n_1772);
  and g3187 (n2601, \A[844] , \A[845] );
  not g3188 (n_1777, \A[845] );
  and g3189 (n2602, \A[844] , n_1777);
  not g3190 (n_1778, \A[844] );
  and g3191 (n2603, n_1778, \A[845] );
  not g3192 (n_1779, n2602);
  not g3193 (n_1780, n2603);
  and g3194 (n2604, n_1779, n_1780);
  not g3195 (n_1782, n2604);
  and g3196 (n2605, \A[846] , n_1782);
  not g3197 (n_1783, n2601);
  not g3198 (n_1784, n2605);
  and g3199 (n2606, n_1783, n_1784);
  and g3200 (n2607, \A[841] , \A[842] );
  not g3201 (n_1787, \A[842] );
  and g3202 (n2608, \A[841] , n_1787);
  not g3203 (n_1788, \A[841] );
  and g3204 (n2609, n_1788, \A[842] );
  not g3205 (n_1789, n2608);
  not g3206 (n_1790, n2609);
  and g3207 (n2610, n_1789, n_1790);
  not g3208 (n_1792, n2610);
  and g3209 (n2611, \A[843] , n_1792);
  not g3210 (n_1793, n2607);
  not g3211 (n_1794, n2611);
  and g3212 (n2612, n_1793, n_1794);
  not g3213 (n_1795, n2606);
  and g3214 (n2613, n_1795, n2612);
  not g3215 (n_1796, n2612);
  and g3216 (n2614, n2606, n_1796);
  not g3217 (n_1797, n2613);
  not g3218 (n_1798, n2614);
  and g3219 (n2615, n_1797, n_1798);
  and g3220 (n2616, \A[843] , n_1789);
  and g3221 (n2617, n_1790, n2616);
  not g3222 (n_1799, \A[843] );
  and g3223 (n2618, n_1799, n_1792);
  not g3224 (n_1800, n2617);
  not g3225 (n_1801, n2618);
  and g3226 (n2619, n_1800, n_1801);
  and g3227 (n2620, \A[846] , n_1779);
  and g3228 (n2621, n_1780, n2620);
  not g3229 (n_1802, \A[846] );
  and g3230 (n2622, n_1802, n_1782);
  not g3231 (n_1803, n2621);
  not g3232 (n_1804, n2622);
  and g3233 (n2623, n_1803, n_1804);
  not g3234 (n_1805, n2619);
  not g3235 (n_1806, n2623);
  and g3236 (n2624, n_1805, n_1806);
  not g3237 (n_1807, n2615);
  and g3238 (n2625, n_1807, n2624);
  and g3239 (n2626, n_1795, n_1796);
  not g3240 (n_1808, n2625);
  not g3241 (n_1809, n2626);
  and g3242 (n2627, n_1808, n_1809);
  and g3243 (n2628, n_1797, n2624);
  and g3244 (n2629, n_1798, n2628);
  not g3245 (n_1810, n2624);
  and g3246 (n2630, n_1807, n_1810);
  not g3247 (n_1811, n2629);
  not g3248 (n_1812, n2630);
  and g3249 (n2631, n_1811, n_1812);
  not g3250 (n_1813, n2627);
  not g3251 (n_1814, n2631);
  and g3252 (n2632, n_1813, n_1814);
  and g3253 (n2633, n_1805, n2623);
  and g3254 (n2634, n2619, n_1806);
  not g3255 (n_1815, n2633);
  not g3256 (n_1816, n2634);
  and g3257 (n2635, n_1815, n_1816);
  not g3258 (n_1817, n2635);
  and g3259 (n2636, n_1771, n_1817);
  not g3260 (n_1818, n2632);
  and g3261 (n2637, n_1818, n2636);
  not g3262 (n_1819, n2600);
  and g3263 (n2638, n_1819, n2637);
  and g3264 (n2639, n_1813, n_1817);
  not g3265 (n_1820, n2639);
  and g3266 (n2640, n_1814, n_1820);
  not g3267 (n_1821, n2638);
  not g3268 (n_1822, n2640);
  and g3269 (n2641, n_1821, n_1822);
  not g3274 (n_1823, n2641);
  not g3275 (n_1824, n2645);
  and g3276 (n2646, n_1823, n_1824);
  not g3277 (n_1825, n2646);
  and g3278 (n2647, n2599, n_1825);
  and g3279 (n2648, n_1821, n2640);
  and g3280 (n2649, n2638, n_1822);
  not g3281 (n_1826, n2648);
  not g3282 (n_1827, n2649);
  and g3283 (n2650, n_1826, n_1827);
  not g3284 (n_1828, n2599);
  not g3285 (n_1829, n2650);
  and g3286 (n2651, n_1828, n_1829);
  and g3287 (n2652, n_1818, n_1817);
  and g3288 (n2653, n_1771, n_1819);
  not g3289 (n_1830, n2652);
  and g3290 (n2654, n_1830, n2653);
  not g3291 (n_1831, n2653);
  and g3292 (n2655, n2652, n_1831);
  not g3293 (n_1832, n2654);
  not g3294 (n_1833, n2655);
  and g3295 (n2656, n_1832, n_1833);
  and g3296 (n2657, n_1717, n_1716);
  and g3297 (n2658, n_1670, n_1718);
  not g3298 (n_1834, n2657);
  and g3299 (n2659, n_1834, n2658);
  not g3300 (n_1835, n2658);
  and g3301 (n2660, n2657, n_1835);
  not g3302 (n_1836, n2659);
  not g3303 (n_1837, n2660);
  and g3304 (n2661, n_1836, n_1837);
  not g3305 (n_1838, n2656);
  not g3306 (n_1839, n2661);
  and g3307 (n2662, n_1838, n_1839);
  not g3308 (n_1840, n2651);
  not g3309 (n_1841, n2662);
  and g3310 (n2663, n_1840, n_1841);
  not g3311 (n_1842, n2647);
  and g3312 (n2664, n_1842, n2663);
  and g3313 (n2665, n_1842, n_1840);
  not g3314 (n_1843, n2665);
  and g3315 (n2666, n2662, n_1843);
  not g3316 (n_1844, n2664);
  not g3317 (n_1845, n2666);
  and g3318 (n2667, n_1844, n_1845);
  not g3319 (n_1846, n2563);
  not g3320 (n_1847, n2667);
  and g3321 (n2668, n_1846, n_1847);
  and g3322 (n2669, n_1840, n2662);
  and g3323 (n2670, n_1842, n2669);
  and g3324 (n2671, n_1841, n_1843);
  not g3325 (n_1848, n2670);
  not g3326 (n_1849, n2671);
  and g3327 (n2672, n_1848, n_1849);
  not g3328 (n_1850, n2672);
  and g3329 (n2673, n2563, n_1850);
  and g3330 (n2674, n_1838, n2661);
  and g3331 (n2675, n2656, n_1839);
  not g3332 (n_1851, n2674);
  not g3333 (n_1852, n2675);
  and g3334 (n2676, n_1851, n_1852);
  and g3335 (n2677, n_1602, n2442);
  and g3336 (n2678, n2367, n_1603);
  not g3337 (n_1853, n2677);
  not g3338 (n_1854, n2678);
  and g3339 (n2679, n_1853, n_1854);
  not g3340 (n_1855, n2676);
  not g3341 (n_1856, n2679);
  and g3342 (n2680, n_1855, n_1856);
  not g3343 (n_1857, n2673);
  not g3344 (n_1858, n2680);
  and g3345 (n2681, n_1857, n_1858);
  not g3346 (n_1859, n2668);
  and g3347 (n2682, n_1859, n2681);
  and g3348 (n2683, n_1859, n_1857);
  not g3349 (n_1860, n2683);
  and g3350 (n2684, n2680, n_1860);
  not g3351 (n_1861, n2682);
  not g3352 (n_1862, n2684);
  and g3353 (n2685, n_1861, n_1862);
  not g3354 (n_1863, n2474);
  not g3355 (n_1864, n2685);
  and g3356 (n2686, n_1863, n_1864);
  and g3357 (n2687, n_1857, n2680);
  and g3358 (n2688, n_1859, n2687);
  and g3359 (n2689, n_1858, n_1860);
  not g3360 (n_1865, n2688);
  not g3361 (n_1866, n2689);
  and g3362 (n2690, n_1865, n_1866);
  not g3363 (n_1867, n2690);
  and g3364 (n2691, n2474, n_1867);
  and g3365 (n2692, n_1855, n2679);
  and g3366 (n2693, n2676, n_1856);
  not g3367 (n_1868, n2692);
  not g3368 (n_1869, n2693);
  and g3369 (n2694, n_1868, n_1869);
  and g3370 (n2695, n_1355, n2211);
  and g3371 (n2696, n2058, n_1356);
  not g3372 (n_1870, n2695);
  not g3373 (n_1871, n2696);
  and g3374 (n2697, n_1870, n_1871);
  not g3375 (n_1872, n2694);
  not g3376 (n_1873, n2697);
  and g3377 (n2698, n_1872, n_1873);
  not g3378 (n_1874, n2691);
  not g3379 (n_1875, n2698);
  and g3380 (n2699, n_1874, n_1875);
  not g3381 (n_1876, n2686);
  and g3382 (n2700, n_1876, n2699);
  and g3383 (n2701, n_1876, n_1874);
  not g3384 (n_1877, n2701);
  and g3385 (n2702, n2698, n_1877);
  not g3386 (n_1878, n2700);
  not g3387 (n_1879, n2702);
  and g3388 (n2703, n_1878, n_1879);
  not g3389 (n_1880, n2274);
  not g3390 (n_1881, n2703);
  and g3391 (n2704, n_1880, n_1881);
  and g3392 (n2705, n_1874, n2698);
  and g3393 (n2706, n_1876, n2705);
  and g3394 (n2707, n_1875, n_1877);
  not g3395 (n_1882, n2706);
  not g3396 (n_1883, n2707);
  and g3397 (n2708, n_1882, n_1883);
  not g3398 (n_1884, n2708);
  and g3399 (n2709, n2274, n_1884);
  and g3400 (n2710, n_1872, n2697);
  and g3401 (n2711, n2694, n_1873);
  not g3402 (n_1885, n2710);
  not g3403 (n_1886, n2711);
  and g3404 (n2712, n_1885, n_1886);
  and g3405 (n2713, n_844, n1731);
  and g3406 (n2714, n1422, n_845);
  not g3407 (n_1887, n2713);
  not g3408 (n_1888, n2714);
  and g3409 (n2715, n_1887, n_1888);
  not g3410 (n_1889, n2712);
  not g3411 (n_1890, n2715);
  and g3412 (n2716, n_1889, n_1890);
  not g3413 (n_1891, n2709);
  not g3414 (n_1892, n2716);
  and g3415 (n2717, n_1891, n_1892);
  not g3416 (n_1893, n2704);
  and g3417 (n2718, n_1893, n2717);
  and g3418 (n2719, n_1893, n_1891);
  not g3419 (n_1894, n2719);
  and g3420 (n2720, n2716, n_1894);
  not g3421 (n_1895, n2718);
  not g3422 (n_1896, n2720);
  and g3423 (n2721, n_1895, n_1896);
  not g3424 (n_1897, n1856);
  not g3425 (n_1898, n2721);
  and g3426 (n2722, n_1897, n_1898);
  and g3427 (n2723, n_1891, n2716);
  and g3428 (n2724, n_1893, n2723);
  and g3429 (n2725, n_1892, n_1894);
  not g3430 (n_1899, n2724);
  not g3431 (n_1900, n2725);
  and g3432 (n2726, n_1899, n_1900);
  not g3433 (n_1901, n2726);
  and g3434 (n2727, n1856, n_1901);
  not g3435 (n_1903, \A[469] );
  and g3436 (n2728, n_1903, \A[470] );
  not g3437 (n_1905, \A[470] );
  and g3438 (n2729, \A[469] , n_1905);
  not g3439 (n_1907, n2729);
  and g3440 (n2730, \A[471] , n_1907);
  not g3441 (n_1908, n2728);
  and g3442 (n2731, n_1908, n2730);
  and g3443 (n2732, n_1908, n_1907);
  not g3444 (n_1909, \A[471] );
  not g3445 (n_1910, n2732);
  and g3446 (n2733, n_1909, n_1910);
  not g3447 (n_1911, n2731);
  not g3448 (n_1912, n2733);
  and g3449 (n2734, n_1911, n_1912);
  not g3450 (n_1914, \A[472] );
  and g3451 (n2735, n_1914, \A[473] );
  not g3452 (n_1916, \A[473] );
  and g3453 (n2736, \A[472] , n_1916);
  not g3454 (n_1918, n2736);
  and g3455 (n2737, \A[474] , n_1918);
  not g3456 (n_1919, n2735);
  and g3457 (n2738, n_1919, n2737);
  and g3458 (n2739, n_1919, n_1918);
  not g3459 (n_1920, \A[474] );
  not g3460 (n_1921, n2739);
  and g3461 (n2740, n_1920, n_1921);
  not g3462 (n_1922, n2738);
  not g3463 (n_1923, n2740);
  and g3464 (n2741, n_1922, n_1923);
  not g3465 (n_1924, n2734);
  and g3466 (n2742, n_1924, n2741);
  not g3467 (n_1925, n2741);
  and g3468 (n2743, n2734, n_1925);
  not g3469 (n_1926, n2742);
  not g3470 (n_1927, n2743);
  and g3471 (n2744, n_1926, n_1927);
  and g3472 (n2745, \A[472] , \A[473] );
  and g3473 (n2746, \A[474] , n_1921);
  not g3474 (n_1928, n2745);
  not g3475 (n_1929, n2746);
  and g3476 (n2747, n_1928, n_1929);
  and g3477 (n2748, \A[469] , \A[470] );
  and g3478 (n2749, \A[471] , n_1910);
  not g3479 (n_1930, n2748);
  not g3480 (n_1931, n2749);
  and g3481 (n2750, n_1930, n_1931);
  not g3482 (n_1932, n2747);
  and g3483 (n2751, n_1932, n2750);
  not g3484 (n_1933, n2750);
  and g3485 (n2752, n2747, n_1933);
  not g3486 (n_1934, n2751);
  not g3487 (n_1935, n2752);
  and g3488 (n2753, n_1934, n_1935);
  and g3489 (n2754, n_1924, n_1925);
  not g3490 (n_1936, n2753);
  and g3491 (n2755, n_1936, n2754);
  and g3492 (n2756, n_1932, n_1933);
  not g3493 (n_1937, n2755);
  not g3494 (n_1938, n2756);
  and g3495 (n2757, n_1937, n_1938);
  and g3496 (n2758, n_1934, n2754);
  and g3497 (n2759, n_1935, n2758);
  not g3498 (n_1939, n2754);
  and g3499 (n2760, n_1936, n_1939);
  not g3500 (n_1940, n2759);
  not g3501 (n_1941, n2760);
  and g3502 (n2761, n_1940, n_1941);
  not g3503 (n_1942, n2757);
  not g3504 (n_1943, n2761);
  and g3505 (n2762, n_1942, n_1943);
  not g3506 (n_1944, n2744);
  not g3507 (n_1945, n2762);
  and g3508 (n2763, n_1944, n_1945);
  not g3509 (n_1947, \A[466] );
  and g3510 (n2764, n_1947, \A[467] );
  not g3511 (n_1949, \A[467] );
  and g3512 (n2765, \A[466] , n_1949);
  not g3513 (n_1951, n2765);
  and g3514 (n2766, \A[468] , n_1951);
  not g3515 (n_1952, n2764);
  and g3516 (n2767, n_1952, n2766);
  and g3517 (n2768, n_1952, n_1951);
  not g3518 (n_1953, \A[468] );
  not g3519 (n_1954, n2768);
  and g3520 (n2769, n_1953, n_1954);
  not g3521 (n_1955, n2767);
  not g3522 (n_1956, n2769);
  and g3523 (n2770, n_1955, n_1956);
  not g3524 (n_1958, \A[463] );
  and g3525 (n2771, n_1958, \A[464] );
  not g3526 (n_1960, \A[464] );
  and g3527 (n2772, \A[463] , n_1960);
  not g3528 (n_1962, n2772);
  and g3529 (n2773, \A[465] , n_1962);
  not g3530 (n_1963, n2771);
  and g3531 (n2774, n_1963, n2773);
  and g3532 (n2775, n_1963, n_1962);
  not g3533 (n_1964, \A[465] );
  not g3534 (n_1965, n2775);
  and g3535 (n2776, n_1964, n_1965);
  not g3536 (n_1966, n2774);
  not g3537 (n_1967, n2776);
  and g3538 (n2777, n_1966, n_1967);
  not g3539 (n_1968, n2770);
  and g3540 (n2778, n_1968, n2777);
  not g3541 (n_1969, n2777);
  and g3542 (n2779, n2770, n_1969);
  not g3543 (n_1970, n2778);
  not g3544 (n_1971, n2779);
  and g3545 (n2780, n_1970, n_1971);
  and g3546 (n2781, \A[466] , \A[467] );
  and g3547 (n2782, \A[468] , n_1954);
  not g3548 (n_1972, n2781);
  not g3549 (n_1973, n2782);
  and g3550 (n2783, n_1972, n_1973);
  and g3551 (n2784, \A[463] , \A[464] );
  and g3552 (n2785, \A[465] , n_1965);
  not g3553 (n_1974, n2784);
  not g3554 (n_1975, n2785);
  and g3555 (n2786, n_1974, n_1975);
  not g3556 (n_1976, n2786);
  and g3557 (n2787, n2783, n_1976);
  not g3558 (n_1977, n2783);
  and g3559 (n2788, n_1977, n2786);
  and g3560 (n2789, n_1968, n_1969);
  not g3561 (n_1978, n2788);
  and g3562 (n2790, n_1978, n2789);
  not g3563 (n_1979, n2787);
  and g3564 (n2791, n_1979, n2790);
  and g3565 (n2792, n_1979, n_1978);
  not g3566 (n_1980, n2789);
  not g3567 (n_1981, n2792);
  and g3568 (n2793, n_1980, n_1981);
  not g3569 (n_1982, n2791);
  not g3570 (n_1983, n2793);
  and g3571 (n2794, n_1982, n_1983);
  and g3572 (n2795, n2789, n_1981);
  and g3573 (n2796, n_1977, n_1976);
  not g3574 (n_1984, n2795);
  not g3575 (n_1985, n2796);
  and g3576 (n2797, n_1984, n_1985);
  not g3577 (n_1986, n2794);
  not g3578 (n_1987, n2797);
  and g3579 (n2798, n_1986, n_1987);
  not g3580 (n_1988, n2780);
  not g3581 (n_1989, n2798);
  and g3582 (n2799, n_1988, n_1989);
  not g3583 (n_1990, n2763);
  and g3584 (n2800, n_1990, n2799);
  not g3585 (n_1991, n2799);
  and g3586 (n2801, n2763, n_1991);
  not g3587 (n_1992, n2800);
  not g3588 (n_1993, n2801);
  and g3589 (n2802, n_1992, n_1993);
  not g3590 (n_1995, \A[481] );
  and g3591 (n2803, n_1995, \A[482] );
  not g3592 (n_1997, \A[482] );
  and g3593 (n2804, \A[481] , n_1997);
  not g3594 (n_1999, n2804);
  and g3595 (n2805, \A[483] , n_1999);
  not g3596 (n_2000, n2803);
  and g3597 (n2806, n_2000, n2805);
  and g3598 (n2807, n_2000, n_1999);
  not g3599 (n_2001, \A[483] );
  not g3600 (n_2002, n2807);
  and g3601 (n2808, n_2001, n_2002);
  not g3602 (n_2003, n2806);
  not g3603 (n_2004, n2808);
  and g3604 (n2809, n_2003, n_2004);
  not g3605 (n_2006, \A[484] );
  and g3606 (n2810, n_2006, \A[485] );
  not g3607 (n_2008, \A[485] );
  and g3608 (n2811, \A[484] , n_2008);
  not g3609 (n_2010, n2811);
  and g3610 (n2812, \A[486] , n_2010);
  not g3611 (n_2011, n2810);
  and g3612 (n2813, n_2011, n2812);
  and g3613 (n2814, n_2011, n_2010);
  not g3614 (n_2012, \A[486] );
  not g3615 (n_2013, n2814);
  and g3616 (n2815, n_2012, n_2013);
  not g3617 (n_2014, n2813);
  not g3618 (n_2015, n2815);
  and g3619 (n2816, n_2014, n_2015);
  not g3620 (n_2016, n2809);
  and g3621 (n2817, n_2016, n2816);
  not g3622 (n_2017, n2816);
  and g3623 (n2818, n2809, n_2017);
  not g3624 (n_2018, n2817);
  not g3625 (n_2019, n2818);
  and g3626 (n2819, n_2018, n_2019);
  and g3627 (n2820, \A[484] , \A[485] );
  and g3628 (n2821, \A[486] , n_2013);
  not g3629 (n_2020, n2820);
  not g3630 (n_2021, n2821);
  and g3631 (n2822, n_2020, n_2021);
  and g3632 (n2823, \A[481] , \A[482] );
  and g3633 (n2824, \A[483] , n_2002);
  not g3634 (n_2022, n2823);
  not g3635 (n_2023, n2824);
  and g3636 (n2825, n_2022, n_2023);
  not g3637 (n_2024, n2822);
  and g3638 (n2826, n_2024, n2825);
  not g3639 (n_2025, n2825);
  and g3640 (n2827, n2822, n_2025);
  not g3641 (n_2026, n2826);
  not g3642 (n_2027, n2827);
  and g3643 (n2828, n_2026, n_2027);
  and g3644 (n2829, n_2016, n_2017);
  not g3645 (n_2028, n2828);
  and g3646 (n2830, n_2028, n2829);
  and g3647 (n2831, n_2024, n_2025);
  not g3648 (n_2029, n2830);
  not g3649 (n_2030, n2831);
  and g3650 (n2832, n_2029, n_2030);
  and g3651 (n2833, n_2026, n2829);
  and g3652 (n2834, n_2027, n2833);
  not g3653 (n_2031, n2829);
  and g3654 (n2835, n_2028, n_2031);
  not g3655 (n_2032, n2834);
  not g3656 (n_2033, n2835);
  and g3657 (n2836, n_2032, n_2033);
  not g3658 (n_2034, n2832);
  not g3659 (n_2035, n2836);
  and g3660 (n2837, n_2034, n_2035);
  not g3661 (n_2036, n2819);
  not g3662 (n_2037, n2837);
  and g3663 (n2838, n_2036, n_2037);
  not g3664 (n_2039, \A[475] );
  and g3665 (n2839, n_2039, \A[476] );
  not g3666 (n_2041, \A[476] );
  and g3667 (n2840, \A[475] , n_2041);
  not g3668 (n_2043, n2840);
  and g3669 (n2841, \A[477] , n_2043);
  not g3670 (n_2044, n2839);
  and g3671 (n2842, n_2044, n2841);
  and g3672 (n2843, n_2044, n_2043);
  not g3673 (n_2045, \A[477] );
  not g3674 (n_2046, n2843);
  and g3675 (n2844, n_2045, n_2046);
  not g3676 (n_2047, n2842);
  not g3677 (n_2048, n2844);
  and g3678 (n2845, n_2047, n_2048);
  not g3679 (n_2050, \A[478] );
  and g3680 (n2846, n_2050, \A[479] );
  not g3681 (n_2052, \A[479] );
  and g3682 (n2847, \A[478] , n_2052);
  not g3683 (n_2054, n2847);
  and g3684 (n2848, \A[480] , n_2054);
  not g3685 (n_2055, n2846);
  and g3686 (n2849, n_2055, n2848);
  and g3687 (n2850, n_2055, n_2054);
  not g3688 (n_2056, \A[480] );
  not g3689 (n_2057, n2850);
  and g3690 (n2851, n_2056, n_2057);
  not g3691 (n_2058, n2849);
  not g3692 (n_2059, n2851);
  and g3693 (n2852, n_2058, n_2059);
  not g3694 (n_2060, n2845);
  and g3695 (n2853, n_2060, n2852);
  not g3696 (n_2061, n2852);
  and g3697 (n2854, n2845, n_2061);
  not g3698 (n_2062, n2853);
  not g3699 (n_2063, n2854);
  and g3700 (n2855, n_2062, n_2063);
  and g3701 (n2856, \A[478] , \A[479] );
  and g3702 (n2857, \A[480] , n_2057);
  not g3703 (n_2064, n2856);
  not g3704 (n_2065, n2857);
  and g3705 (n2858, n_2064, n_2065);
  and g3706 (n2859, \A[475] , \A[476] );
  and g3707 (n2860, \A[477] , n_2046);
  not g3708 (n_2066, n2859);
  not g3709 (n_2067, n2860);
  and g3710 (n2861, n_2066, n_2067);
  not g3711 (n_2068, n2858);
  and g3712 (n2862, n_2068, n2861);
  not g3713 (n_2069, n2861);
  and g3714 (n2863, n2858, n_2069);
  not g3715 (n_2070, n2862);
  not g3716 (n_2071, n2863);
  and g3717 (n2864, n_2070, n_2071);
  and g3718 (n2865, n_2060, n_2061);
  not g3719 (n_2072, n2864);
  and g3720 (n2866, n_2072, n2865);
  and g3721 (n2867, n_2068, n_2069);
  not g3722 (n_2073, n2866);
  not g3723 (n_2074, n2867);
  and g3724 (n2868, n_2073, n_2074);
  and g3725 (n2869, n_2070, n2865);
  and g3726 (n2870, n_2071, n2869);
  not g3727 (n_2075, n2865);
  and g3728 (n2871, n_2072, n_2075);
  not g3729 (n_2076, n2870);
  not g3730 (n_2077, n2871);
  and g3731 (n2872, n_2076, n_2077);
  not g3732 (n_2078, n2868);
  not g3733 (n_2079, n2872);
  and g3734 (n2873, n_2078, n_2079);
  not g3735 (n_2080, n2855);
  not g3736 (n_2081, n2873);
  and g3737 (n2874, n_2080, n_2081);
  not g3738 (n_2082, n2838);
  and g3739 (n2875, n_2082, n2874);
  not g3740 (n_2083, n2874);
  and g3741 (n2876, n2838, n_2083);
  not g3742 (n_2084, n2875);
  not g3743 (n_2085, n2876);
  and g3744 (n2877, n_2084, n_2085);
  not g3745 (n_2086, n2802);
  and g3746 (n2878, n_2086, n2877);
  not g3747 (n_2087, n2877);
  and g3748 (n2879, n2802, n_2087);
  not g3749 (n_2088, n2878);
  not g3750 (n_2089, n2879);
  and g3751 (n2880, n_2088, n_2089);
  not g3752 (n_2091, \A[505] );
  and g3753 (n2881, n_2091, \A[506] );
  not g3754 (n_2093, \A[506] );
  and g3755 (n2882, \A[505] , n_2093);
  not g3756 (n_2095, n2882);
  and g3757 (n2883, \A[507] , n_2095);
  not g3758 (n_2096, n2881);
  and g3759 (n2884, n_2096, n2883);
  and g3760 (n2885, n_2096, n_2095);
  not g3761 (n_2097, \A[507] );
  not g3762 (n_2098, n2885);
  and g3763 (n2886, n_2097, n_2098);
  not g3764 (n_2099, n2884);
  not g3765 (n_2100, n2886);
  and g3766 (n2887, n_2099, n_2100);
  not g3767 (n_2102, \A[508] );
  and g3768 (n2888, n_2102, \A[509] );
  not g3769 (n_2104, \A[509] );
  and g3770 (n2889, \A[508] , n_2104);
  not g3771 (n_2106, n2889);
  and g3772 (n2890, \A[510] , n_2106);
  not g3773 (n_2107, n2888);
  and g3774 (n2891, n_2107, n2890);
  and g3775 (n2892, n_2107, n_2106);
  not g3776 (n_2108, \A[510] );
  not g3777 (n_2109, n2892);
  and g3778 (n2893, n_2108, n_2109);
  not g3779 (n_2110, n2891);
  not g3780 (n_2111, n2893);
  and g3781 (n2894, n_2110, n_2111);
  not g3782 (n_2112, n2887);
  and g3783 (n2895, n_2112, n2894);
  not g3784 (n_2113, n2894);
  and g3785 (n2896, n2887, n_2113);
  not g3786 (n_2114, n2895);
  not g3787 (n_2115, n2896);
  and g3788 (n2897, n_2114, n_2115);
  and g3789 (n2898, \A[508] , \A[509] );
  and g3790 (n2899, \A[510] , n_2109);
  not g3791 (n_2116, n2898);
  not g3792 (n_2117, n2899);
  and g3793 (n2900, n_2116, n_2117);
  and g3794 (n2901, \A[505] , \A[506] );
  and g3795 (n2902, \A[507] , n_2098);
  not g3796 (n_2118, n2901);
  not g3797 (n_2119, n2902);
  and g3798 (n2903, n_2118, n_2119);
  not g3799 (n_2120, n2900);
  and g3800 (n2904, n_2120, n2903);
  not g3801 (n_2121, n2903);
  and g3802 (n2905, n2900, n_2121);
  not g3803 (n_2122, n2904);
  not g3804 (n_2123, n2905);
  and g3805 (n2906, n_2122, n_2123);
  and g3806 (n2907, n_2112, n_2113);
  not g3807 (n_2124, n2906);
  and g3808 (n2908, n_2124, n2907);
  and g3809 (n2909, n_2120, n_2121);
  not g3810 (n_2125, n2908);
  not g3811 (n_2126, n2909);
  and g3812 (n2910, n_2125, n_2126);
  and g3813 (n2911, n_2122, n2907);
  and g3814 (n2912, n_2123, n2911);
  not g3815 (n_2127, n2907);
  and g3816 (n2913, n_2124, n_2127);
  not g3817 (n_2128, n2912);
  not g3818 (n_2129, n2913);
  and g3819 (n2914, n_2128, n_2129);
  not g3820 (n_2130, n2910);
  not g3821 (n_2131, n2914);
  and g3822 (n2915, n_2130, n_2131);
  not g3823 (n_2132, n2897);
  not g3824 (n_2133, n2915);
  and g3825 (n2916, n_2132, n_2133);
  not g3826 (n_2135, \A[499] );
  and g3827 (n2917, n_2135, \A[500] );
  not g3828 (n_2137, \A[500] );
  and g3829 (n2918, \A[499] , n_2137);
  not g3830 (n_2139, n2918);
  and g3831 (n2919, \A[501] , n_2139);
  not g3832 (n_2140, n2917);
  and g3833 (n2920, n_2140, n2919);
  and g3834 (n2921, n_2140, n_2139);
  not g3835 (n_2141, \A[501] );
  not g3836 (n_2142, n2921);
  and g3837 (n2922, n_2141, n_2142);
  not g3838 (n_2143, n2920);
  not g3839 (n_2144, n2922);
  and g3840 (n2923, n_2143, n_2144);
  not g3841 (n_2146, \A[502] );
  and g3842 (n2924, n_2146, \A[503] );
  not g3843 (n_2148, \A[503] );
  and g3844 (n2925, \A[502] , n_2148);
  not g3845 (n_2150, n2925);
  and g3846 (n2926, \A[504] , n_2150);
  not g3847 (n_2151, n2924);
  and g3848 (n2927, n_2151, n2926);
  and g3849 (n2928, n_2151, n_2150);
  not g3850 (n_2152, \A[504] );
  not g3851 (n_2153, n2928);
  and g3852 (n2929, n_2152, n_2153);
  not g3853 (n_2154, n2927);
  not g3854 (n_2155, n2929);
  and g3855 (n2930, n_2154, n_2155);
  not g3856 (n_2156, n2923);
  and g3857 (n2931, n_2156, n2930);
  not g3858 (n_2157, n2930);
  and g3859 (n2932, n2923, n_2157);
  not g3860 (n_2158, n2931);
  not g3861 (n_2159, n2932);
  and g3862 (n2933, n_2158, n_2159);
  and g3863 (n2934, \A[502] , \A[503] );
  and g3864 (n2935, \A[504] , n_2153);
  not g3865 (n_2160, n2934);
  not g3866 (n_2161, n2935);
  and g3867 (n2936, n_2160, n_2161);
  and g3868 (n2937, \A[499] , \A[500] );
  and g3869 (n2938, \A[501] , n_2142);
  not g3870 (n_2162, n2937);
  not g3871 (n_2163, n2938);
  and g3872 (n2939, n_2162, n_2163);
  not g3873 (n_2164, n2936);
  and g3874 (n2940, n_2164, n2939);
  not g3875 (n_2165, n2939);
  and g3876 (n2941, n2936, n_2165);
  not g3877 (n_2166, n2940);
  not g3878 (n_2167, n2941);
  and g3879 (n2942, n_2166, n_2167);
  and g3880 (n2943, n_2156, n_2157);
  not g3881 (n_2168, n2942);
  and g3882 (n2944, n_2168, n2943);
  and g3883 (n2945, n_2164, n_2165);
  not g3884 (n_2169, n2944);
  not g3885 (n_2170, n2945);
  and g3886 (n2946, n_2169, n_2170);
  and g3887 (n2947, n_2166, n2943);
  and g3888 (n2948, n_2167, n2947);
  not g3889 (n_2171, n2943);
  and g3890 (n2949, n_2168, n_2171);
  not g3891 (n_2172, n2948);
  not g3892 (n_2173, n2949);
  and g3893 (n2950, n_2172, n_2173);
  not g3894 (n_2174, n2946);
  not g3895 (n_2175, n2950);
  and g3896 (n2951, n_2174, n_2175);
  not g3897 (n_2176, n2933);
  not g3898 (n_2177, n2951);
  and g3899 (n2952, n_2176, n_2177);
  not g3900 (n_2178, n2916);
  and g3901 (n2953, n_2178, n2952);
  not g3902 (n_2179, n2952);
  and g3903 (n2954, n2916, n_2179);
  not g3904 (n_2180, n2953);
  not g3905 (n_2181, n2954);
  and g3906 (n2955, n_2180, n_2181);
  not g3907 (n_2183, \A[493] );
  and g3908 (n2956, n_2183, \A[494] );
  not g3909 (n_2185, \A[494] );
  and g3910 (n2957, \A[493] , n_2185);
  not g3911 (n_2187, n2957);
  and g3912 (n2958, \A[495] , n_2187);
  not g3913 (n_2188, n2956);
  and g3914 (n2959, n_2188, n2958);
  and g3915 (n2960, n_2188, n_2187);
  not g3916 (n_2189, \A[495] );
  not g3917 (n_2190, n2960);
  and g3918 (n2961, n_2189, n_2190);
  not g3919 (n_2191, n2959);
  not g3920 (n_2192, n2961);
  and g3921 (n2962, n_2191, n_2192);
  not g3922 (n_2194, \A[496] );
  and g3923 (n2963, n_2194, \A[497] );
  not g3924 (n_2196, \A[497] );
  and g3925 (n2964, \A[496] , n_2196);
  not g3926 (n_2198, n2964);
  and g3927 (n2965, \A[498] , n_2198);
  not g3928 (n_2199, n2963);
  and g3929 (n2966, n_2199, n2965);
  and g3930 (n2967, n_2199, n_2198);
  not g3931 (n_2200, \A[498] );
  not g3932 (n_2201, n2967);
  and g3933 (n2968, n_2200, n_2201);
  not g3934 (n_2202, n2966);
  not g3935 (n_2203, n2968);
  and g3936 (n2969, n_2202, n_2203);
  not g3937 (n_2204, n2962);
  and g3938 (n2970, n_2204, n2969);
  not g3939 (n_2205, n2969);
  and g3940 (n2971, n2962, n_2205);
  not g3941 (n_2206, n2970);
  not g3942 (n_2207, n2971);
  and g3943 (n2972, n_2206, n_2207);
  and g3944 (n2973, \A[496] , \A[497] );
  and g3945 (n2974, \A[498] , n_2201);
  not g3946 (n_2208, n2973);
  not g3947 (n_2209, n2974);
  and g3948 (n2975, n_2208, n_2209);
  and g3949 (n2976, \A[493] , \A[494] );
  and g3950 (n2977, \A[495] , n_2190);
  not g3951 (n_2210, n2976);
  not g3952 (n_2211, n2977);
  and g3953 (n2978, n_2210, n_2211);
  not g3954 (n_2212, n2975);
  and g3955 (n2979, n_2212, n2978);
  not g3956 (n_2213, n2978);
  and g3957 (n2980, n2975, n_2213);
  not g3958 (n_2214, n2979);
  not g3959 (n_2215, n2980);
  and g3960 (n2981, n_2214, n_2215);
  and g3961 (n2982, n_2204, n_2205);
  not g3962 (n_2216, n2981);
  and g3963 (n2983, n_2216, n2982);
  and g3964 (n2984, n_2212, n_2213);
  not g3965 (n_2217, n2983);
  not g3966 (n_2218, n2984);
  and g3967 (n2985, n_2217, n_2218);
  and g3968 (n2986, n_2214, n2982);
  and g3969 (n2987, n_2215, n2986);
  not g3970 (n_2219, n2982);
  and g3971 (n2988, n_2216, n_2219);
  not g3972 (n_2220, n2987);
  not g3973 (n_2221, n2988);
  and g3974 (n2989, n_2220, n_2221);
  not g3975 (n_2222, n2985);
  not g3976 (n_2223, n2989);
  and g3977 (n2990, n_2222, n_2223);
  not g3978 (n_2224, n2972);
  not g3979 (n_2225, n2990);
  and g3980 (n2991, n_2224, n_2225);
  not g3981 (n_2227, \A[487] );
  and g3982 (n2992, n_2227, \A[488] );
  not g3983 (n_2229, \A[488] );
  and g3984 (n2993, \A[487] , n_2229);
  not g3985 (n_2231, n2993);
  and g3986 (n2994, \A[489] , n_2231);
  not g3987 (n_2232, n2992);
  and g3988 (n2995, n_2232, n2994);
  and g3989 (n2996, n_2232, n_2231);
  not g3990 (n_2233, \A[489] );
  not g3991 (n_2234, n2996);
  and g3992 (n2997, n_2233, n_2234);
  not g3993 (n_2235, n2995);
  not g3994 (n_2236, n2997);
  and g3995 (n2998, n_2235, n_2236);
  not g3996 (n_2238, \A[490] );
  and g3997 (n2999, n_2238, \A[491] );
  not g3998 (n_2240, \A[491] );
  and g3999 (n3000, \A[490] , n_2240);
  not g4000 (n_2242, n3000);
  and g4001 (n3001, \A[492] , n_2242);
  not g4002 (n_2243, n2999);
  and g4003 (n3002, n_2243, n3001);
  and g4004 (n3003, n_2243, n_2242);
  not g4005 (n_2244, \A[492] );
  not g4006 (n_2245, n3003);
  and g4007 (n3004, n_2244, n_2245);
  not g4008 (n_2246, n3002);
  not g4009 (n_2247, n3004);
  and g4010 (n3005, n_2246, n_2247);
  not g4011 (n_2248, n2998);
  and g4012 (n3006, n_2248, n3005);
  not g4013 (n_2249, n3005);
  and g4014 (n3007, n2998, n_2249);
  not g4015 (n_2250, n3006);
  not g4016 (n_2251, n3007);
  and g4017 (n3008, n_2250, n_2251);
  and g4018 (n3009, \A[490] , \A[491] );
  and g4019 (n3010, \A[492] , n_2245);
  not g4020 (n_2252, n3009);
  not g4021 (n_2253, n3010);
  and g4022 (n3011, n_2252, n_2253);
  and g4023 (n3012, \A[487] , \A[488] );
  and g4024 (n3013, \A[489] , n_2234);
  not g4025 (n_2254, n3012);
  not g4026 (n_2255, n3013);
  and g4027 (n3014, n_2254, n_2255);
  not g4028 (n_2256, n3011);
  and g4029 (n3015, n_2256, n3014);
  not g4030 (n_2257, n3014);
  and g4031 (n3016, n3011, n_2257);
  not g4032 (n_2258, n3015);
  not g4033 (n_2259, n3016);
  and g4034 (n3017, n_2258, n_2259);
  and g4035 (n3018, n_2248, n_2249);
  not g4036 (n_2260, n3017);
  and g4037 (n3019, n_2260, n3018);
  and g4038 (n3020, n_2256, n_2257);
  not g4039 (n_2261, n3019);
  not g4040 (n_2262, n3020);
  and g4041 (n3021, n_2261, n_2262);
  and g4042 (n3022, n_2258, n3018);
  and g4043 (n3023, n_2259, n3022);
  not g4044 (n_2263, n3018);
  and g4045 (n3024, n_2260, n_2263);
  not g4046 (n_2264, n3023);
  not g4047 (n_2265, n3024);
  and g4048 (n3025, n_2264, n_2265);
  not g4049 (n_2266, n3021);
  not g4050 (n_2267, n3025);
  and g4051 (n3026, n_2266, n_2267);
  not g4052 (n_2268, n3008);
  not g4053 (n_2269, n3026);
  and g4054 (n3027, n_2268, n_2269);
  not g4055 (n_2270, n2991);
  and g4056 (n3028, n_2270, n3027);
  not g4057 (n_2271, n3027);
  and g4058 (n3029, n2991, n_2271);
  not g4059 (n_2272, n3028);
  not g4060 (n_2273, n3029);
  and g4061 (n3030, n_2272, n_2273);
  not g4062 (n_2274, n2955);
  and g4063 (n3031, n_2274, n3030);
  not g4064 (n_2275, n3030);
  and g4065 (n3032, n2955, n_2275);
  not g4066 (n_2276, n3031);
  not g4067 (n_2277, n3032);
  and g4068 (n3033, n_2276, n_2277);
  not g4069 (n_2278, n2880);
  and g4070 (n3034, n_2278, n3033);
  not g4071 (n_2279, n3033);
  and g4072 (n3035, n2880, n_2279);
  not g4073 (n_2280, n3034);
  not g4074 (n_2281, n3035);
  and g4075 (n3036, n_2280, n_2281);
  not g4076 (n_2283, \A[553] );
  and g4077 (n3037, n_2283, \A[554] );
  not g4078 (n_2285, \A[554] );
  and g4079 (n3038, \A[553] , n_2285);
  not g4080 (n_2287, n3038);
  and g4081 (n3039, \A[555] , n_2287);
  not g4082 (n_2288, n3037);
  and g4083 (n3040, n_2288, n3039);
  and g4084 (n3041, n_2288, n_2287);
  not g4085 (n_2289, \A[555] );
  not g4086 (n_2290, n3041);
  and g4087 (n3042, n_2289, n_2290);
  not g4088 (n_2291, n3040);
  not g4089 (n_2292, n3042);
  and g4090 (n3043, n_2291, n_2292);
  not g4091 (n_2294, \A[556] );
  and g4092 (n3044, n_2294, \A[557] );
  not g4093 (n_2296, \A[557] );
  and g4094 (n3045, \A[556] , n_2296);
  not g4095 (n_2298, n3045);
  and g4096 (n3046, \A[558] , n_2298);
  not g4097 (n_2299, n3044);
  and g4098 (n3047, n_2299, n3046);
  and g4099 (n3048, n_2299, n_2298);
  not g4100 (n_2300, \A[558] );
  not g4101 (n_2301, n3048);
  and g4102 (n3049, n_2300, n_2301);
  not g4103 (n_2302, n3047);
  not g4104 (n_2303, n3049);
  and g4105 (n3050, n_2302, n_2303);
  not g4106 (n_2304, n3043);
  and g4107 (n3051, n_2304, n3050);
  not g4108 (n_2305, n3050);
  and g4109 (n3052, n3043, n_2305);
  not g4110 (n_2306, n3051);
  not g4111 (n_2307, n3052);
  and g4112 (n3053, n_2306, n_2307);
  and g4113 (n3054, \A[556] , \A[557] );
  and g4114 (n3055, \A[558] , n_2301);
  not g4115 (n_2308, n3054);
  not g4116 (n_2309, n3055);
  and g4117 (n3056, n_2308, n_2309);
  and g4118 (n3057, \A[553] , \A[554] );
  and g4119 (n3058, \A[555] , n_2290);
  not g4120 (n_2310, n3057);
  not g4121 (n_2311, n3058);
  and g4122 (n3059, n_2310, n_2311);
  not g4123 (n_2312, n3056);
  and g4124 (n3060, n_2312, n3059);
  not g4125 (n_2313, n3059);
  and g4126 (n3061, n3056, n_2313);
  not g4127 (n_2314, n3060);
  not g4128 (n_2315, n3061);
  and g4129 (n3062, n_2314, n_2315);
  and g4130 (n3063, n_2304, n_2305);
  not g4131 (n_2316, n3062);
  and g4132 (n3064, n_2316, n3063);
  and g4133 (n3065, n_2312, n_2313);
  not g4134 (n_2317, n3064);
  not g4135 (n_2318, n3065);
  and g4136 (n3066, n_2317, n_2318);
  and g4137 (n3067, n_2314, n3063);
  and g4138 (n3068, n_2315, n3067);
  not g4139 (n_2319, n3063);
  and g4140 (n3069, n_2316, n_2319);
  not g4141 (n_2320, n3068);
  not g4142 (n_2321, n3069);
  and g4143 (n3070, n_2320, n_2321);
  not g4144 (n_2322, n3066);
  not g4145 (n_2323, n3070);
  and g4146 (n3071, n_2322, n_2323);
  not g4147 (n_2324, n3053);
  not g4148 (n_2325, n3071);
  and g4149 (n3072, n_2324, n_2325);
  not g4150 (n_2327, \A[547] );
  and g4151 (n3073, n_2327, \A[548] );
  not g4152 (n_2329, \A[548] );
  and g4153 (n3074, \A[547] , n_2329);
  not g4154 (n_2331, n3074);
  and g4155 (n3075, \A[549] , n_2331);
  not g4156 (n_2332, n3073);
  and g4157 (n3076, n_2332, n3075);
  and g4158 (n3077, n_2332, n_2331);
  not g4159 (n_2333, \A[549] );
  not g4160 (n_2334, n3077);
  and g4161 (n3078, n_2333, n_2334);
  not g4162 (n_2335, n3076);
  not g4163 (n_2336, n3078);
  and g4164 (n3079, n_2335, n_2336);
  not g4165 (n_2338, \A[550] );
  and g4166 (n3080, n_2338, \A[551] );
  not g4167 (n_2340, \A[551] );
  and g4168 (n3081, \A[550] , n_2340);
  not g4169 (n_2342, n3081);
  and g4170 (n3082, \A[552] , n_2342);
  not g4171 (n_2343, n3080);
  and g4172 (n3083, n_2343, n3082);
  and g4173 (n3084, n_2343, n_2342);
  not g4174 (n_2344, \A[552] );
  not g4175 (n_2345, n3084);
  and g4176 (n3085, n_2344, n_2345);
  not g4177 (n_2346, n3083);
  not g4178 (n_2347, n3085);
  and g4179 (n3086, n_2346, n_2347);
  not g4180 (n_2348, n3079);
  and g4181 (n3087, n_2348, n3086);
  not g4182 (n_2349, n3086);
  and g4183 (n3088, n3079, n_2349);
  not g4184 (n_2350, n3087);
  not g4185 (n_2351, n3088);
  and g4186 (n3089, n_2350, n_2351);
  and g4187 (n3090, \A[550] , \A[551] );
  and g4188 (n3091, \A[552] , n_2345);
  not g4189 (n_2352, n3090);
  not g4190 (n_2353, n3091);
  and g4191 (n3092, n_2352, n_2353);
  and g4192 (n3093, \A[547] , \A[548] );
  and g4193 (n3094, \A[549] , n_2334);
  not g4194 (n_2354, n3093);
  not g4195 (n_2355, n3094);
  and g4196 (n3095, n_2354, n_2355);
  not g4197 (n_2356, n3092);
  and g4198 (n3096, n_2356, n3095);
  not g4199 (n_2357, n3095);
  and g4200 (n3097, n3092, n_2357);
  not g4201 (n_2358, n3096);
  not g4202 (n_2359, n3097);
  and g4203 (n3098, n_2358, n_2359);
  and g4204 (n3099, n_2348, n_2349);
  not g4205 (n_2360, n3098);
  and g4206 (n3100, n_2360, n3099);
  and g4207 (n3101, n_2356, n_2357);
  not g4208 (n_2361, n3100);
  not g4209 (n_2362, n3101);
  and g4210 (n3102, n_2361, n_2362);
  and g4211 (n3103, n_2358, n3099);
  and g4212 (n3104, n_2359, n3103);
  not g4213 (n_2363, n3099);
  and g4214 (n3105, n_2360, n_2363);
  not g4215 (n_2364, n3104);
  not g4216 (n_2365, n3105);
  and g4217 (n3106, n_2364, n_2365);
  not g4218 (n_2366, n3102);
  not g4219 (n_2367, n3106);
  and g4220 (n3107, n_2366, n_2367);
  not g4221 (n_2368, n3089);
  not g4222 (n_2369, n3107);
  and g4223 (n3108, n_2368, n_2369);
  not g4224 (n_2370, n3072);
  and g4225 (n3109, n_2370, n3108);
  not g4226 (n_2371, n3108);
  and g4227 (n3110, n3072, n_2371);
  not g4228 (n_2372, n3109);
  not g4229 (n_2373, n3110);
  and g4230 (n3111, n_2372, n_2373);
  not g4231 (n_2375, \A[541] );
  and g4232 (n3112, n_2375, \A[542] );
  not g4233 (n_2377, \A[542] );
  and g4234 (n3113, \A[541] , n_2377);
  not g4235 (n_2379, n3113);
  and g4236 (n3114, \A[543] , n_2379);
  not g4237 (n_2380, n3112);
  and g4238 (n3115, n_2380, n3114);
  and g4239 (n3116, n_2380, n_2379);
  not g4240 (n_2381, \A[543] );
  not g4241 (n_2382, n3116);
  and g4242 (n3117, n_2381, n_2382);
  not g4243 (n_2383, n3115);
  not g4244 (n_2384, n3117);
  and g4245 (n3118, n_2383, n_2384);
  not g4246 (n_2386, \A[544] );
  and g4247 (n3119, n_2386, \A[545] );
  not g4248 (n_2388, \A[545] );
  and g4249 (n3120, \A[544] , n_2388);
  not g4250 (n_2390, n3120);
  and g4251 (n3121, \A[546] , n_2390);
  not g4252 (n_2391, n3119);
  and g4253 (n3122, n_2391, n3121);
  and g4254 (n3123, n_2391, n_2390);
  not g4255 (n_2392, \A[546] );
  not g4256 (n_2393, n3123);
  and g4257 (n3124, n_2392, n_2393);
  not g4258 (n_2394, n3122);
  not g4259 (n_2395, n3124);
  and g4260 (n3125, n_2394, n_2395);
  not g4261 (n_2396, n3118);
  and g4262 (n3126, n_2396, n3125);
  not g4263 (n_2397, n3125);
  and g4264 (n3127, n3118, n_2397);
  not g4265 (n_2398, n3126);
  not g4266 (n_2399, n3127);
  and g4267 (n3128, n_2398, n_2399);
  and g4268 (n3129, \A[544] , \A[545] );
  and g4269 (n3130, \A[546] , n_2393);
  not g4270 (n_2400, n3129);
  not g4271 (n_2401, n3130);
  and g4272 (n3131, n_2400, n_2401);
  and g4273 (n3132, \A[541] , \A[542] );
  and g4274 (n3133, \A[543] , n_2382);
  not g4275 (n_2402, n3132);
  not g4276 (n_2403, n3133);
  and g4277 (n3134, n_2402, n_2403);
  not g4278 (n_2404, n3131);
  and g4279 (n3135, n_2404, n3134);
  not g4280 (n_2405, n3134);
  and g4281 (n3136, n3131, n_2405);
  not g4282 (n_2406, n3135);
  not g4283 (n_2407, n3136);
  and g4284 (n3137, n_2406, n_2407);
  and g4285 (n3138, n_2396, n_2397);
  not g4286 (n_2408, n3137);
  and g4287 (n3139, n_2408, n3138);
  and g4288 (n3140, n_2404, n_2405);
  not g4289 (n_2409, n3139);
  not g4290 (n_2410, n3140);
  and g4291 (n3141, n_2409, n_2410);
  and g4292 (n3142, n_2406, n3138);
  and g4293 (n3143, n_2407, n3142);
  not g4294 (n_2411, n3138);
  and g4295 (n3144, n_2408, n_2411);
  not g4296 (n_2412, n3143);
  not g4297 (n_2413, n3144);
  and g4298 (n3145, n_2412, n_2413);
  not g4299 (n_2414, n3141);
  not g4300 (n_2415, n3145);
  and g4301 (n3146, n_2414, n_2415);
  not g4302 (n_2416, n3128);
  not g4303 (n_2417, n3146);
  and g4304 (n3147, n_2416, n_2417);
  not g4305 (n_2419, \A[535] );
  and g4306 (n3148, n_2419, \A[536] );
  not g4307 (n_2421, \A[536] );
  and g4308 (n3149, \A[535] , n_2421);
  not g4309 (n_2423, n3149);
  and g4310 (n3150, \A[537] , n_2423);
  not g4311 (n_2424, n3148);
  and g4312 (n3151, n_2424, n3150);
  and g4313 (n3152, n_2424, n_2423);
  not g4314 (n_2425, \A[537] );
  not g4315 (n_2426, n3152);
  and g4316 (n3153, n_2425, n_2426);
  not g4317 (n_2427, n3151);
  not g4318 (n_2428, n3153);
  and g4319 (n3154, n_2427, n_2428);
  not g4320 (n_2430, \A[538] );
  and g4321 (n3155, n_2430, \A[539] );
  not g4322 (n_2432, \A[539] );
  and g4323 (n3156, \A[538] , n_2432);
  not g4324 (n_2434, n3156);
  and g4325 (n3157, \A[540] , n_2434);
  not g4326 (n_2435, n3155);
  and g4327 (n3158, n_2435, n3157);
  and g4328 (n3159, n_2435, n_2434);
  not g4329 (n_2436, \A[540] );
  not g4330 (n_2437, n3159);
  and g4331 (n3160, n_2436, n_2437);
  not g4332 (n_2438, n3158);
  not g4333 (n_2439, n3160);
  and g4334 (n3161, n_2438, n_2439);
  not g4335 (n_2440, n3154);
  and g4336 (n3162, n_2440, n3161);
  not g4337 (n_2441, n3161);
  and g4338 (n3163, n3154, n_2441);
  not g4339 (n_2442, n3162);
  not g4340 (n_2443, n3163);
  and g4341 (n3164, n_2442, n_2443);
  and g4342 (n3165, \A[538] , \A[539] );
  and g4343 (n3166, \A[540] , n_2437);
  not g4344 (n_2444, n3165);
  not g4345 (n_2445, n3166);
  and g4346 (n3167, n_2444, n_2445);
  and g4347 (n3168, \A[535] , \A[536] );
  and g4348 (n3169, \A[537] , n_2426);
  not g4349 (n_2446, n3168);
  not g4350 (n_2447, n3169);
  and g4351 (n3170, n_2446, n_2447);
  not g4352 (n_2448, n3167);
  and g4353 (n3171, n_2448, n3170);
  not g4354 (n_2449, n3170);
  and g4355 (n3172, n3167, n_2449);
  not g4356 (n_2450, n3171);
  not g4357 (n_2451, n3172);
  and g4358 (n3173, n_2450, n_2451);
  and g4359 (n3174, n_2440, n_2441);
  not g4360 (n_2452, n3173);
  and g4361 (n3175, n_2452, n3174);
  and g4362 (n3176, n_2448, n_2449);
  not g4363 (n_2453, n3175);
  not g4364 (n_2454, n3176);
  and g4365 (n3177, n_2453, n_2454);
  and g4366 (n3178, n_2450, n3174);
  and g4367 (n3179, n_2451, n3178);
  not g4368 (n_2455, n3174);
  and g4369 (n3180, n_2452, n_2455);
  not g4370 (n_2456, n3179);
  not g4371 (n_2457, n3180);
  and g4372 (n3181, n_2456, n_2457);
  not g4373 (n_2458, n3177);
  not g4374 (n_2459, n3181);
  and g4375 (n3182, n_2458, n_2459);
  not g4376 (n_2460, n3164);
  not g4377 (n_2461, n3182);
  and g4378 (n3183, n_2460, n_2461);
  not g4379 (n_2462, n3147);
  and g4380 (n3184, n_2462, n3183);
  not g4381 (n_2463, n3183);
  and g4382 (n3185, n3147, n_2463);
  not g4383 (n_2464, n3184);
  not g4384 (n_2465, n3185);
  and g4385 (n3186, n_2464, n_2465);
  not g4386 (n_2466, n3111);
  and g4387 (n3187, n_2466, n3186);
  not g4388 (n_2467, n3186);
  and g4389 (n3188, n3111, n_2467);
  not g4390 (n_2468, n3187);
  not g4391 (n_2469, n3188);
  and g4392 (n3189, n_2468, n_2469);
  not g4393 (n_2471, \A[529] );
  and g4394 (n3190, n_2471, \A[530] );
  not g4395 (n_2473, \A[530] );
  and g4396 (n3191, \A[529] , n_2473);
  not g4397 (n_2475, n3191);
  and g4398 (n3192, \A[531] , n_2475);
  not g4399 (n_2476, n3190);
  and g4400 (n3193, n_2476, n3192);
  and g4401 (n3194, n_2476, n_2475);
  not g4402 (n_2477, \A[531] );
  not g4403 (n_2478, n3194);
  and g4404 (n3195, n_2477, n_2478);
  not g4405 (n_2479, n3193);
  not g4406 (n_2480, n3195);
  and g4407 (n3196, n_2479, n_2480);
  not g4408 (n_2482, \A[532] );
  and g4409 (n3197, n_2482, \A[533] );
  not g4410 (n_2484, \A[533] );
  and g4411 (n3198, \A[532] , n_2484);
  not g4412 (n_2486, n3198);
  and g4413 (n3199, \A[534] , n_2486);
  not g4414 (n_2487, n3197);
  and g4415 (n3200, n_2487, n3199);
  and g4416 (n3201, n_2487, n_2486);
  not g4417 (n_2488, \A[534] );
  not g4418 (n_2489, n3201);
  and g4419 (n3202, n_2488, n_2489);
  not g4420 (n_2490, n3200);
  not g4421 (n_2491, n3202);
  and g4422 (n3203, n_2490, n_2491);
  not g4423 (n_2492, n3196);
  and g4424 (n3204, n_2492, n3203);
  not g4425 (n_2493, n3203);
  and g4426 (n3205, n3196, n_2493);
  not g4427 (n_2494, n3204);
  not g4428 (n_2495, n3205);
  and g4429 (n3206, n_2494, n_2495);
  and g4430 (n3207, \A[532] , \A[533] );
  and g4431 (n3208, \A[534] , n_2489);
  not g4432 (n_2496, n3207);
  not g4433 (n_2497, n3208);
  and g4434 (n3209, n_2496, n_2497);
  and g4435 (n3210, \A[529] , \A[530] );
  and g4436 (n3211, \A[531] , n_2478);
  not g4437 (n_2498, n3210);
  not g4438 (n_2499, n3211);
  and g4439 (n3212, n_2498, n_2499);
  not g4440 (n_2500, n3209);
  and g4441 (n3213, n_2500, n3212);
  not g4442 (n_2501, n3212);
  and g4443 (n3214, n3209, n_2501);
  not g4444 (n_2502, n3213);
  not g4445 (n_2503, n3214);
  and g4446 (n3215, n_2502, n_2503);
  and g4447 (n3216, n_2492, n_2493);
  not g4448 (n_2504, n3215);
  and g4449 (n3217, n_2504, n3216);
  and g4450 (n3218, n_2500, n_2501);
  not g4451 (n_2505, n3217);
  not g4452 (n_2506, n3218);
  and g4453 (n3219, n_2505, n_2506);
  and g4454 (n3220, n_2502, n3216);
  and g4455 (n3221, n_2503, n3220);
  not g4456 (n_2507, n3216);
  and g4457 (n3222, n_2504, n_2507);
  not g4458 (n_2508, n3221);
  not g4459 (n_2509, n3222);
  and g4460 (n3223, n_2508, n_2509);
  not g4461 (n_2510, n3219);
  not g4462 (n_2511, n3223);
  and g4463 (n3224, n_2510, n_2511);
  not g4464 (n_2512, n3206);
  not g4465 (n_2513, n3224);
  and g4466 (n3225, n_2512, n_2513);
  not g4467 (n_2515, \A[523] );
  and g4468 (n3226, n_2515, \A[524] );
  not g4469 (n_2517, \A[524] );
  and g4470 (n3227, \A[523] , n_2517);
  not g4471 (n_2519, n3227);
  and g4472 (n3228, \A[525] , n_2519);
  not g4473 (n_2520, n3226);
  and g4474 (n3229, n_2520, n3228);
  and g4475 (n3230, n_2520, n_2519);
  not g4476 (n_2521, \A[525] );
  not g4477 (n_2522, n3230);
  and g4478 (n3231, n_2521, n_2522);
  not g4479 (n_2523, n3229);
  not g4480 (n_2524, n3231);
  and g4481 (n3232, n_2523, n_2524);
  not g4482 (n_2526, \A[526] );
  and g4483 (n3233, n_2526, \A[527] );
  not g4484 (n_2528, \A[527] );
  and g4485 (n3234, \A[526] , n_2528);
  not g4486 (n_2530, n3234);
  and g4487 (n3235, \A[528] , n_2530);
  not g4488 (n_2531, n3233);
  and g4489 (n3236, n_2531, n3235);
  and g4490 (n3237, n_2531, n_2530);
  not g4491 (n_2532, \A[528] );
  not g4492 (n_2533, n3237);
  and g4493 (n3238, n_2532, n_2533);
  not g4494 (n_2534, n3236);
  not g4495 (n_2535, n3238);
  and g4496 (n3239, n_2534, n_2535);
  not g4497 (n_2536, n3232);
  and g4498 (n3240, n_2536, n3239);
  not g4499 (n_2537, n3239);
  and g4500 (n3241, n3232, n_2537);
  not g4501 (n_2538, n3240);
  not g4502 (n_2539, n3241);
  and g4503 (n3242, n_2538, n_2539);
  and g4504 (n3243, \A[526] , \A[527] );
  and g4505 (n3244, \A[528] , n_2533);
  not g4506 (n_2540, n3243);
  not g4507 (n_2541, n3244);
  and g4508 (n3245, n_2540, n_2541);
  and g4509 (n3246, \A[523] , \A[524] );
  and g4510 (n3247, \A[525] , n_2522);
  not g4511 (n_2542, n3246);
  not g4512 (n_2543, n3247);
  and g4513 (n3248, n_2542, n_2543);
  not g4514 (n_2544, n3245);
  and g4515 (n3249, n_2544, n3248);
  not g4516 (n_2545, n3248);
  and g4517 (n3250, n3245, n_2545);
  not g4518 (n_2546, n3249);
  not g4519 (n_2547, n3250);
  and g4520 (n3251, n_2546, n_2547);
  and g4521 (n3252, n_2536, n_2537);
  not g4522 (n_2548, n3251);
  and g4523 (n3253, n_2548, n3252);
  and g4524 (n3254, n_2544, n_2545);
  not g4525 (n_2549, n3253);
  not g4526 (n_2550, n3254);
  and g4527 (n3255, n_2549, n_2550);
  and g4528 (n3256, n_2546, n3252);
  and g4529 (n3257, n_2547, n3256);
  not g4530 (n_2551, n3252);
  and g4531 (n3258, n_2548, n_2551);
  not g4532 (n_2552, n3257);
  not g4533 (n_2553, n3258);
  and g4534 (n3259, n_2552, n_2553);
  not g4535 (n_2554, n3255);
  not g4536 (n_2555, n3259);
  and g4537 (n3260, n_2554, n_2555);
  not g4538 (n_2556, n3242);
  not g4539 (n_2557, n3260);
  and g4540 (n3261, n_2556, n_2557);
  not g4541 (n_2558, n3225);
  and g4542 (n3262, n_2558, n3261);
  not g4543 (n_2559, n3261);
  and g4544 (n3263, n3225, n_2559);
  not g4545 (n_2560, n3262);
  not g4546 (n_2561, n3263);
  and g4547 (n3264, n_2560, n_2561);
  not g4548 (n_2563, \A[517] );
  and g4549 (n3265, n_2563, \A[518] );
  not g4550 (n_2565, \A[518] );
  and g4551 (n3266, \A[517] , n_2565);
  not g4552 (n_2567, n3266);
  and g4553 (n3267, \A[519] , n_2567);
  not g4554 (n_2568, n3265);
  and g4555 (n3268, n_2568, n3267);
  and g4556 (n3269, n_2568, n_2567);
  not g4557 (n_2569, \A[519] );
  not g4558 (n_2570, n3269);
  and g4559 (n3270, n_2569, n_2570);
  not g4560 (n_2571, n3268);
  not g4561 (n_2572, n3270);
  and g4562 (n3271, n_2571, n_2572);
  not g4563 (n_2574, \A[520] );
  and g4564 (n3272, n_2574, \A[521] );
  not g4565 (n_2576, \A[521] );
  and g4566 (n3273, \A[520] , n_2576);
  not g4567 (n_2578, n3273);
  and g4568 (n3274, \A[522] , n_2578);
  not g4569 (n_2579, n3272);
  and g4570 (n3275, n_2579, n3274);
  and g4571 (n3276, n_2579, n_2578);
  not g4572 (n_2580, \A[522] );
  not g4573 (n_2581, n3276);
  and g4574 (n3277, n_2580, n_2581);
  not g4575 (n_2582, n3275);
  not g4576 (n_2583, n3277);
  and g4577 (n3278, n_2582, n_2583);
  not g4578 (n_2584, n3271);
  and g4579 (n3279, n_2584, n3278);
  not g4580 (n_2585, n3278);
  and g4581 (n3280, n3271, n_2585);
  not g4582 (n_2586, n3279);
  not g4583 (n_2587, n3280);
  and g4584 (n3281, n_2586, n_2587);
  and g4585 (n3282, \A[520] , \A[521] );
  and g4586 (n3283, \A[522] , n_2581);
  not g4587 (n_2588, n3282);
  not g4588 (n_2589, n3283);
  and g4589 (n3284, n_2588, n_2589);
  and g4590 (n3285, \A[517] , \A[518] );
  and g4591 (n3286, \A[519] , n_2570);
  not g4592 (n_2590, n3285);
  not g4593 (n_2591, n3286);
  and g4594 (n3287, n_2590, n_2591);
  not g4595 (n_2592, n3284);
  and g4596 (n3288, n_2592, n3287);
  not g4597 (n_2593, n3287);
  and g4598 (n3289, n3284, n_2593);
  not g4599 (n_2594, n3288);
  not g4600 (n_2595, n3289);
  and g4601 (n3290, n_2594, n_2595);
  and g4602 (n3291, n_2584, n_2585);
  not g4603 (n_2596, n3290);
  and g4604 (n3292, n_2596, n3291);
  and g4605 (n3293, n_2592, n_2593);
  not g4606 (n_2597, n3292);
  not g4607 (n_2598, n3293);
  and g4608 (n3294, n_2597, n_2598);
  and g4609 (n3295, n_2594, n3291);
  and g4610 (n3296, n_2595, n3295);
  not g4611 (n_2599, n3291);
  and g4612 (n3297, n_2596, n_2599);
  not g4613 (n_2600, n3296);
  not g4614 (n_2601, n3297);
  and g4615 (n3298, n_2600, n_2601);
  not g4616 (n_2602, n3294);
  not g4617 (n_2603, n3298);
  and g4618 (n3299, n_2602, n_2603);
  not g4619 (n_2604, n3281);
  not g4620 (n_2605, n3299);
  and g4621 (n3300, n_2604, n_2605);
  not g4622 (n_2607, \A[511] );
  and g4623 (n3301, n_2607, \A[512] );
  not g4624 (n_2609, \A[512] );
  and g4625 (n3302, \A[511] , n_2609);
  not g4626 (n_2611, n3302);
  and g4627 (n3303, \A[513] , n_2611);
  not g4628 (n_2612, n3301);
  and g4629 (n3304, n_2612, n3303);
  and g4630 (n3305, n_2612, n_2611);
  not g4631 (n_2613, \A[513] );
  not g4632 (n_2614, n3305);
  and g4633 (n3306, n_2613, n_2614);
  not g4634 (n_2615, n3304);
  not g4635 (n_2616, n3306);
  and g4636 (n3307, n_2615, n_2616);
  not g4637 (n_2618, \A[514] );
  and g4638 (n3308, n_2618, \A[515] );
  not g4639 (n_2620, \A[515] );
  and g4640 (n3309, \A[514] , n_2620);
  not g4641 (n_2622, n3309);
  and g4642 (n3310, \A[516] , n_2622);
  not g4643 (n_2623, n3308);
  and g4644 (n3311, n_2623, n3310);
  and g4645 (n3312, n_2623, n_2622);
  not g4646 (n_2624, \A[516] );
  not g4647 (n_2625, n3312);
  and g4648 (n3313, n_2624, n_2625);
  not g4649 (n_2626, n3311);
  not g4650 (n_2627, n3313);
  and g4651 (n3314, n_2626, n_2627);
  not g4652 (n_2628, n3307);
  and g4653 (n3315, n_2628, n3314);
  not g4654 (n_2629, n3314);
  and g4655 (n3316, n3307, n_2629);
  not g4656 (n_2630, n3315);
  not g4657 (n_2631, n3316);
  and g4658 (n3317, n_2630, n_2631);
  and g4659 (n3318, \A[514] , \A[515] );
  and g4660 (n3319, \A[516] , n_2625);
  not g4661 (n_2632, n3318);
  not g4662 (n_2633, n3319);
  and g4663 (n3320, n_2632, n_2633);
  and g4664 (n3321, \A[511] , \A[512] );
  and g4665 (n3322, \A[513] , n_2614);
  not g4666 (n_2634, n3321);
  not g4667 (n_2635, n3322);
  and g4668 (n3323, n_2634, n_2635);
  not g4669 (n_2636, n3320);
  and g4670 (n3324, n_2636, n3323);
  not g4671 (n_2637, n3323);
  and g4672 (n3325, n3320, n_2637);
  not g4673 (n_2638, n3324);
  not g4674 (n_2639, n3325);
  and g4675 (n3326, n_2638, n_2639);
  and g4676 (n3327, n_2628, n_2629);
  not g4677 (n_2640, n3326);
  and g4678 (n3328, n_2640, n3327);
  and g4679 (n3329, n_2636, n_2637);
  not g4680 (n_2641, n3328);
  not g4681 (n_2642, n3329);
  and g4682 (n3330, n_2641, n_2642);
  and g4683 (n3331, n_2638, n3327);
  and g4684 (n3332, n_2639, n3331);
  not g4685 (n_2643, n3327);
  and g4686 (n3333, n_2640, n_2643);
  not g4687 (n_2644, n3332);
  not g4688 (n_2645, n3333);
  and g4689 (n3334, n_2644, n_2645);
  not g4690 (n_2646, n3330);
  not g4691 (n_2647, n3334);
  and g4692 (n3335, n_2646, n_2647);
  not g4693 (n_2648, n3317);
  not g4694 (n_2649, n3335);
  and g4695 (n3336, n_2648, n_2649);
  not g4696 (n_2650, n3300);
  and g4697 (n3337, n_2650, n3336);
  not g4698 (n_2651, n3336);
  and g4699 (n3338, n3300, n_2651);
  not g4700 (n_2652, n3337);
  not g4701 (n_2653, n3338);
  and g4702 (n3339, n_2652, n_2653);
  not g4703 (n_2654, n3264);
  and g4704 (n3340, n_2654, n3339);
  not g4705 (n_2655, n3339);
  and g4706 (n3341, n3264, n_2655);
  not g4707 (n_2656, n3340);
  not g4708 (n_2657, n3341);
  and g4709 (n3342, n_2656, n_2657);
  not g4710 (n_2658, n3189);
  and g4711 (n3343, n_2658, n3342);
  not g4712 (n_2659, n3342);
  and g4713 (n3344, n3189, n_2659);
  not g4714 (n_2660, n3343);
  not g4715 (n_2661, n3344);
  and g4716 (n3345, n_2660, n_2661);
  not g4717 (n_2662, n3036);
  and g4718 (n3346, n_2662, n3345);
  not g4719 (n_2663, n3345);
  and g4720 (n3347, n3036, n_2663);
  not g4721 (n_2664, n3346);
  not g4722 (n_2665, n3347);
  and g4723 (n3348, n_2664, n_2665);
  not g4724 (n_2667, \A[649] );
  and g4725 (n3349, n_2667, \A[650] );
  not g4726 (n_2669, \A[650] );
  and g4727 (n3350, \A[649] , n_2669);
  not g4728 (n_2671, n3350);
  and g4729 (n3351, \A[651] , n_2671);
  not g4730 (n_2672, n3349);
  and g4731 (n3352, n_2672, n3351);
  and g4732 (n3353, n_2672, n_2671);
  not g4733 (n_2673, \A[651] );
  not g4734 (n_2674, n3353);
  and g4735 (n3354, n_2673, n_2674);
  not g4736 (n_2675, n3352);
  not g4737 (n_2676, n3354);
  and g4738 (n3355, n_2675, n_2676);
  not g4739 (n_2678, \A[652] );
  and g4740 (n3356, n_2678, \A[653] );
  not g4741 (n_2680, \A[653] );
  and g4742 (n3357, \A[652] , n_2680);
  not g4743 (n_2682, n3357);
  and g4744 (n3358, \A[654] , n_2682);
  not g4745 (n_2683, n3356);
  and g4746 (n3359, n_2683, n3358);
  and g4747 (n3360, n_2683, n_2682);
  not g4748 (n_2684, \A[654] );
  not g4749 (n_2685, n3360);
  and g4750 (n3361, n_2684, n_2685);
  not g4751 (n_2686, n3359);
  not g4752 (n_2687, n3361);
  and g4753 (n3362, n_2686, n_2687);
  not g4754 (n_2688, n3355);
  and g4755 (n3363, n_2688, n3362);
  not g4756 (n_2689, n3362);
  and g4757 (n3364, n3355, n_2689);
  not g4758 (n_2690, n3363);
  not g4759 (n_2691, n3364);
  and g4760 (n3365, n_2690, n_2691);
  and g4761 (n3366, \A[652] , \A[653] );
  and g4762 (n3367, \A[654] , n_2685);
  not g4763 (n_2692, n3366);
  not g4764 (n_2693, n3367);
  and g4765 (n3368, n_2692, n_2693);
  and g4766 (n3369, \A[649] , \A[650] );
  and g4767 (n3370, \A[651] , n_2674);
  not g4768 (n_2694, n3369);
  not g4769 (n_2695, n3370);
  and g4770 (n3371, n_2694, n_2695);
  not g4771 (n_2696, n3368);
  and g4772 (n3372, n_2696, n3371);
  not g4773 (n_2697, n3371);
  and g4774 (n3373, n3368, n_2697);
  not g4775 (n_2698, n3372);
  not g4776 (n_2699, n3373);
  and g4777 (n3374, n_2698, n_2699);
  and g4778 (n3375, n_2688, n_2689);
  not g4779 (n_2700, n3374);
  and g4780 (n3376, n_2700, n3375);
  and g4781 (n3377, n_2696, n_2697);
  not g4782 (n_2701, n3376);
  not g4783 (n_2702, n3377);
  and g4784 (n3378, n_2701, n_2702);
  and g4785 (n3379, n_2698, n3375);
  and g4786 (n3380, n_2699, n3379);
  not g4787 (n_2703, n3375);
  and g4788 (n3381, n_2700, n_2703);
  not g4789 (n_2704, n3380);
  not g4790 (n_2705, n3381);
  and g4791 (n3382, n_2704, n_2705);
  not g4792 (n_2706, n3378);
  not g4793 (n_2707, n3382);
  and g4794 (n3383, n_2706, n_2707);
  not g4795 (n_2708, n3365);
  not g4796 (n_2709, n3383);
  and g4797 (n3384, n_2708, n_2709);
  not g4798 (n_2711, \A[643] );
  and g4799 (n3385, n_2711, \A[644] );
  not g4800 (n_2713, \A[644] );
  and g4801 (n3386, \A[643] , n_2713);
  not g4802 (n_2715, n3386);
  and g4803 (n3387, \A[645] , n_2715);
  not g4804 (n_2716, n3385);
  and g4805 (n3388, n_2716, n3387);
  and g4806 (n3389, n_2716, n_2715);
  not g4807 (n_2717, \A[645] );
  not g4808 (n_2718, n3389);
  and g4809 (n3390, n_2717, n_2718);
  not g4810 (n_2719, n3388);
  not g4811 (n_2720, n3390);
  and g4812 (n3391, n_2719, n_2720);
  not g4813 (n_2722, \A[646] );
  and g4814 (n3392, n_2722, \A[647] );
  not g4815 (n_2724, \A[647] );
  and g4816 (n3393, \A[646] , n_2724);
  not g4817 (n_2726, n3393);
  and g4818 (n3394, \A[648] , n_2726);
  not g4819 (n_2727, n3392);
  and g4820 (n3395, n_2727, n3394);
  and g4821 (n3396, n_2727, n_2726);
  not g4822 (n_2728, \A[648] );
  not g4823 (n_2729, n3396);
  and g4824 (n3397, n_2728, n_2729);
  not g4825 (n_2730, n3395);
  not g4826 (n_2731, n3397);
  and g4827 (n3398, n_2730, n_2731);
  not g4828 (n_2732, n3391);
  and g4829 (n3399, n_2732, n3398);
  not g4830 (n_2733, n3398);
  and g4831 (n3400, n3391, n_2733);
  not g4832 (n_2734, n3399);
  not g4833 (n_2735, n3400);
  and g4834 (n3401, n_2734, n_2735);
  and g4835 (n3402, \A[646] , \A[647] );
  and g4836 (n3403, \A[648] , n_2729);
  not g4837 (n_2736, n3402);
  not g4838 (n_2737, n3403);
  and g4839 (n3404, n_2736, n_2737);
  and g4840 (n3405, \A[643] , \A[644] );
  and g4841 (n3406, \A[645] , n_2718);
  not g4842 (n_2738, n3405);
  not g4843 (n_2739, n3406);
  and g4844 (n3407, n_2738, n_2739);
  not g4845 (n_2740, n3404);
  and g4846 (n3408, n_2740, n3407);
  not g4847 (n_2741, n3407);
  and g4848 (n3409, n3404, n_2741);
  not g4849 (n_2742, n3408);
  not g4850 (n_2743, n3409);
  and g4851 (n3410, n_2742, n_2743);
  and g4852 (n3411, n_2732, n_2733);
  not g4853 (n_2744, n3410);
  and g4854 (n3412, n_2744, n3411);
  and g4855 (n3413, n_2740, n_2741);
  not g4856 (n_2745, n3412);
  not g4857 (n_2746, n3413);
  and g4858 (n3414, n_2745, n_2746);
  and g4859 (n3415, n_2742, n3411);
  and g4860 (n3416, n_2743, n3415);
  not g4861 (n_2747, n3411);
  and g4862 (n3417, n_2744, n_2747);
  not g4863 (n_2748, n3416);
  not g4864 (n_2749, n3417);
  and g4865 (n3418, n_2748, n_2749);
  not g4866 (n_2750, n3414);
  not g4867 (n_2751, n3418);
  and g4868 (n3419, n_2750, n_2751);
  not g4869 (n_2752, n3401);
  not g4870 (n_2753, n3419);
  and g4871 (n3420, n_2752, n_2753);
  not g4872 (n_2754, n3384);
  and g4873 (n3421, n_2754, n3420);
  not g4874 (n_2755, n3420);
  and g4875 (n3422, n3384, n_2755);
  not g4876 (n_2756, n3421);
  not g4877 (n_2757, n3422);
  and g4878 (n3423, n_2756, n_2757);
  not g4879 (n_2759, \A[637] );
  and g4880 (n3424, n_2759, \A[638] );
  not g4881 (n_2761, \A[638] );
  and g4882 (n3425, \A[637] , n_2761);
  not g4883 (n_2763, n3425);
  and g4884 (n3426, \A[639] , n_2763);
  not g4885 (n_2764, n3424);
  and g4886 (n3427, n_2764, n3426);
  and g4887 (n3428, n_2764, n_2763);
  not g4888 (n_2765, \A[639] );
  not g4889 (n_2766, n3428);
  and g4890 (n3429, n_2765, n_2766);
  not g4891 (n_2767, n3427);
  not g4892 (n_2768, n3429);
  and g4893 (n3430, n_2767, n_2768);
  not g4894 (n_2770, \A[640] );
  and g4895 (n3431, n_2770, \A[641] );
  not g4896 (n_2772, \A[641] );
  and g4897 (n3432, \A[640] , n_2772);
  not g4898 (n_2774, n3432);
  and g4899 (n3433, \A[642] , n_2774);
  not g4900 (n_2775, n3431);
  and g4901 (n3434, n_2775, n3433);
  and g4902 (n3435, n_2775, n_2774);
  not g4903 (n_2776, \A[642] );
  not g4904 (n_2777, n3435);
  and g4905 (n3436, n_2776, n_2777);
  not g4906 (n_2778, n3434);
  not g4907 (n_2779, n3436);
  and g4908 (n3437, n_2778, n_2779);
  not g4909 (n_2780, n3430);
  and g4910 (n3438, n_2780, n3437);
  not g4911 (n_2781, n3437);
  and g4912 (n3439, n3430, n_2781);
  not g4913 (n_2782, n3438);
  not g4914 (n_2783, n3439);
  and g4915 (n3440, n_2782, n_2783);
  and g4916 (n3441, \A[640] , \A[641] );
  and g4917 (n3442, \A[642] , n_2777);
  not g4918 (n_2784, n3441);
  not g4919 (n_2785, n3442);
  and g4920 (n3443, n_2784, n_2785);
  and g4921 (n3444, \A[637] , \A[638] );
  and g4922 (n3445, \A[639] , n_2766);
  not g4923 (n_2786, n3444);
  not g4924 (n_2787, n3445);
  and g4925 (n3446, n_2786, n_2787);
  not g4926 (n_2788, n3443);
  and g4927 (n3447, n_2788, n3446);
  not g4928 (n_2789, n3446);
  and g4929 (n3448, n3443, n_2789);
  not g4930 (n_2790, n3447);
  not g4931 (n_2791, n3448);
  and g4932 (n3449, n_2790, n_2791);
  and g4933 (n3450, n_2780, n_2781);
  not g4934 (n_2792, n3449);
  and g4935 (n3451, n_2792, n3450);
  and g4936 (n3452, n_2788, n_2789);
  not g4937 (n_2793, n3451);
  not g4938 (n_2794, n3452);
  and g4939 (n3453, n_2793, n_2794);
  and g4940 (n3454, n_2790, n3450);
  and g4941 (n3455, n_2791, n3454);
  not g4942 (n_2795, n3450);
  and g4943 (n3456, n_2792, n_2795);
  not g4944 (n_2796, n3455);
  not g4945 (n_2797, n3456);
  and g4946 (n3457, n_2796, n_2797);
  not g4947 (n_2798, n3453);
  not g4948 (n_2799, n3457);
  and g4949 (n3458, n_2798, n_2799);
  not g4950 (n_2800, n3440);
  not g4951 (n_2801, n3458);
  and g4952 (n3459, n_2800, n_2801);
  not g4953 (n_2803, \A[631] );
  and g4954 (n3460, n_2803, \A[632] );
  not g4955 (n_2805, \A[632] );
  and g4956 (n3461, \A[631] , n_2805);
  not g4957 (n_2807, n3461);
  and g4958 (n3462, \A[633] , n_2807);
  not g4959 (n_2808, n3460);
  and g4960 (n3463, n_2808, n3462);
  and g4961 (n3464, n_2808, n_2807);
  not g4962 (n_2809, \A[633] );
  not g4963 (n_2810, n3464);
  and g4964 (n3465, n_2809, n_2810);
  not g4965 (n_2811, n3463);
  not g4966 (n_2812, n3465);
  and g4967 (n3466, n_2811, n_2812);
  not g4968 (n_2814, \A[634] );
  and g4969 (n3467, n_2814, \A[635] );
  not g4970 (n_2816, \A[635] );
  and g4971 (n3468, \A[634] , n_2816);
  not g4972 (n_2818, n3468);
  and g4973 (n3469, \A[636] , n_2818);
  not g4974 (n_2819, n3467);
  and g4975 (n3470, n_2819, n3469);
  and g4976 (n3471, n_2819, n_2818);
  not g4977 (n_2820, \A[636] );
  not g4978 (n_2821, n3471);
  and g4979 (n3472, n_2820, n_2821);
  not g4980 (n_2822, n3470);
  not g4981 (n_2823, n3472);
  and g4982 (n3473, n_2822, n_2823);
  not g4983 (n_2824, n3466);
  and g4984 (n3474, n_2824, n3473);
  not g4985 (n_2825, n3473);
  and g4986 (n3475, n3466, n_2825);
  not g4987 (n_2826, n3474);
  not g4988 (n_2827, n3475);
  and g4989 (n3476, n_2826, n_2827);
  and g4990 (n3477, \A[634] , \A[635] );
  and g4991 (n3478, \A[636] , n_2821);
  not g4992 (n_2828, n3477);
  not g4993 (n_2829, n3478);
  and g4994 (n3479, n_2828, n_2829);
  and g4995 (n3480, \A[631] , \A[632] );
  and g4996 (n3481, \A[633] , n_2810);
  not g4997 (n_2830, n3480);
  not g4998 (n_2831, n3481);
  and g4999 (n3482, n_2830, n_2831);
  not g5000 (n_2832, n3479);
  and g5001 (n3483, n_2832, n3482);
  not g5002 (n_2833, n3482);
  and g5003 (n3484, n3479, n_2833);
  not g5004 (n_2834, n3483);
  not g5005 (n_2835, n3484);
  and g5006 (n3485, n_2834, n_2835);
  and g5007 (n3486, n_2824, n_2825);
  not g5008 (n_2836, n3485);
  and g5009 (n3487, n_2836, n3486);
  and g5010 (n3488, n_2832, n_2833);
  not g5011 (n_2837, n3487);
  not g5012 (n_2838, n3488);
  and g5013 (n3489, n_2837, n_2838);
  and g5014 (n3490, n_2834, n3486);
  and g5015 (n3491, n_2835, n3490);
  not g5016 (n_2839, n3486);
  and g5017 (n3492, n_2836, n_2839);
  not g5018 (n_2840, n3491);
  not g5019 (n_2841, n3492);
  and g5020 (n3493, n_2840, n_2841);
  not g5021 (n_2842, n3489);
  not g5022 (n_2843, n3493);
  and g5023 (n3494, n_2842, n_2843);
  not g5024 (n_2844, n3476);
  not g5025 (n_2845, n3494);
  and g5026 (n3495, n_2844, n_2845);
  not g5027 (n_2846, n3459);
  and g5028 (n3496, n_2846, n3495);
  not g5029 (n_2847, n3495);
  and g5030 (n3497, n3459, n_2847);
  not g5031 (n_2848, n3496);
  not g5032 (n_2849, n3497);
  and g5033 (n3498, n_2848, n_2849);
  not g5034 (n_2850, n3423);
  and g5035 (n3499, n_2850, n3498);
  not g5036 (n_2851, n3498);
  and g5037 (n3500, n3423, n_2851);
  not g5038 (n_2852, n3499);
  not g5039 (n_2853, n3500);
  and g5040 (n3501, n_2852, n_2853);
  not g5041 (n_2855, \A[625] );
  and g5042 (n3502, n_2855, \A[626] );
  not g5043 (n_2857, \A[626] );
  and g5044 (n3503, \A[625] , n_2857);
  not g5045 (n_2859, n3503);
  and g5046 (n3504, \A[627] , n_2859);
  not g5047 (n_2860, n3502);
  and g5048 (n3505, n_2860, n3504);
  and g5049 (n3506, n_2860, n_2859);
  not g5050 (n_2861, \A[627] );
  not g5051 (n_2862, n3506);
  and g5052 (n3507, n_2861, n_2862);
  not g5053 (n_2863, n3505);
  not g5054 (n_2864, n3507);
  and g5055 (n3508, n_2863, n_2864);
  not g5056 (n_2866, \A[628] );
  and g5057 (n3509, n_2866, \A[629] );
  not g5058 (n_2868, \A[629] );
  and g5059 (n3510, \A[628] , n_2868);
  not g5060 (n_2870, n3510);
  and g5061 (n3511, \A[630] , n_2870);
  not g5062 (n_2871, n3509);
  and g5063 (n3512, n_2871, n3511);
  and g5064 (n3513, n_2871, n_2870);
  not g5065 (n_2872, \A[630] );
  not g5066 (n_2873, n3513);
  and g5067 (n3514, n_2872, n_2873);
  not g5068 (n_2874, n3512);
  not g5069 (n_2875, n3514);
  and g5070 (n3515, n_2874, n_2875);
  not g5071 (n_2876, n3508);
  and g5072 (n3516, n_2876, n3515);
  not g5073 (n_2877, n3515);
  and g5074 (n3517, n3508, n_2877);
  not g5075 (n_2878, n3516);
  not g5076 (n_2879, n3517);
  and g5077 (n3518, n_2878, n_2879);
  and g5078 (n3519, \A[628] , \A[629] );
  and g5079 (n3520, \A[630] , n_2873);
  not g5080 (n_2880, n3519);
  not g5081 (n_2881, n3520);
  and g5082 (n3521, n_2880, n_2881);
  and g5083 (n3522, \A[625] , \A[626] );
  and g5084 (n3523, \A[627] , n_2862);
  not g5085 (n_2882, n3522);
  not g5086 (n_2883, n3523);
  and g5087 (n3524, n_2882, n_2883);
  not g5088 (n_2884, n3521);
  and g5089 (n3525, n_2884, n3524);
  not g5090 (n_2885, n3524);
  and g5091 (n3526, n3521, n_2885);
  not g5092 (n_2886, n3525);
  not g5093 (n_2887, n3526);
  and g5094 (n3527, n_2886, n_2887);
  and g5095 (n3528, n_2876, n_2877);
  not g5096 (n_2888, n3527);
  and g5097 (n3529, n_2888, n3528);
  and g5098 (n3530, n_2884, n_2885);
  not g5099 (n_2889, n3529);
  not g5100 (n_2890, n3530);
  and g5101 (n3531, n_2889, n_2890);
  and g5102 (n3532, n_2886, n3528);
  and g5103 (n3533, n_2887, n3532);
  not g5104 (n_2891, n3528);
  and g5105 (n3534, n_2888, n_2891);
  not g5106 (n_2892, n3533);
  not g5107 (n_2893, n3534);
  and g5108 (n3535, n_2892, n_2893);
  not g5109 (n_2894, n3531);
  not g5110 (n_2895, n3535);
  and g5111 (n3536, n_2894, n_2895);
  not g5112 (n_2896, n3518);
  not g5113 (n_2897, n3536);
  and g5114 (n3537, n_2896, n_2897);
  not g5115 (n_2899, \A[619] );
  and g5116 (n3538, n_2899, \A[620] );
  not g5117 (n_2901, \A[620] );
  and g5118 (n3539, \A[619] , n_2901);
  not g5119 (n_2903, n3539);
  and g5120 (n3540, \A[621] , n_2903);
  not g5121 (n_2904, n3538);
  and g5122 (n3541, n_2904, n3540);
  and g5123 (n3542, n_2904, n_2903);
  not g5124 (n_2905, \A[621] );
  not g5125 (n_2906, n3542);
  and g5126 (n3543, n_2905, n_2906);
  not g5127 (n_2907, n3541);
  not g5128 (n_2908, n3543);
  and g5129 (n3544, n_2907, n_2908);
  not g5130 (n_2910, \A[622] );
  and g5131 (n3545, n_2910, \A[623] );
  not g5132 (n_2912, \A[623] );
  and g5133 (n3546, \A[622] , n_2912);
  not g5134 (n_2914, n3546);
  and g5135 (n3547, \A[624] , n_2914);
  not g5136 (n_2915, n3545);
  and g5137 (n3548, n_2915, n3547);
  and g5138 (n3549, n_2915, n_2914);
  not g5139 (n_2916, \A[624] );
  not g5140 (n_2917, n3549);
  and g5141 (n3550, n_2916, n_2917);
  not g5142 (n_2918, n3548);
  not g5143 (n_2919, n3550);
  and g5144 (n3551, n_2918, n_2919);
  not g5145 (n_2920, n3544);
  and g5146 (n3552, n_2920, n3551);
  not g5147 (n_2921, n3551);
  and g5148 (n3553, n3544, n_2921);
  not g5149 (n_2922, n3552);
  not g5150 (n_2923, n3553);
  and g5151 (n3554, n_2922, n_2923);
  and g5152 (n3555, \A[622] , \A[623] );
  and g5153 (n3556, \A[624] , n_2917);
  not g5154 (n_2924, n3555);
  not g5155 (n_2925, n3556);
  and g5156 (n3557, n_2924, n_2925);
  and g5157 (n3558, \A[619] , \A[620] );
  and g5158 (n3559, \A[621] , n_2906);
  not g5159 (n_2926, n3558);
  not g5160 (n_2927, n3559);
  and g5161 (n3560, n_2926, n_2927);
  not g5162 (n_2928, n3557);
  and g5163 (n3561, n_2928, n3560);
  not g5164 (n_2929, n3560);
  and g5165 (n3562, n3557, n_2929);
  not g5166 (n_2930, n3561);
  not g5167 (n_2931, n3562);
  and g5168 (n3563, n_2930, n_2931);
  and g5169 (n3564, n_2920, n_2921);
  not g5170 (n_2932, n3563);
  and g5171 (n3565, n_2932, n3564);
  and g5172 (n3566, n_2928, n_2929);
  not g5173 (n_2933, n3565);
  not g5174 (n_2934, n3566);
  and g5175 (n3567, n_2933, n_2934);
  and g5176 (n3568, n_2930, n3564);
  and g5177 (n3569, n_2931, n3568);
  not g5178 (n_2935, n3564);
  and g5179 (n3570, n_2932, n_2935);
  not g5180 (n_2936, n3569);
  not g5181 (n_2937, n3570);
  and g5182 (n3571, n_2936, n_2937);
  not g5183 (n_2938, n3567);
  not g5184 (n_2939, n3571);
  and g5185 (n3572, n_2938, n_2939);
  not g5186 (n_2940, n3554);
  not g5187 (n_2941, n3572);
  and g5188 (n3573, n_2940, n_2941);
  not g5189 (n_2942, n3537);
  and g5190 (n3574, n_2942, n3573);
  not g5191 (n_2943, n3573);
  and g5192 (n3575, n3537, n_2943);
  not g5193 (n_2944, n3574);
  not g5194 (n_2945, n3575);
  and g5195 (n3576, n_2944, n_2945);
  not g5196 (n_2947, \A[613] );
  and g5197 (n3577, n_2947, \A[614] );
  not g5198 (n_2949, \A[614] );
  and g5199 (n3578, \A[613] , n_2949);
  not g5200 (n_2951, n3578);
  and g5201 (n3579, \A[615] , n_2951);
  not g5202 (n_2952, n3577);
  and g5203 (n3580, n_2952, n3579);
  and g5204 (n3581, n_2952, n_2951);
  not g5205 (n_2953, \A[615] );
  not g5206 (n_2954, n3581);
  and g5207 (n3582, n_2953, n_2954);
  not g5208 (n_2955, n3580);
  not g5209 (n_2956, n3582);
  and g5210 (n3583, n_2955, n_2956);
  not g5211 (n_2958, \A[616] );
  and g5212 (n3584, n_2958, \A[617] );
  not g5213 (n_2960, \A[617] );
  and g5214 (n3585, \A[616] , n_2960);
  not g5215 (n_2962, n3585);
  and g5216 (n3586, \A[618] , n_2962);
  not g5217 (n_2963, n3584);
  and g5218 (n3587, n_2963, n3586);
  and g5219 (n3588, n_2963, n_2962);
  not g5220 (n_2964, \A[618] );
  not g5221 (n_2965, n3588);
  and g5222 (n3589, n_2964, n_2965);
  not g5223 (n_2966, n3587);
  not g5224 (n_2967, n3589);
  and g5225 (n3590, n_2966, n_2967);
  not g5226 (n_2968, n3583);
  and g5227 (n3591, n_2968, n3590);
  not g5228 (n_2969, n3590);
  and g5229 (n3592, n3583, n_2969);
  not g5230 (n_2970, n3591);
  not g5231 (n_2971, n3592);
  and g5232 (n3593, n_2970, n_2971);
  and g5233 (n3594, \A[616] , \A[617] );
  and g5234 (n3595, \A[618] , n_2965);
  not g5235 (n_2972, n3594);
  not g5236 (n_2973, n3595);
  and g5237 (n3596, n_2972, n_2973);
  and g5238 (n3597, \A[613] , \A[614] );
  and g5239 (n3598, \A[615] , n_2954);
  not g5240 (n_2974, n3597);
  not g5241 (n_2975, n3598);
  and g5242 (n3599, n_2974, n_2975);
  not g5243 (n_2976, n3596);
  and g5244 (n3600, n_2976, n3599);
  not g5245 (n_2977, n3599);
  and g5246 (n3601, n3596, n_2977);
  not g5247 (n_2978, n3600);
  not g5248 (n_2979, n3601);
  and g5249 (n3602, n_2978, n_2979);
  and g5250 (n3603, n_2968, n_2969);
  not g5251 (n_2980, n3602);
  and g5252 (n3604, n_2980, n3603);
  and g5253 (n3605, n_2976, n_2977);
  not g5254 (n_2981, n3604);
  not g5255 (n_2982, n3605);
  and g5256 (n3606, n_2981, n_2982);
  and g5257 (n3607, n_2978, n3603);
  and g5258 (n3608, n_2979, n3607);
  not g5259 (n_2983, n3603);
  and g5260 (n3609, n_2980, n_2983);
  not g5261 (n_2984, n3608);
  not g5262 (n_2985, n3609);
  and g5263 (n3610, n_2984, n_2985);
  not g5264 (n_2986, n3606);
  not g5265 (n_2987, n3610);
  and g5266 (n3611, n_2986, n_2987);
  not g5267 (n_2988, n3593);
  not g5268 (n_2989, n3611);
  and g5269 (n3612, n_2988, n_2989);
  not g5270 (n_2991, \A[607] );
  and g5271 (n3613, n_2991, \A[608] );
  not g5272 (n_2993, \A[608] );
  and g5273 (n3614, \A[607] , n_2993);
  not g5274 (n_2995, n3614);
  and g5275 (n3615, \A[609] , n_2995);
  not g5276 (n_2996, n3613);
  and g5277 (n3616, n_2996, n3615);
  and g5278 (n3617, n_2996, n_2995);
  not g5279 (n_2997, \A[609] );
  not g5280 (n_2998, n3617);
  and g5281 (n3618, n_2997, n_2998);
  not g5282 (n_2999, n3616);
  not g5283 (n_3000, n3618);
  and g5284 (n3619, n_2999, n_3000);
  not g5285 (n_3002, \A[610] );
  and g5286 (n3620, n_3002, \A[611] );
  not g5287 (n_3004, \A[611] );
  and g5288 (n3621, \A[610] , n_3004);
  not g5289 (n_3006, n3621);
  and g5290 (n3622, \A[612] , n_3006);
  not g5291 (n_3007, n3620);
  and g5292 (n3623, n_3007, n3622);
  and g5293 (n3624, n_3007, n_3006);
  not g5294 (n_3008, \A[612] );
  not g5295 (n_3009, n3624);
  and g5296 (n3625, n_3008, n_3009);
  not g5297 (n_3010, n3623);
  not g5298 (n_3011, n3625);
  and g5299 (n3626, n_3010, n_3011);
  not g5300 (n_3012, n3619);
  and g5301 (n3627, n_3012, n3626);
  not g5302 (n_3013, n3626);
  and g5303 (n3628, n3619, n_3013);
  not g5304 (n_3014, n3627);
  not g5305 (n_3015, n3628);
  and g5306 (n3629, n_3014, n_3015);
  and g5307 (n3630, \A[610] , \A[611] );
  and g5308 (n3631, \A[612] , n_3009);
  not g5309 (n_3016, n3630);
  not g5310 (n_3017, n3631);
  and g5311 (n3632, n_3016, n_3017);
  and g5312 (n3633, \A[607] , \A[608] );
  and g5313 (n3634, \A[609] , n_2998);
  not g5314 (n_3018, n3633);
  not g5315 (n_3019, n3634);
  and g5316 (n3635, n_3018, n_3019);
  not g5317 (n_3020, n3632);
  and g5318 (n3636, n_3020, n3635);
  not g5319 (n_3021, n3635);
  and g5320 (n3637, n3632, n_3021);
  not g5321 (n_3022, n3636);
  not g5322 (n_3023, n3637);
  and g5323 (n3638, n_3022, n_3023);
  and g5324 (n3639, n_3012, n_3013);
  not g5325 (n_3024, n3638);
  and g5326 (n3640, n_3024, n3639);
  and g5327 (n3641, n_3020, n_3021);
  not g5328 (n_3025, n3640);
  not g5329 (n_3026, n3641);
  and g5330 (n3642, n_3025, n_3026);
  and g5331 (n3643, n_3022, n3639);
  and g5332 (n3644, n_3023, n3643);
  not g5333 (n_3027, n3639);
  and g5334 (n3645, n_3024, n_3027);
  not g5335 (n_3028, n3644);
  not g5336 (n_3029, n3645);
  and g5337 (n3646, n_3028, n_3029);
  not g5338 (n_3030, n3642);
  not g5339 (n_3031, n3646);
  and g5340 (n3647, n_3030, n_3031);
  not g5341 (n_3032, n3629);
  not g5342 (n_3033, n3647);
  and g5343 (n3648, n_3032, n_3033);
  not g5344 (n_3034, n3612);
  and g5345 (n3649, n_3034, n3648);
  not g5346 (n_3035, n3648);
  and g5347 (n3650, n3612, n_3035);
  not g5348 (n_3036, n3649);
  not g5349 (n_3037, n3650);
  and g5350 (n3651, n_3036, n_3037);
  not g5351 (n_3038, n3576);
  and g5352 (n3652, n_3038, n3651);
  not g5353 (n_3039, n3651);
  and g5354 (n3653, n3576, n_3039);
  not g5355 (n_3040, n3652);
  not g5356 (n_3041, n3653);
  and g5357 (n3654, n_3040, n_3041);
  not g5358 (n_3042, n3501);
  and g5359 (n3655, n_3042, n3654);
  not g5360 (n_3043, n3654);
  and g5361 (n3656, n3501, n_3043);
  not g5362 (n_3044, n3655);
  not g5363 (n_3045, n3656);
  and g5364 (n3657, n_3044, n_3045);
  not g5365 (n_3047, \A[601] );
  and g5366 (n3658, n_3047, \A[602] );
  not g5367 (n_3049, \A[602] );
  and g5368 (n3659, \A[601] , n_3049);
  not g5369 (n_3051, n3659);
  and g5370 (n3660, \A[603] , n_3051);
  not g5371 (n_3052, n3658);
  and g5372 (n3661, n_3052, n3660);
  and g5373 (n3662, n_3052, n_3051);
  not g5374 (n_3053, \A[603] );
  not g5375 (n_3054, n3662);
  and g5376 (n3663, n_3053, n_3054);
  not g5377 (n_3055, n3661);
  not g5378 (n_3056, n3663);
  and g5379 (n3664, n_3055, n_3056);
  not g5380 (n_3058, \A[604] );
  and g5381 (n3665, n_3058, \A[605] );
  not g5382 (n_3060, \A[605] );
  and g5383 (n3666, \A[604] , n_3060);
  not g5384 (n_3062, n3666);
  and g5385 (n3667, \A[606] , n_3062);
  not g5386 (n_3063, n3665);
  and g5387 (n3668, n_3063, n3667);
  and g5388 (n3669, n_3063, n_3062);
  not g5389 (n_3064, \A[606] );
  not g5390 (n_3065, n3669);
  and g5391 (n3670, n_3064, n_3065);
  not g5392 (n_3066, n3668);
  not g5393 (n_3067, n3670);
  and g5394 (n3671, n_3066, n_3067);
  not g5395 (n_3068, n3664);
  and g5396 (n3672, n_3068, n3671);
  not g5397 (n_3069, n3671);
  and g5398 (n3673, n3664, n_3069);
  not g5399 (n_3070, n3672);
  not g5400 (n_3071, n3673);
  and g5401 (n3674, n_3070, n_3071);
  and g5402 (n3675, \A[604] , \A[605] );
  and g5403 (n3676, \A[606] , n_3065);
  not g5404 (n_3072, n3675);
  not g5405 (n_3073, n3676);
  and g5406 (n3677, n_3072, n_3073);
  and g5407 (n3678, \A[601] , \A[602] );
  and g5408 (n3679, \A[603] , n_3054);
  not g5409 (n_3074, n3678);
  not g5410 (n_3075, n3679);
  and g5411 (n3680, n_3074, n_3075);
  not g5412 (n_3076, n3677);
  and g5413 (n3681, n_3076, n3680);
  not g5414 (n_3077, n3680);
  and g5415 (n3682, n3677, n_3077);
  not g5416 (n_3078, n3681);
  not g5417 (n_3079, n3682);
  and g5418 (n3683, n_3078, n_3079);
  and g5419 (n3684, n_3068, n_3069);
  not g5420 (n_3080, n3683);
  and g5421 (n3685, n_3080, n3684);
  and g5422 (n3686, n_3076, n_3077);
  not g5423 (n_3081, n3685);
  not g5424 (n_3082, n3686);
  and g5425 (n3687, n_3081, n_3082);
  and g5426 (n3688, n_3078, n3684);
  and g5427 (n3689, n_3079, n3688);
  not g5428 (n_3083, n3684);
  and g5429 (n3690, n_3080, n_3083);
  not g5430 (n_3084, n3689);
  not g5431 (n_3085, n3690);
  and g5432 (n3691, n_3084, n_3085);
  not g5433 (n_3086, n3687);
  not g5434 (n_3087, n3691);
  and g5435 (n3692, n_3086, n_3087);
  not g5436 (n_3088, n3674);
  not g5437 (n_3089, n3692);
  and g5438 (n3693, n_3088, n_3089);
  not g5439 (n_3091, \A[595] );
  and g5440 (n3694, n_3091, \A[596] );
  not g5441 (n_3093, \A[596] );
  and g5442 (n3695, \A[595] , n_3093);
  not g5443 (n_3095, n3695);
  and g5444 (n3696, \A[597] , n_3095);
  not g5445 (n_3096, n3694);
  and g5446 (n3697, n_3096, n3696);
  and g5447 (n3698, n_3096, n_3095);
  not g5448 (n_3097, \A[597] );
  not g5449 (n_3098, n3698);
  and g5450 (n3699, n_3097, n_3098);
  not g5451 (n_3099, n3697);
  not g5452 (n_3100, n3699);
  and g5453 (n3700, n_3099, n_3100);
  not g5454 (n_3102, \A[598] );
  and g5455 (n3701, n_3102, \A[599] );
  not g5456 (n_3104, \A[599] );
  and g5457 (n3702, \A[598] , n_3104);
  not g5458 (n_3106, n3702);
  and g5459 (n3703, \A[600] , n_3106);
  not g5460 (n_3107, n3701);
  and g5461 (n3704, n_3107, n3703);
  and g5462 (n3705, n_3107, n_3106);
  not g5463 (n_3108, \A[600] );
  not g5464 (n_3109, n3705);
  and g5465 (n3706, n_3108, n_3109);
  not g5466 (n_3110, n3704);
  not g5467 (n_3111, n3706);
  and g5468 (n3707, n_3110, n_3111);
  not g5469 (n_3112, n3700);
  and g5470 (n3708, n_3112, n3707);
  not g5471 (n_3113, n3707);
  and g5472 (n3709, n3700, n_3113);
  not g5473 (n_3114, n3708);
  not g5474 (n_3115, n3709);
  and g5475 (n3710, n_3114, n_3115);
  and g5476 (n3711, \A[598] , \A[599] );
  and g5477 (n3712, \A[600] , n_3109);
  not g5478 (n_3116, n3711);
  not g5479 (n_3117, n3712);
  and g5480 (n3713, n_3116, n_3117);
  and g5481 (n3714, \A[595] , \A[596] );
  and g5482 (n3715, \A[597] , n_3098);
  not g5483 (n_3118, n3714);
  not g5484 (n_3119, n3715);
  and g5485 (n3716, n_3118, n_3119);
  not g5486 (n_3120, n3713);
  and g5487 (n3717, n_3120, n3716);
  not g5488 (n_3121, n3716);
  and g5489 (n3718, n3713, n_3121);
  not g5490 (n_3122, n3717);
  not g5491 (n_3123, n3718);
  and g5492 (n3719, n_3122, n_3123);
  and g5493 (n3720, n_3112, n_3113);
  not g5494 (n_3124, n3719);
  and g5495 (n3721, n_3124, n3720);
  and g5496 (n3722, n_3120, n_3121);
  not g5497 (n_3125, n3721);
  not g5498 (n_3126, n3722);
  and g5499 (n3723, n_3125, n_3126);
  and g5500 (n3724, n_3122, n3720);
  and g5501 (n3725, n_3123, n3724);
  not g5502 (n_3127, n3720);
  and g5503 (n3726, n_3124, n_3127);
  not g5504 (n_3128, n3725);
  not g5505 (n_3129, n3726);
  and g5506 (n3727, n_3128, n_3129);
  not g5507 (n_3130, n3723);
  not g5508 (n_3131, n3727);
  and g5509 (n3728, n_3130, n_3131);
  not g5510 (n_3132, n3710);
  not g5511 (n_3133, n3728);
  and g5512 (n3729, n_3132, n_3133);
  not g5513 (n_3134, n3693);
  and g5514 (n3730, n_3134, n3729);
  not g5515 (n_3135, n3729);
  and g5516 (n3731, n3693, n_3135);
  not g5517 (n_3136, n3730);
  not g5518 (n_3137, n3731);
  and g5519 (n3732, n_3136, n_3137);
  not g5520 (n_3139, \A[589] );
  and g5521 (n3733, n_3139, \A[590] );
  not g5522 (n_3141, \A[590] );
  and g5523 (n3734, \A[589] , n_3141);
  not g5524 (n_3143, n3734);
  and g5525 (n3735, \A[591] , n_3143);
  not g5526 (n_3144, n3733);
  and g5527 (n3736, n_3144, n3735);
  and g5528 (n3737, n_3144, n_3143);
  not g5529 (n_3145, \A[591] );
  not g5530 (n_3146, n3737);
  and g5531 (n3738, n_3145, n_3146);
  not g5532 (n_3147, n3736);
  not g5533 (n_3148, n3738);
  and g5534 (n3739, n_3147, n_3148);
  not g5535 (n_3150, \A[592] );
  and g5536 (n3740, n_3150, \A[593] );
  not g5537 (n_3152, \A[593] );
  and g5538 (n3741, \A[592] , n_3152);
  not g5539 (n_3154, n3741);
  and g5540 (n3742, \A[594] , n_3154);
  not g5541 (n_3155, n3740);
  and g5542 (n3743, n_3155, n3742);
  and g5543 (n3744, n_3155, n_3154);
  not g5544 (n_3156, \A[594] );
  not g5545 (n_3157, n3744);
  and g5546 (n3745, n_3156, n_3157);
  not g5547 (n_3158, n3743);
  not g5548 (n_3159, n3745);
  and g5549 (n3746, n_3158, n_3159);
  not g5550 (n_3160, n3739);
  and g5551 (n3747, n_3160, n3746);
  not g5552 (n_3161, n3746);
  and g5553 (n3748, n3739, n_3161);
  not g5554 (n_3162, n3747);
  not g5555 (n_3163, n3748);
  and g5556 (n3749, n_3162, n_3163);
  and g5557 (n3750, \A[592] , \A[593] );
  and g5558 (n3751, \A[594] , n_3157);
  not g5559 (n_3164, n3750);
  not g5560 (n_3165, n3751);
  and g5561 (n3752, n_3164, n_3165);
  and g5562 (n3753, \A[589] , \A[590] );
  and g5563 (n3754, \A[591] , n_3146);
  not g5564 (n_3166, n3753);
  not g5565 (n_3167, n3754);
  and g5566 (n3755, n_3166, n_3167);
  not g5567 (n_3168, n3752);
  and g5568 (n3756, n_3168, n3755);
  not g5569 (n_3169, n3755);
  and g5570 (n3757, n3752, n_3169);
  not g5571 (n_3170, n3756);
  not g5572 (n_3171, n3757);
  and g5573 (n3758, n_3170, n_3171);
  and g5574 (n3759, n_3160, n_3161);
  not g5575 (n_3172, n3758);
  and g5576 (n3760, n_3172, n3759);
  and g5577 (n3761, n_3168, n_3169);
  not g5578 (n_3173, n3760);
  not g5579 (n_3174, n3761);
  and g5580 (n3762, n_3173, n_3174);
  and g5581 (n3763, n_3170, n3759);
  and g5582 (n3764, n_3171, n3763);
  not g5583 (n_3175, n3759);
  and g5584 (n3765, n_3172, n_3175);
  not g5585 (n_3176, n3764);
  not g5586 (n_3177, n3765);
  and g5587 (n3766, n_3176, n_3177);
  not g5588 (n_3178, n3762);
  not g5589 (n_3179, n3766);
  and g5590 (n3767, n_3178, n_3179);
  not g5591 (n_3180, n3749);
  not g5592 (n_3181, n3767);
  and g5593 (n3768, n_3180, n_3181);
  not g5594 (n_3183, \A[583] );
  and g5595 (n3769, n_3183, \A[584] );
  not g5596 (n_3185, \A[584] );
  and g5597 (n3770, \A[583] , n_3185);
  not g5598 (n_3187, n3770);
  and g5599 (n3771, \A[585] , n_3187);
  not g5600 (n_3188, n3769);
  and g5601 (n3772, n_3188, n3771);
  and g5602 (n3773, n_3188, n_3187);
  not g5603 (n_3189, \A[585] );
  not g5604 (n_3190, n3773);
  and g5605 (n3774, n_3189, n_3190);
  not g5606 (n_3191, n3772);
  not g5607 (n_3192, n3774);
  and g5608 (n3775, n_3191, n_3192);
  not g5609 (n_3194, \A[586] );
  and g5610 (n3776, n_3194, \A[587] );
  not g5611 (n_3196, \A[587] );
  and g5612 (n3777, \A[586] , n_3196);
  not g5613 (n_3198, n3777);
  and g5614 (n3778, \A[588] , n_3198);
  not g5615 (n_3199, n3776);
  and g5616 (n3779, n_3199, n3778);
  and g5617 (n3780, n_3199, n_3198);
  not g5618 (n_3200, \A[588] );
  not g5619 (n_3201, n3780);
  and g5620 (n3781, n_3200, n_3201);
  not g5621 (n_3202, n3779);
  not g5622 (n_3203, n3781);
  and g5623 (n3782, n_3202, n_3203);
  not g5624 (n_3204, n3775);
  and g5625 (n3783, n_3204, n3782);
  not g5626 (n_3205, n3782);
  and g5627 (n3784, n3775, n_3205);
  not g5628 (n_3206, n3783);
  not g5629 (n_3207, n3784);
  and g5630 (n3785, n_3206, n_3207);
  and g5631 (n3786, \A[586] , \A[587] );
  and g5632 (n3787, \A[588] , n_3201);
  not g5633 (n_3208, n3786);
  not g5634 (n_3209, n3787);
  and g5635 (n3788, n_3208, n_3209);
  and g5636 (n3789, \A[583] , \A[584] );
  and g5637 (n3790, \A[585] , n_3190);
  not g5638 (n_3210, n3789);
  not g5639 (n_3211, n3790);
  and g5640 (n3791, n_3210, n_3211);
  not g5641 (n_3212, n3788);
  and g5642 (n3792, n_3212, n3791);
  not g5643 (n_3213, n3791);
  and g5644 (n3793, n3788, n_3213);
  not g5645 (n_3214, n3792);
  not g5646 (n_3215, n3793);
  and g5647 (n3794, n_3214, n_3215);
  and g5648 (n3795, n_3204, n_3205);
  not g5649 (n_3216, n3794);
  and g5650 (n3796, n_3216, n3795);
  and g5651 (n3797, n_3212, n_3213);
  not g5652 (n_3217, n3796);
  not g5653 (n_3218, n3797);
  and g5654 (n3798, n_3217, n_3218);
  and g5655 (n3799, n_3214, n3795);
  and g5656 (n3800, n_3215, n3799);
  not g5657 (n_3219, n3795);
  and g5658 (n3801, n_3216, n_3219);
  not g5659 (n_3220, n3800);
  not g5660 (n_3221, n3801);
  and g5661 (n3802, n_3220, n_3221);
  not g5662 (n_3222, n3798);
  not g5663 (n_3223, n3802);
  and g5664 (n3803, n_3222, n_3223);
  not g5665 (n_3224, n3785);
  not g5666 (n_3225, n3803);
  and g5667 (n3804, n_3224, n_3225);
  not g5668 (n_3226, n3768);
  and g5669 (n3805, n_3226, n3804);
  not g5670 (n_3227, n3804);
  and g5671 (n3806, n3768, n_3227);
  not g5672 (n_3228, n3805);
  not g5673 (n_3229, n3806);
  and g5674 (n3807, n_3228, n_3229);
  not g5675 (n_3230, n3732);
  and g5676 (n3808, n_3230, n3807);
  not g5677 (n_3231, n3807);
  and g5678 (n3809, n3732, n_3231);
  not g5679 (n_3232, n3808);
  not g5680 (n_3233, n3809);
  and g5681 (n3810, n_3232, n_3233);
  not g5682 (n_3235, \A[577] );
  and g5683 (n3811, n_3235, \A[578] );
  not g5684 (n_3237, \A[578] );
  and g5685 (n3812, \A[577] , n_3237);
  not g5686 (n_3239, n3812);
  and g5687 (n3813, \A[579] , n_3239);
  not g5688 (n_3240, n3811);
  and g5689 (n3814, n_3240, n3813);
  and g5690 (n3815, n_3240, n_3239);
  not g5691 (n_3241, \A[579] );
  not g5692 (n_3242, n3815);
  and g5693 (n3816, n_3241, n_3242);
  not g5694 (n_3243, n3814);
  not g5695 (n_3244, n3816);
  and g5696 (n3817, n_3243, n_3244);
  not g5697 (n_3246, \A[580] );
  and g5698 (n3818, n_3246, \A[581] );
  not g5699 (n_3248, \A[581] );
  and g5700 (n3819, \A[580] , n_3248);
  not g5701 (n_3250, n3819);
  and g5702 (n3820, \A[582] , n_3250);
  not g5703 (n_3251, n3818);
  and g5704 (n3821, n_3251, n3820);
  and g5705 (n3822, n_3251, n_3250);
  not g5706 (n_3252, \A[582] );
  not g5707 (n_3253, n3822);
  and g5708 (n3823, n_3252, n_3253);
  not g5709 (n_3254, n3821);
  not g5710 (n_3255, n3823);
  and g5711 (n3824, n_3254, n_3255);
  not g5712 (n_3256, n3817);
  and g5713 (n3825, n_3256, n3824);
  not g5714 (n_3257, n3824);
  and g5715 (n3826, n3817, n_3257);
  not g5716 (n_3258, n3825);
  not g5717 (n_3259, n3826);
  and g5718 (n3827, n_3258, n_3259);
  and g5719 (n3828, \A[580] , \A[581] );
  and g5720 (n3829, \A[582] , n_3253);
  not g5721 (n_3260, n3828);
  not g5722 (n_3261, n3829);
  and g5723 (n3830, n_3260, n_3261);
  and g5724 (n3831, \A[577] , \A[578] );
  and g5725 (n3832, \A[579] , n_3242);
  not g5726 (n_3262, n3831);
  not g5727 (n_3263, n3832);
  and g5728 (n3833, n_3262, n_3263);
  not g5729 (n_3264, n3830);
  and g5730 (n3834, n_3264, n3833);
  not g5731 (n_3265, n3833);
  and g5732 (n3835, n3830, n_3265);
  not g5733 (n_3266, n3834);
  not g5734 (n_3267, n3835);
  and g5735 (n3836, n_3266, n_3267);
  and g5736 (n3837, n_3256, n_3257);
  not g5737 (n_3268, n3836);
  and g5738 (n3838, n_3268, n3837);
  and g5739 (n3839, n_3264, n_3265);
  not g5740 (n_3269, n3838);
  not g5741 (n_3270, n3839);
  and g5742 (n3840, n_3269, n_3270);
  and g5743 (n3841, n_3266, n3837);
  and g5744 (n3842, n_3267, n3841);
  not g5745 (n_3271, n3837);
  and g5746 (n3843, n_3268, n_3271);
  not g5747 (n_3272, n3842);
  not g5748 (n_3273, n3843);
  and g5749 (n3844, n_3272, n_3273);
  not g5750 (n_3274, n3840);
  not g5751 (n_3275, n3844);
  and g5752 (n3845, n_3274, n_3275);
  not g5753 (n_3276, n3827);
  not g5754 (n_3277, n3845);
  and g5755 (n3846, n_3276, n_3277);
  not g5756 (n_3279, \A[571] );
  and g5757 (n3847, n_3279, \A[572] );
  not g5758 (n_3281, \A[572] );
  and g5759 (n3848, \A[571] , n_3281);
  not g5760 (n_3283, n3848);
  and g5761 (n3849, \A[573] , n_3283);
  not g5762 (n_3284, n3847);
  and g5763 (n3850, n_3284, n3849);
  and g5764 (n3851, n_3284, n_3283);
  not g5765 (n_3285, \A[573] );
  not g5766 (n_3286, n3851);
  and g5767 (n3852, n_3285, n_3286);
  not g5768 (n_3287, n3850);
  not g5769 (n_3288, n3852);
  and g5770 (n3853, n_3287, n_3288);
  not g5771 (n_3290, \A[574] );
  and g5772 (n3854, n_3290, \A[575] );
  not g5773 (n_3292, \A[575] );
  and g5774 (n3855, \A[574] , n_3292);
  not g5775 (n_3294, n3855);
  and g5776 (n3856, \A[576] , n_3294);
  not g5777 (n_3295, n3854);
  and g5778 (n3857, n_3295, n3856);
  and g5779 (n3858, n_3295, n_3294);
  not g5780 (n_3296, \A[576] );
  not g5781 (n_3297, n3858);
  and g5782 (n3859, n_3296, n_3297);
  not g5783 (n_3298, n3857);
  not g5784 (n_3299, n3859);
  and g5785 (n3860, n_3298, n_3299);
  not g5786 (n_3300, n3853);
  and g5787 (n3861, n_3300, n3860);
  not g5788 (n_3301, n3860);
  and g5789 (n3862, n3853, n_3301);
  not g5790 (n_3302, n3861);
  not g5791 (n_3303, n3862);
  and g5792 (n3863, n_3302, n_3303);
  and g5793 (n3864, \A[574] , \A[575] );
  and g5794 (n3865, \A[576] , n_3297);
  not g5795 (n_3304, n3864);
  not g5796 (n_3305, n3865);
  and g5797 (n3866, n_3304, n_3305);
  and g5798 (n3867, \A[571] , \A[572] );
  and g5799 (n3868, \A[573] , n_3286);
  not g5800 (n_3306, n3867);
  not g5801 (n_3307, n3868);
  and g5802 (n3869, n_3306, n_3307);
  not g5803 (n_3308, n3866);
  and g5804 (n3870, n_3308, n3869);
  not g5805 (n_3309, n3869);
  and g5806 (n3871, n3866, n_3309);
  not g5807 (n_3310, n3870);
  not g5808 (n_3311, n3871);
  and g5809 (n3872, n_3310, n_3311);
  and g5810 (n3873, n_3300, n_3301);
  not g5811 (n_3312, n3872);
  and g5812 (n3874, n_3312, n3873);
  and g5813 (n3875, n_3308, n_3309);
  not g5814 (n_3313, n3874);
  not g5815 (n_3314, n3875);
  and g5816 (n3876, n_3313, n_3314);
  and g5817 (n3877, n_3310, n3873);
  and g5818 (n3878, n_3311, n3877);
  not g5819 (n_3315, n3873);
  and g5820 (n3879, n_3312, n_3315);
  not g5821 (n_3316, n3878);
  not g5822 (n_3317, n3879);
  and g5823 (n3880, n_3316, n_3317);
  not g5824 (n_3318, n3876);
  not g5825 (n_3319, n3880);
  and g5826 (n3881, n_3318, n_3319);
  not g5827 (n_3320, n3863);
  not g5828 (n_3321, n3881);
  and g5829 (n3882, n_3320, n_3321);
  not g5830 (n_3322, n3846);
  and g5831 (n3883, n_3322, n3882);
  not g5832 (n_3323, n3882);
  and g5833 (n3884, n3846, n_3323);
  not g5834 (n_3324, n3883);
  not g5835 (n_3325, n3884);
  and g5836 (n3885, n_3324, n_3325);
  not g5837 (n_3327, \A[565] );
  and g5838 (n3886, n_3327, \A[566] );
  not g5839 (n_3329, \A[566] );
  and g5840 (n3887, \A[565] , n_3329);
  not g5841 (n_3331, n3887);
  and g5842 (n3888, \A[567] , n_3331);
  not g5843 (n_3332, n3886);
  and g5844 (n3889, n_3332, n3888);
  and g5845 (n3890, n_3332, n_3331);
  not g5846 (n_3333, \A[567] );
  not g5847 (n_3334, n3890);
  and g5848 (n3891, n_3333, n_3334);
  not g5849 (n_3335, n3889);
  not g5850 (n_3336, n3891);
  and g5851 (n3892, n_3335, n_3336);
  not g5852 (n_3338, \A[568] );
  and g5853 (n3893, n_3338, \A[569] );
  not g5854 (n_3340, \A[569] );
  and g5855 (n3894, \A[568] , n_3340);
  not g5856 (n_3342, n3894);
  and g5857 (n3895, \A[570] , n_3342);
  not g5858 (n_3343, n3893);
  and g5859 (n3896, n_3343, n3895);
  and g5860 (n3897, n_3343, n_3342);
  not g5861 (n_3344, \A[570] );
  not g5862 (n_3345, n3897);
  and g5863 (n3898, n_3344, n_3345);
  not g5864 (n_3346, n3896);
  not g5865 (n_3347, n3898);
  and g5866 (n3899, n_3346, n_3347);
  not g5867 (n_3348, n3892);
  and g5868 (n3900, n_3348, n3899);
  not g5869 (n_3349, n3899);
  and g5870 (n3901, n3892, n_3349);
  not g5871 (n_3350, n3900);
  not g5872 (n_3351, n3901);
  and g5873 (n3902, n_3350, n_3351);
  and g5874 (n3903, \A[568] , \A[569] );
  and g5875 (n3904, \A[570] , n_3345);
  not g5876 (n_3352, n3903);
  not g5877 (n_3353, n3904);
  and g5878 (n3905, n_3352, n_3353);
  and g5879 (n3906, \A[565] , \A[566] );
  and g5880 (n3907, \A[567] , n_3334);
  not g5881 (n_3354, n3906);
  not g5882 (n_3355, n3907);
  and g5883 (n3908, n_3354, n_3355);
  not g5884 (n_3356, n3905);
  and g5885 (n3909, n_3356, n3908);
  not g5886 (n_3357, n3908);
  and g5887 (n3910, n3905, n_3357);
  not g5888 (n_3358, n3909);
  not g5889 (n_3359, n3910);
  and g5890 (n3911, n_3358, n_3359);
  and g5891 (n3912, n_3348, n_3349);
  not g5892 (n_3360, n3911);
  and g5893 (n3913, n_3360, n3912);
  and g5894 (n3914, n_3356, n_3357);
  not g5895 (n_3361, n3913);
  not g5896 (n_3362, n3914);
  and g5897 (n3915, n_3361, n_3362);
  and g5898 (n3916, n_3358, n3912);
  and g5899 (n3917, n_3359, n3916);
  not g5900 (n_3363, n3912);
  and g5901 (n3918, n_3360, n_3363);
  not g5902 (n_3364, n3917);
  not g5903 (n_3365, n3918);
  and g5904 (n3919, n_3364, n_3365);
  not g5905 (n_3366, n3915);
  not g5906 (n_3367, n3919);
  and g5907 (n3920, n_3366, n_3367);
  not g5908 (n_3368, n3902);
  not g5909 (n_3369, n3920);
  and g5910 (n3921, n_3368, n_3369);
  not g5911 (n_3371, \A[559] );
  and g5912 (n3922, n_3371, \A[560] );
  not g5913 (n_3373, \A[560] );
  and g5914 (n3923, \A[559] , n_3373);
  not g5915 (n_3375, n3923);
  and g5916 (n3924, \A[561] , n_3375);
  not g5917 (n_3376, n3922);
  and g5918 (n3925, n_3376, n3924);
  and g5919 (n3926, n_3376, n_3375);
  not g5920 (n_3377, \A[561] );
  not g5921 (n_3378, n3926);
  and g5922 (n3927, n_3377, n_3378);
  not g5923 (n_3379, n3925);
  not g5924 (n_3380, n3927);
  and g5925 (n3928, n_3379, n_3380);
  not g5926 (n_3382, \A[562] );
  and g5927 (n3929, n_3382, \A[563] );
  not g5928 (n_3384, \A[563] );
  and g5929 (n3930, \A[562] , n_3384);
  not g5930 (n_3386, n3930);
  and g5931 (n3931, \A[564] , n_3386);
  not g5932 (n_3387, n3929);
  and g5933 (n3932, n_3387, n3931);
  and g5934 (n3933, n_3387, n_3386);
  not g5935 (n_3388, \A[564] );
  not g5936 (n_3389, n3933);
  and g5937 (n3934, n_3388, n_3389);
  not g5938 (n_3390, n3932);
  not g5939 (n_3391, n3934);
  and g5940 (n3935, n_3390, n_3391);
  not g5941 (n_3392, n3928);
  and g5942 (n3936, n_3392, n3935);
  not g5943 (n_3393, n3935);
  and g5944 (n3937, n3928, n_3393);
  not g5945 (n_3394, n3936);
  not g5946 (n_3395, n3937);
  and g5947 (n3938, n_3394, n_3395);
  and g5948 (n3939, \A[562] , \A[563] );
  and g5949 (n3940, \A[564] , n_3389);
  not g5950 (n_3396, n3939);
  not g5951 (n_3397, n3940);
  and g5952 (n3941, n_3396, n_3397);
  and g5953 (n3942, \A[559] , \A[560] );
  and g5954 (n3943, \A[561] , n_3378);
  not g5955 (n_3398, n3942);
  not g5956 (n_3399, n3943);
  and g5957 (n3944, n_3398, n_3399);
  not g5958 (n_3400, n3941);
  and g5959 (n3945, n_3400, n3944);
  not g5960 (n_3401, n3944);
  and g5961 (n3946, n3941, n_3401);
  not g5962 (n_3402, n3945);
  not g5963 (n_3403, n3946);
  and g5964 (n3947, n_3402, n_3403);
  and g5965 (n3948, n_3392, n_3393);
  not g5966 (n_3404, n3947);
  and g5967 (n3949, n_3404, n3948);
  and g5968 (n3950, n_3400, n_3401);
  not g5969 (n_3405, n3949);
  not g5970 (n_3406, n3950);
  and g5971 (n3951, n_3405, n_3406);
  and g5972 (n3952, n_3402, n3948);
  and g5973 (n3953, n_3403, n3952);
  not g5974 (n_3407, n3948);
  and g5975 (n3954, n_3404, n_3407);
  not g5976 (n_3408, n3953);
  not g5977 (n_3409, n3954);
  and g5978 (n3955, n_3408, n_3409);
  not g5979 (n_3410, n3951);
  not g5980 (n_3411, n3955);
  and g5981 (n3956, n_3410, n_3411);
  not g5982 (n_3412, n3938);
  not g5983 (n_3413, n3956);
  and g5984 (n3957, n_3412, n_3413);
  not g5985 (n_3414, n3921);
  and g5986 (n3958, n_3414, n3957);
  not g5987 (n_3415, n3957);
  and g5988 (n3959, n3921, n_3415);
  not g5989 (n_3416, n3958);
  not g5990 (n_3417, n3959);
  and g5991 (n3960, n_3416, n_3417);
  not g5992 (n_3418, n3885);
  and g5993 (n3961, n_3418, n3960);
  not g5994 (n_3419, n3960);
  and g5995 (n3962, n3885, n_3419);
  not g5996 (n_3420, n3961);
  not g5997 (n_3421, n3962);
  and g5998 (n3963, n_3420, n_3421);
  not g5999 (n_3422, n3810);
  and g6000 (n3964, n_3422, n3963);
  not g6001 (n_3423, n3963);
  and g6002 (n3965, n3810, n_3423);
  not g6003 (n_3424, n3964);
  not g6004 (n_3425, n3965);
  and g6005 (n3966, n_3424, n_3425);
  not g6006 (n_3426, n3657);
  and g6007 (n3967, n_3426, n3966);
  not g6008 (n_3427, n3966);
  and g6009 (n3968, n3657, n_3427);
  not g6010 (n_3428, n3967);
  not g6011 (n_3429, n3968);
  and g6012 (n3969, n_3428, n_3429);
  not g6013 (n_3430, n3348);
  and g6014 (n3970, n_3430, n3969);
  not g6015 (n_3431, n3969);
  and g6016 (n3971, n3348, n_3431);
  not g6017 (n_3432, n3970);
  not g6018 (n_3433, n3971);
  and g6019 (n3972, n_3432, n_3433);
  and g6020 (n3973, n_1889, n2715);
  and g6021 (n3974, n2712, n_1890);
  not g6022 (n_3434, n3973);
  not g6023 (n_3435, n3974);
  and g6024 (n3975, n_3434, n_3435);
  not g6025 (n_3436, n3972);
  not g6026 (n_3437, n3975);
  and g6027 (n3976, n_3436, n_3437);
  not g6028 (n_3438, n2727);
  and g6029 (n3977, n_3438, n3976);
  not g6030 (n_3439, n2722);
  and g6031 (n3978, n_3439, n3977);
  and g6032 (n3979, n_3439, n_3438);
  not g6033 (n_3440, n3976);
  not g6034 (n_3441, n3979);
  and g6035 (n3980, n_3440, n_3441);
  not g6036 (n_3442, n3978);
  not g6037 (n_3443, n3980);
  and g6038 (n3981, n_3442, n_3443);
  and g6039 (n3982, n_3224, n_3222);
  not g6040 (n_3444, n3982);
  and g6041 (n3983, n_3223, n_3444);
  and g6042 (n3984, n_3180, n_3224);
  and g6043 (n3985, n_3181, n3984);
  and g6044 (n3986, n_3225, n3985);
  and g6045 (n3987, n_3180, n_3178);
  not g6046 (n_3445, n3987);
  and g6047 (n3988, n_3179, n_3445);
  not g6048 (n_3446, n3986);
  and g6049 (n3989, n_3446, n3988);
  not g6050 (n_3447, n3988);
  and g6051 (n3990, n3986, n_3447);
  not g6052 (n_3448, n3989);
  not g6053 (n_3449, n3990);
  and g6054 (n3991, n_3448, n_3449);
  not g6055 (n_3450, n3983);
  not g6056 (n_3451, n3991);
  and g6057 (n3992, n_3450, n_3451);
  and g6058 (n3993, n_3446, n_3447);
  not g6063 (n_3452, n3993);
  not g6064 (n_3453, n3997);
  and g6065 (n3998, n_3452, n_3453);
  not g6066 (n_3454, n3998);
  and g6067 (n3999, n3983, n_3454);
  not g6068 (n_3455, n3992);
  not g6069 (n_3456, n3999);
  and g6070 (n4000, n_3455, n_3456);
  and g6071 (n4001, n_3132, n_3130);
  not g6072 (n_3457, n4001);
  and g6073 (n4002, n_3131, n_3457);
  and g6074 (n4003, n_3088, n_3132);
  and g6075 (n4004, n_3089, n4003);
  and g6076 (n4005, n_3133, n4004);
  and g6077 (n4006, n_3088, n_3086);
  not g6078 (n_3458, n4006);
  and g6079 (n4007, n_3087, n_3458);
  not g6080 (n_3459, n4005);
  not g6081 (n_3460, n4007);
  and g6082 (n4008, n_3459, n_3460);
  not g6087 (n_3461, n4008);
  not g6088 (n_3462, n4012);
  and g6089 (n4013, n_3461, n_3462);
  not g6090 (n_3463, n4013);
  and g6091 (n4014, n4002, n_3463);
  and g6092 (n4015, n_3459, n4007);
  and g6093 (n4016, n4005, n_3460);
  not g6094 (n_3464, n4015);
  not g6095 (n_3465, n4016);
  and g6096 (n4017, n_3464, n_3465);
  not g6097 (n_3466, n4002);
  not g6098 (n_3467, n4017);
  and g6099 (n4018, n_3466, n_3467);
  and g6100 (n4019, n_3230, n_3231);
  not g6101 (n_3468, n4018);
  not g6102 (n_3469, n4019);
  and g6103 (n4020, n_3468, n_3469);
  not g6104 (n_3470, n4014);
  and g6105 (n4021, n_3470, n4020);
  and g6106 (n4022, n_3470, n_3468);
  not g6107 (n_3471, n4022);
  and g6108 (n4023, n4019, n_3471);
  not g6109 (n_3472, n4021);
  not g6110 (n_3473, n4023);
  and g6111 (n4024, n_3472, n_3473);
  not g6112 (n_3474, n4000);
  not g6113 (n_3475, n4024);
  and g6114 (n4025, n_3474, n_3475);
  and g6115 (n4026, n_3468, n4019);
  and g6116 (n4027, n_3470, n4026);
  and g6117 (n4028, n_3469, n_3471);
  not g6118 (n_3476, n4027);
  not g6119 (n_3477, n4028);
  and g6120 (n4029, n_3476, n_3477);
  not g6121 (n_3478, n4029);
  and g6122 (n4030, n4000, n_3478);
  and g6123 (n4031, n_3422, n_3423);
  not g6124 (n_3479, n4030);
  and g6125 (n4032, n_3479, n4031);
  not g6126 (n_3480, n4025);
  and g6127 (n4033, n_3480, n4032);
  and g6128 (n4034, n_3480, n_3479);
  not g6129 (n_3481, n4031);
  not g6130 (n_3482, n4034);
  and g6131 (n4035, n_3481, n_3482);
  not g6132 (n_3483, n4033);
  not g6133 (n_3484, n4035);
  and g6134 (n4036, n_3483, n_3484);
  and g6135 (n4037, n_3320, n_3318);
  not g6136 (n_3485, n4037);
  and g6137 (n4038, n_3319, n_3485);
  and g6138 (n4039, n_3276, n_3320);
  and g6139 (n4040, n_3277, n4039);
  and g6140 (n4041, n_3321, n4040);
  and g6141 (n4042, n_3276, n_3274);
  not g6142 (n_3486, n4042);
  and g6143 (n4043, n_3275, n_3486);
  not g6144 (n_3487, n4041);
  not g6145 (n_3488, n4043);
  and g6146 (n4044, n_3487, n_3488);
  not g6151 (n_3489, n4044);
  not g6152 (n_3490, n4048);
  and g6153 (n4049, n_3489, n_3490);
  not g6154 (n_3491, n4049);
  and g6155 (n4050, n4038, n_3491);
  and g6156 (n4051, n_3487, n4043);
  and g6157 (n4052, n4041, n_3488);
  not g6158 (n_3492, n4051);
  not g6159 (n_3493, n4052);
  and g6160 (n4053, n_3492, n_3493);
  not g6161 (n_3494, n4038);
  not g6162 (n_3495, n4053);
  and g6163 (n4054, n_3494, n_3495);
  and g6164 (n4055, n_3418, n_3419);
  not g6165 (n_3496, n4054);
  and g6166 (n4056, n_3496, n4055);
  not g6167 (n_3497, n4050);
  and g6168 (n4057, n_3497, n4056);
  and g6169 (n4058, n_3497, n_3496);
  not g6170 (n_3498, n4055);
  not g6171 (n_3499, n4058);
  and g6172 (n4059, n_3498, n_3499);
  not g6173 (n_3500, n4057);
  not g6174 (n_3501, n4059);
  and g6175 (n4060, n_3500, n_3501);
  and g6176 (n4061, n_3412, n_3410);
  not g6177 (n_3502, n4061);
  and g6178 (n4062, n_3411, n_3502);
  and g6179 (n4063, n_3368, n_3412);
  and g6180 (n4064, n_3369, n4063);
  and g6181 (n4065, n_3413, n4064);
  and g6182 (n4066, n_3368, n_3366);
  not g6183 (n_3503, n4066);
  and g6184 (n4067, n_3367, n_3503);
  not g6185 (n_3504, n4065);
  and g6186 (n4068, n_3504, n4067);
  not g6187 (n_3505, n4067);
  and g6188 (n4069, n4065, n_3505);
  not g6189 (n_3506, n4068);
  not g6190 (n_3507, n4069);
  and g6191 (n4070, n_3506, n_3507);
  not g6192 (n_3508, n4062);
  not g6193 (n_3509, n4070);
  and g6194 (n4071, n_3508, n_3509);
  and g6195 (n4072, n_3504, n_3505);
  not g6200 (n_3510, n4072);
  not g6201 (n_3511, n4076);
  and g6202 (n4077, n_3510, n_3511);
  not g6203 (n_3512, n4077);
  and g6204 (n4078, n4062, n_3512);
  not g6205 (n_3513, n4071);
  not g6206 (n_3514, n4078);
  and g6207 (n4079, n_3513, n_3514);
  not g6208 (n_3515, n4060);
  and g6209 (n4080, n_3515, n4079);
  and g6210 (n4081, n_3496, n_3498);
  and g6211 (n4082, n_3497, n4081);
  and g6212 (n4083, n4055, n_3499);
  not g6213 (n_3516, n4082);
  not g6214 (n_3517, n4083);
  and g6215 (n4084, n_3516, n_3517);
  not g6216 (n_3518, n4079);
  not g6217 (n_3519, n4084);
  and g6218 (n4085, n_3518, n_3519);
  not g6219 (n_3520, n4080);
  not g6220 (n_3521, n4085);
  and g6221 (n4086, n_3520, n_3521);
  not g6222 (n_3522, n4036);
  and g6223 (n4087, n_3522, n4086);
  and g6224 (n4088, n_3479, n_3481);
  and g6225 (n4089, n_3480, n4088);
  and g6226 (n4090, n4031, n_3482);
  not g6227 (n_3523, n4089);
  not g6228 (n_3524, n4090);
  and g6229 (n4091, n_3523, n_3524);
  not g6230 (n_3525, n4086);
  not g6231 (n_3526, n4091);
  and g6232 (n4092, n_3525, n_3526);
  not g6233 (n_3527, n4087);
  not g6234 (n_3528, n4092);
  and g6235 (n4093, n_3527, n_3528);
  and g6236 (n4094, n_2940, n_2938);
  not g6237 (n_3529, n4094);
  and g6238 (n4095, n_2939, n_3529);
  and g6239 (n4096, n_2896, n_2940);
  and g6240 (n4097, n_2897, n4096);
  and g6241 (n4098, n_2941, n4097);
  and g6242 (n4099, n_2896, n_2894);
  not g6243 (n_3530, n4099);
  and g6244 (n4100, n_2895, n_3530);
  not g6245 (n_3531, n4098);
  not g6246 (n_3532, n4100);
  and g6247 (n4101, n_3531, n_3532);
  not g6252 (n_3533, n4101);
  not g6253 (n_3534, n4105);
  and g6254 (n4106, n_3533, n_3534);
  not g6255 (n_3535, n4106);
  and g6256 (n4107, n4095, n_3535);
  and g6257 (n4108, n_3531, n4100);
  and g6258 (n4109, n4098, n_3532);
  not g6259 (n_3536, n4108);
  not g6260 (n_3537, n4109);
  and g6261 (n4110, n_3536, n_3537);
  not g6262 (n_3538, n4095);
  not g6263 (n_3539, n4110);
  and g6264 (n4111, n_3538, n_3539);
  and g6265 (n4112, n_3038, n_3039);
  not g6266 (n_3540, n4111);
  and g6267 (n4113, n_3540, n4112);
  not g6268 (n_3541, n4107);
  and g6269 (n4114, n_3541, n4113);
  and g6270 (n4115, n_3541, n_3540);
  not g6271 (n_3542, n4112);
  not g6272 (n_3543, n4115);
  and g6273 (n4116, n_3542, n_3543);
  not g6274 (n_3544, n4114);
  not g6275 (n_3545, n4116);
  and g6276 (n4117, n_3544, n_3545);
  and g6277 (n4118, n_3032, n_3030);
  not g6278 (n_3546, n4118);
  and g6279 (n4119, n_3031, n_3546);
  and g6280 (n4120, n_2988, n_3032);
  and g6281 (n4121, n_2989, n4120);
  and g6282 (n4122, n_3033, n4121);
  and g6283 (n4123, n_2988, n_2986);
  not g6284 (n_3547, n4123);
  and g6285 (n4124, n_2987, n_3547);
  not g6286 (n_3548, n4122);
  and g6287 (n4125, n_3548, n4124);
  not g6288 (n_3549, n4124);
  and g6289 (n4126, n4122, n_3549);
  not g6290 (n_3550, n4125);
  not g6291 (n_3551, n4126);
  and g6292 (n4127, n_3550, n_3551);
  not g6293 (n_3552, n4119);
  not g6294 (n_3553, n4127);
  and g6295 (n4128, n_3552, n_3553);
  and g6296 (n4129, n_3548, n_3549);
  not g6301 (n_3554, n4129);
  not g6302 (n_3555, n4133);
  and g6303 (n4134, n_3554, n_3555);
  not g6304 (n_3556, n4134);
  and g6305 (n4135, n4119, n_3556);
  not g6306 (n_3557, n4128);
  not g6307 (n_3558, n4135);
  and g6308 (n4136, n_3557, n_3558);
  not g6309 (n_3559, n4117);
  and g6310 (n4137, n_3559, n4136);
  and g6311 (n4138, n_3540, n_3542);
  and g6312 (n4139, n_3541, n4138);
  and g6313 (n4140, n4112, n_3543);
  not g6314 (n_3560, n4139);
  not g6315 (n_3561, n4140);
  and g6316 (n4141, n_3560, n_3561);
  not g6317 (n_3562, n4136);
  not g6318 (n_3563, n4141);
  and g6319 (n4142, n_3562, n_3563);
  not g6320 (n_3564, n4137);
  not g6321 (n_3565, n4142);
  and g6322 (n4143, n_3564, n_3565);
  and g6323 (n4144, n_2844, n_2842);
  not g6324 (n_3566, n4144);
  and g6325 (n4145, n_2843, n_3566);
  and g6326 (n4146, n_2800, n_2844);
  and g6327 (n4147, n_2801, n4146);
  and g6328 (n4148, n_2845, n4147);
  and g6329 (n4149, n_2800, n_2798);
  not g6330 (n_3567, n4149);
  and g6331 (n4150, n_2799, n_3567);
  not g6332 (n_3568, n4148);
  and g6333 (n4151, n_3568, n4150);
  not g6334 (n_3569, n4150);
  and g6335 (n4152, n4148, n_3569);
  not g6336 (n_3570, n4151);
  not g6337 (n_3571, n4152);
  and g6338 (n4153, n_3570, n_3571);
  not g6339 (n_3572, n4145);
  not g6340 (n_3573, n4153);
  and g6341 (n4154, n_3572, n_3573);
  and g6342 (n4155, n_3568, n_3569);
  not g6347 (n_3574, n4155);
  not g6348 (n_3575, n4159);
  and g6349 (n4160, n_3574, n_3575);
  not g6350 (n_3576, n4160);
  and g6351 (n4161, n4145, n_3576);
  not g6352 (n_3577, n4154);
  not g6353 (n_3578, n4161);
  and g6354 (n4162, n_3577, n_3578);
  and g6355 (n4163, n_2752, n_2750);
  not g6356 (n_3579, n4163);
  and g6357 (n4164, n_2751, n_3579);
  and g6358 (n4165, n_2708, n_2752);
  and g6359 (n4166, n_2709, n4165);
  and g6360 (n4167, n_2753, n4166);
  and g6361 (n4168, n_2708, n_2706);
  not g6362 (n_3580, n4168);
  and g6363 (n4169, n_2707, n_3580);
  not g6364 (n_3581, n4167);
  not g6365 (n_3582, n4169);
  and g6366 (n4170, n_3581, n_3582);
  not g6371 (n_3583, n4170);
  not g6372 (n_3584, n4174);
  and g6373 (n4175, n_3583, n_3584);
  not g6374 (n_3585, n4175);
  and g6375 (n4176, n4164, n_3585);
  and g6376 (n4177, n_3581, n4169);
  and g6377 (n4178, n4167, n_3582);
  not g6378 (n_3586, n4177);
  not g6379 (n_3587, n4178);
  and g6380 (n4179, n_3586, n_3587);
  not g6381 (n_3588, n4164);
  not g6382 (n_3589, n4179);
  and g6383 (n4180, n_3588, n_3589);
  and g6384 (n4181, n_2850, n_2851);
  not g6385 (n_3590, n4180);
  not g6386 (n_3591, n4181);
  and g6387 (n4182, n_3590, n_3591);
  not g6388 (n_3592, n4176);
  and g6389 (n4183, n_3592, n4182);
  and g6390 (n4184, n_3592, n_3590);
  not g6391 (n_3593, n4184);
  and g6392 (n4185, n4181, n_3593);
  not g6393 (n_3594, n4183);
  not g6394 (n_3595, n4185);
  and g6395 (n4186, n_3594, n_3595);
  not g6396 (n_3596, n4162);
  not g6397 (n_3597, n4186);
  and g6398 (n4187, n_3596, n_3597);
  and g6399 (n4188, n_3590, n4181);
  and g6400 (n4189, n_3592, n4188);
  and g6401 (n4190, n_3591, n_3593);
  not g6402 (n_3598, n4189);
  not g6403 (n_3599, n4190);
  and g6404 (n4191, n_3598, n_3599);
  not g6405 (n_3600, n4191);
  and g6406 (n4192, n4162, n_3600);
  and g6407 (n4193, n_3042, n_3043);
  not g6408 (n_3601, n4192);
  not g6409 (n_3602, n4193);
  and g6410 (n4194, n_3601, n_3602);
  not g6411 (n_3603, n4187);
  and g6412 (n4195, n_3603, n4194);
  and g6413 (n4196, n_3603, n_3601);
  not g6414 (n_3604, n4196);
  and g6415 (n4197, n4193, n_3604);
  not g6416 (n_3605, n4195);
  not g6417 (n_3606, n4197);
  and g6418 (n4198, n_3605, n_3606);
  not g6419 (n_3607, n4143);
  not g6420 (n_3608, n4198);
  and g6421 (n4199, n_3607, n_3608);
  and g6422 (n4200, n_3601, n4193);
  and g6423 (n4201, n_3603, n4200);
  and g6424 (n4202, n_3602, n_3604);
  not g6425 (n_3609, n4201);
  not g6426 (n_3610, n4202);
  and g6427 (n4203, n_3609, n_3610);
  not g6428 (n_3611, n4203);
  and g6429 (n4204, n4143, n_3611);
  and g6430 (n4205, n_3426, n_3427);
  not g6431 (n_3612, n4204);
  not g6432 (n_3613, n4205);
  and g6433 (n4206, n_3612, n_3613);
  not g6434 (n_3614, n4199);
  and g6435 (n4207, n_3614, n4206);
  and g6436 (n4208, n_3614, n_3612);
  not g6437 (n_3615, n4208);
  and g6438 (n4209, n4205, n_3615);
  not g6439 (n_3616, n4207);
  not g6440 (n_3617, n4209);
  and g6441 (n4210, n_3616, n_3617);
  not g6442 (n_3618, n4093);
  not g6443 (n_3619, n4210);
  and g6444 (n4211, n_3618, n_3619);
  and g6445 (n4212, n_3612, n4205);
  and g6446 (n4213, n_3614, n4212);
  and g6447 (n4214, n_3613, n_3615);
  not g6448 (n_3620, n4213);
  not g6449 (n_3621, n4214);
  and g6450 (n4215, n_3620, n_3621);
  not g6451 (n_3622, n4215);
  and g6452 (n4216, n4093, n_3622);
  and g6453 (n4217, n_3430, n_3431);
  not g6454 (n_3623, n4216);
  and g6455 (n4218, n_3623, n4217);
  not g6456 (n_3624, n4211);
  and g6457 (n4219, n_3624, n4218);
  and g6458 (n4220, n_3624, n_3623);
  not g6459 (n_3625, n4217);
  not g6460 (n_3626, n4220);
  and g6461 (n4221, n_3625, n_3626);
  not g6462 (n_3627, n4219);
  not g6463 (n_3628, n4221);
  and g6464 (n4222, n_3627, n_3628);
  and g6465 (n4223, n_2556, n_2554);
  not g6466 (n_3629, n4223);
  and g6467 (n4224, n_2555, n_3629);
  and g6468 (n4225, n_2512, n_2556);
  and g6469 (n4226, n_2513, n4225);
  and g6470 (n4227, n_2557, n4226);
  and g6471 (n4228, n_2512, n_2510);
  not g6472 (n_3630, n4228);
  and g6473 (n4229, n_2511, n_3630);
  not g6474 (n_3631, n4227);
  not g6475 (n_3632, n4229);
  and g6476 (n4230, n_3631, n_3632);
  not g6481 (n_3633, n4230);
  not g6482 (n_3634, n4234);
  and g6483 (n4235, n_3633, n_3634);
  not g6484 (n_3635, n4235);
  and g6485 (n4236, n4224, n_3635);
  and g6486 (n4237, n_3631, n4229);
  and g6487 (n4238, n4227, n_3632);
  not g6488 (n_3636, n4237);
  not g6489 (n_3637, n4238);
  and g6490 (n4239, n_3636, n_3637);
  not g6491 (n_3638, n4224);
  not g6492 (n_3639, n4239);
  and g6493 (n4240, n_3638, n_3639);
  and g6494 (n4241, n_2654, n_2655);
  not g6495 (n_3640, n4240);
  and g6496 (n4242, n_3640, n4241);
  not g6497 (n_3641, n4236);
  and g6498 (n4243, n_3641, n4242);
  and g6499 (n4244, n_3641, n_3640);
  not g6500 (n_3642, n4241);
  not g6501 (n_3643, n4244);
  and g6502 (n4245, n_3642, n_3643);
  not g6503 (n_3644, n4243);
  not g6504 (n_3645, n4245);
  and g6505 (n4246, n_3644, n_3645);
  and g6506 (n4247, n_2648, n_2646);
  not g6507 (n_3646, n4247);
  and g6508 (n4248, n_2647, n_3646);
  and g6509 (n4249, n_2604, n_2648);
  and g6510 (n4250, n_2605, n4249);
  and g6511 (n4251, n_2649, n4250);
  and g6512 (n4252, n_2604, n_2602);
  not g6513 (n_3647, n4252);
  and g6514 (n4253, n_2603, n_3647);
  not g6515 (n_3648, n4251);
  and g6516 (n4254, n_3648, n4253);
  not g6517 (n_3649, n4253);
  and g6518 (n4255, n4251, n_3649);
  not g6519 (n_3650, n4254);
  not g6520 (n_3651, n4255);
  and g6521 (n4256, n_3650, n_3651);
  not g6522 (n_3652, n4248);
  not g6523 (n_3653, n4256);
  and g6524 (n4257, n_3652, n_3653);
  and g6525 (n4258, n_3648, n_3649);
  not g6530 (n_3654, n4258);
  not g6531 (n_3655, n4262);
  and g6532 (n4263, n_3654, n_3655);
  not g6533 (n_3656, n4263);
  and g6534 (n4264, n4248, n_3656);
  not g6535 (n_3657, n4257);
  not g6536 (n_3658, n4264);
  and g6537 (n4265, n_3657, n_3658);
  not g6538 (n_3659, n4246);
  and g6539 (n4266, n_3659, n4265);
  and g6540 (n4267, n_3640, n_3642);
  and g6541 (n4268, n_3641, n4267);
  and g6542 (n4269, n4241, n_3643);
  not g6543 (n_3660, n4268);
  not g6544 (n_3661, n4269);
  and g6545 (n4270, n_3660, n_3661);
  not g6546 (n_3662, n4265);
  not g6547 (n_3663, n4270);
  and g6548 (n4271, n_3662, n_3663);
  not g6549 (n_3664, n4266);
  not g6550 (n_3665, n4271);
  and g6551 (n4272, n_3664, n_3665);
  and g6552 (n4273, n_2460, n_2458);
  not g6553 (n_3666, n4273);
  and g6554 (n4274, n_2459, n_3666);
  and g6555 (n4275, n_2416, n_2460);
  and g6556 (n4276, n_2417, n4275);
  and g6557 (n4277, n_2461, n4276);
  and g6558 (n4278, n_2416, n_2414);
  not g6559 (n_3667, n4278);
  and g6560 (n4279, n_2415, n_3667);
  not g6561 (n_3668, n4277);
  and g6562 (n4280, n_3668, n4279);
  not g6563 (n_3669, n4279);
  and g6564 (n4281, n4277, n_3669);
  not g6565 (n_3670, n4280);
  not g6566 (n_3671, n4281);
  and g6567 (n4282, n_3670, n_3671);
  not g6568 (n_3672, n4274);
  not g6569 (n_3673, n4282);
  and g6570 (n4283, n_3672, n_3673);
  and g6571 (n4284, n_3668, n_3669);
  not g6576 (n_3674, n4284);
  not g6577 (n_3675, n4288);
  and g6578 (n4289, n_3674, n_3675);
  not g6579 (n_3676, n4289);
  and g6580 (n4290, n4274, n_3676);
  not g6581 (n_3677, n4283);
  not g6582 (n_3678, n4290);
  and g6583 (n4291, n_3677, n_3678);
  and g6584 (n4292, n_2368, n_2366);
  not g6585 (n_3679, n4292);
  and g6586 (n4293, n_2367, n_3679);
  and g6587 (n4294, n_2324, n_2368);
  and g6588 (n4295, n_2325, n4294);
  and g6589 (n4296, n_2369, n4295);
  and g6590 (n4297, n_2324, n_2322);
  not g6591 (n_3680, n4297);
  and g6592 (n4298, n_2323, n_3680);
  not g6593 (n_3681, n4296);
  not g6594 (n_3682, n4298);
  and g6595 (n4299, n_3681, n_3682);
  not g6600 (n_3683, n4299);
  not g6601 (n_3684, n4303);
  and g6602 (n4304, n_3683, n_3684);
  not g6603 (n_3685, n4304);
  and g6604 (n4305, n4293, n_3685);
  and g6605 (n4306, n_3681, n4298);
  and g6606 (n4307, n4296, n_3682);
  not g6607 (n_3686, n4306);
  not g6608 (n_3687, n4307);
  and g6609 (n4308, n_3686, n_3687);
  not g6610 (n_3688, n4293);
  not g6611 (n_3689, n4308);
  and g6612 (n4309, n_3688, n_3689);
  and g6613 (n4310, n_2466, n_2467);
  not g6614 (n_3690, n4309);
  not g6615 (n_3691, n4310);
  and g6616 (n4311, n_3690, n_3691);
  not g6617 (n_3692, n4305);
  and g6618 (n4312, n_3692, n4311);
  and g6619 (n4313, n_3692, n_3690);
  not g6620 (n_3693, n4313);
  and g6621 (n4314, n4310, n_3693);
  not g6622 (n_3694, n4312);
  not g6623 (n_3695, n4314);
  and g6624 (n4315, n_3694, n_3695);
  not g6625 (n_3696, n4291);
  not g6626 (n_3697, n4315);
  and g6627 (n4316, n_3696, n_3697);
  and g6628 (n4317, n_3690, n4310);
  and g6629 (n4318, n_3692, n4317);
  and g6630 (n4319, n_3691, n_3693);
  not g6631 (n_3698, n4318);
  not g6632 (n_3699, n4319);
  and g6633 (n4320, n_3698, n_3699);
  not g6634 (n_3700, n4320);
  and g6635 (n4321, n4291, n_3700);
  and g6636 (n4322, n_2658, n_2659);
  not g6637 (n_3701, n4321);
  not g6638 (n_3702, n4322);
  and g6639 (n4323, n_3701, n_3702);
  not g6640 (n_3703, n4316);
  and g6641 (n4324, n_3703, n4323);
  and g6642 (n4325, n_3703, n_3701);
  not g6643 (n_3704, n4325);
  and g6644 (n4326, n4322, n_3704);
  not g6645 (n_3705, n4324);
  not g6646 (n_3706, n4326);
  and g6647 (n4327, n_3705, n_3706);
  not g6648 (n_3707, n4272);
  not g6649 (n_3708, n4327);
  and g6650 (n4328, n_3707, n_3708);
  and g6651 (n4329, n_3701, n4322);
  and g6652 (n4330, n_3703, n4329);
  and g6653 (n4331, n_3702, n_3704);
  not g6654 (n_3709, n4330);
  not g6655 (n_3710, n4331);
  and g6656 (n4332, n_3709, n_3710);
  not g6657 (n_3711, n4332);
  and g6658 (n4333, n4272, n_3711);
  and g6659 (n4334, n_2662, n_2663);
  not g6660 (n_3712, n4333);
  and g6661 (n4335, n_3712, n4334);
  not g6662 (n_3713, n4328);
  and g6663 (n4336, n_3713, n4335);
  and g6664 (n4337, n_3713, n_3712);
  not g6665 (n_3714, n4334);
  not g6666 (n_3715, n4337);
  and g6667 (n4338, n_3714, n_3715);
  not g6668 (n_3716, n4336);
  not g6669 (n_3717, n4338);
  and g6670 (n4339, n_3716, n_3717);
  and g6671 (n4340, n_2268, n_2266);
  not g6672 (n_3718, n4340);
  and g6673 (n4341, n_2267, n_3718);
  and g6674 (n4342, n_2224, n_2268);
  and g6675 (n4343, n_2225, n4342);
  and g6676 (n4344, n_2269, n4343);
  and g6677 (n4345, n_2224, n_2222);
  not g6678 (n_3719, n4345);
  and g6679 (n4346, n_2223, n_3719);
  not g6680 (n_3720, n4344);
  and g6681 (n4347, n_3720, n4346);
  not g6682 (n_3721, n4346);
  and g6683 (n4348, n4344, n_3721);
  not g6684 (n_3722, n4347);
  not g6685 (n_3723, n4348);
  and g6686 (n4349, n_3722, n_3723);
  not g6687 (n_3724, n4341);
  not g6688 (n_3725, n4349);
  and g6689 (n4350, n_3724, n_3725);
  and g6690 (n4351, n_3720, n_3721);
  not g6695 (n_3726, n4351);
  not g6696 (n_3727, n4355);
  and g6697 (n4356, n_3726, n_3727);
  not g6698 (n_3728, n4356);
  and g6699 (n4357, n4341, n_3728);
  not g6700 (n_3729, n4350);
  not g6701 (n_3730, n4357);
  and g6702 (n4358, n_3729, n_3730);
  and g6703 (n4359, n_2176, n_2174);
  not g6704 (n_3731, n4359);
  and g6705 (n4360, n_2175, n_3731);
  and g6706 (n4361, n_2132, n_2176);
  and g6707 (n4362, n_2133, n4361);
  and g6708 (n4363, n_2177, n4362);
  and g6709 (n4364, n_2132, n_2130);
  not g6710 (n_3732, n4364);
  and g6711 (n4365, n_2131, n_3732);
  not g6712 (n_3733, n4363);
  not g6713 (n_3734, n4365);
  and g6714 (n4366, n_3733, n_3734);
  not g6719 (n_3735, n4366);
  not g6720 (n_3736, n4370);
  and g6721 (n4371, n_3735, n_3736);
  not g6722 (n_3737, n4371);
  and g6723 (n4372, n4360, n_3737);
  and g6724 (n4373, n_3733, n4365);
  and g6725 (n4374, n4363, n_3734);
  not g6726 (n_3738, n4373);
  not g6727 (n_3739, n4374);
  and g6728 (n4375, n_3738, n_3739);
  not g6729 (n_3740, n4360);
  not g6730 (n_3741, n4375);
  and g6731 (n4376, n_3740, n_3741);
  and g6732 (n4377, n_2274, n_2275);
  not g6733 (n_3742, n4376);
  not g6734 (n_3743, n4377);
  and g6735 (n4378, n_3742, n_3743);
  not g6736 (n_3744, n4372);
  and g6737 (n4379, n_3744, n4378);
  and g6738 (n4380, n_3744, n_3742);
  not g6739 (n_3745, n4380);
  and g6740 (n4381, n4377, n_3745);
  not g6741 (n_3746, n4379);
  not g6742 (n_3747, n4381);
  and g6743 (n4382, n_3746, n_3747);
  not g6744 (n_3748, n4358);
  not g6745 (n_3749, n4382);
  and g6746 (n4383, n_3748, n_3749);
  and g6747 (n4384, n_3742, n4377);
  and g6748 (n4385, n_3744, n4384);
  and g6749 (n4386, n_3743, n_3745);
  not g6750 (n_3750, n4385);
  not g6751 (n_3751, n4386);
  and g6752 (n4387, n_3750, n_3751);
  not g6753 (n_3752, n4387);
  and g6754 (n4388, n4358, n_3752);
  and g6755 (n4389, n_2278, n_2279);
  not g6756 (n_3753, n4388);
  and g6757 (n4390, n_3753, n4389);
  not g6758 (n_3754, n4383);
  and g6759 (n4391, n_3754, n4390);
  and g6760 (n4392, n_3754, n_3753);
  not g6761 (n_3755, n4389);
  not g6762 (n_3756, n4392);
  and g6763 (n4393, n_3755, n_3756);
  not g6764 (n_3757, n4391);
  not g6765 (n_3758, n4393);
  and g6766 (n4394, n_3757, n_3758);
  and g6767 (n4395, n_2080, n_2078);
  not g6768 (n_3759, n4395);
  and g6769 (n4396, n_2079, n_3759);
  and g6770 (n4397, n_2036, n_2080);
  and g6771 (n4398, n_2037, n4397);
  and g6772 (n4399, n_2081, n4398);
  and g6773 (n4400, n_2036, n_2034);
  not g6774 (n_3760, n4400);
  and g6775 (n4401, n_2035, n_3760);
  not g6776 (n_3761, n4399);
  not g6777 (n_3762, n4401);
  and g6778 (n4402, n_3761, n_3762);
  not g6783 (n_3763, n4402);
  not g6784 (n_3764, n4406);
  and g6785 (n4407, n_3763, n_3764);
  not g6786 (n_3765, n4407);
  and g6787 (n4408, n4396, n_3765);
  and g6788 (n4409, n_3761, n4401);
  and g6789 (n4410, n4399, n_3762);
  not g6790 (n_3766, n4409);
  not g6791 (n_3767, n4410);
  and g6792 (n4411, n_3766, n_3767);
  not g6793 (n_3768, n4396);
  not g6794 (n_3769, n4411);
  and g6795 (n4412, n_3768, n_3769);
  and g6796 (n4413, n_2086, n_2087);
  not g6797 (n_3770, n4412);
  and g6798 (n4414, n_3770, n4413);
  not g6799 (n_3771, n4408);
  and g6800 (n4415, n_3771, n4414);
  and g6801 (n4416, n_3771, n_3770);
  not g6802 (n_3772, n4413);
  not g6803 (n_3773, n4416);
  and g6804 (n4417, n_3772, n_3773);
  not g6805 (n_3774, n4415);
  not g6806 (n_3775, n4417);
  and g6807 (n4418, n_3774, n_3775);
  and g6808 (n4419, n_1988, n_1987);
  not g6809 (n_3776, n4419);
  and g6810 (n4420, n_1986, n_3776);
  and g6811 (n4421, n_1944, n_1988);
  and g6812 (n4422, n_1945, n4421);
  and g6813 (n4423, n_1989, n4422);
  and g6814 (n4424, n_1944, n_1942);
  not g6815 (n_3777, n4424);
  and g6816 (n4425, n_1943, n_3777);
  not g6817 (n_3778, n4423);
  and g6818 (n4426, n_3778, n4425);
  not g6819 (n_3779, n4425);
  and g6820 (n4427, n4423, n_3779);
  not g6821 (n_3780, n4426);
  not g6822 (n_3781, n4427);
  and g6823 (n4428, n_3780, n_3781);
  not g6824 (n_3782, n4420);
  not g6825 (n_3783, n4428);
  and g6826 (n4429, n_3782, n_3783);
  and g6827 (n4430, n_3778, n_3779);
  not g6832 (n_3784, n4430);
  not g6833 (n_3785, n4434);
  and g6834 (n4435, n_3784, n_3785);
  not g6835 (n_3786, n4435);
  and g6836 (n4436, n4420, n_3786);
  not g6837 (n_3787, n4429);
  not g6838 (n_3788, n4436);
  and g6839 (n4437, n_3787, n_3788);
  not g6840 (n_3789, n4418);
  and g6841 (n4438, n_3789, n4437);
  and g6842 (n4439, n_3770, n_3772);
  and g6843 (n4440, n_3771, n4439);
  and g6844 (n4441, n4413, n_3773);
  not g6845 (n_3790, n4440);
  not g6846 (n_3791, n4441);
  and g6847 (n4442, n_3790, n_3791);
  not g6848 (n_3792, n4437);
  not g6849 (n_3793, n4442);
  and g6850 (n4443, n_3792, n_3793);
  not g6851 (n_3794, n4438);
  not g6852 (n_3795, n4443);
  and g6853 (n4444, n_3794, n_3795);
  not g6854 (n_3796, n4394);
  and g6855 (n4445, n_3796, n4444);
  and g6856 (n4446, n_3753, n_3755);
  and g6857 (n4447, n_3754, n4446);
  and g6858 (n4448, n4389, n_3756);
  not g6859 (n_3797, n4447);
  not g6860 (n_3798, n4448);
  and g6861 (n4449, n_3797, n_3798);
  not g6862 (n_3799, n4444);
  not g6863 (n_3800, n4449);
  and g6864 (n4450, n_3799, n_3800);
  not g6865 (n_3801, n4445);
  not g6866 (n_3802, n4450);
  and g6867 (n4451, n_3801, n_3802);
  not g6868 (n_3803, n4339);
  and g6869 (n4452, n_3803, n4451);
  and g6870 (n4453, n_3712, n_3714);
  and g6871 (n4454, n_3713, n4453);
  and g6872 (n4455, n4334, n_3715);
  not g6873 (n_3804, n4454);
  not g6874 (n_3805, n4455);
  and g6875 (n4456, n_3804, n_3805);
  not g6876 (n_3806, n4451);
  not g6877 (n_3807, n4456);
  and g6878 (n4457, n_3806, n_3807);
  not g6879 (n_3808, n4452);
  not g6880 (n_3809, n4457);
  and g6881 (n4458, n_3808, n_3809);
  not g6882 (n_3810, n4222);
  and g6883 (n4459, n_3810, n4458);
  and g6884 (n4460, n_3623, n_3625);
  and g6885 (n4461, n_3624, n4460);
  and g6886 (n4462, n4217, n_3626);
  not g6887 (n_3811, n4461);
  not g6888 (n_3812, n4462);
  and g6889 (n4463, n_3811, n_3812);
  not g6890 (n_3813, n4458);
  not g6891 (n_3814, n4463);
  and g6892 (n4464, n_3813, n_3814);
  not g6893 (n_3815, n4459);
  not g6894 (n_3816, n4464);
  and g6895 (n4465, n_3815, n_3816);
  not g6896 (n_3817, n3981);
  and g6897 (n4466, n_3817, n4465);
  and g6898 (n4467, n_3438, n_3440);
  and g6899 (n4468, n_3439, n4467);
  and g6900 (n4469, n3976, n_3441);
  not g6901 (n_3818, n4468);
  not g6902 (n_3819, n4469);
  and g6903 (n4470, n_3818, n_3819);
  not g6904 (n_3820, n4465);
  not g6905 (n_3821, n4470);
  and g6906 (n4471, n_3820, n_3821);
  not g6907 (n_3822, n4466);
  not g6908 (n_3823, n4471);
  and g6909 (n4472, n_3822, n_3823);
  and g6910 (n4473, \A[970] , \A[971] );
  not g6911 (n_3826, \A[971] );
  and g6912 (n4474, \A[970] , n_3826);
  not g6913 (n_3827, \A[970] );
  and g6914 (n4475, n_3827, \A[971] );
  not g6915 (n_3828, n4474);
  not g6916 (n_3829, n4475);
  and g6917 (n4476, n_3828, n_3829);
  not g6918 (n_3831, n4476);
  and g6919 (n4477, \A[972] , n_3831);
  not g6920 (n_3832, n4473);
  not g6921 (n_3833, n4477);
  and g6922 (n4478, n_3832, n_3833);
  and g6923 (n4479, \A[967] , \A[968] );
  not g6924 (n_3836, \A[968] );
  and g6925 (n4480, \A[967] , n_3836);
  not g6926 (n_3837, \A[967] );
  and g6927 (n4481, n_3837, \A[968] );
  not g6928 (n_3838, n4480);
  not g6929 (n_3839, n4481);
  and g6930 (n4482, n_3838, n_3839);
  not g6931 (n_3841, n4482);
  and g6932 (n4483, \A[969] , n_3841);
  not g6933 (n_3842, n4479);
  not g6934 (n_3843, n4483);
  and g6935 (n4484, n_3842, n_3843);
  not g6936 (n_3844, n4484);
  and g6937 (n4485, n4478, n_3844);
  not g6938 (n_3845, n4478);
  and g6939 (n4486, n_3845, n4484);
  and g6940 (n4487, \A[969] , n_3838);
  and g6941 (n4488, n_3839, n4487);
  not g6942 (n_3846, \A[969] );
  and g6943 (n4489, n_3846, n_3841);
  not g6944 (n_3847, n4488);
  not g6945 (n_3848, n4489);
  and g6946 (n4490, n_3847, n_3848);
  and g6947 (n4491, \A[972] , n_3828);
  and g6948 (n4492, n_3829, n4491);
  not g6949 (n_3849, \A[972] );
  and g6950 (n4493, n_3849, n_3831);
  not g6951 (n_3850, n4492);
  not g6952 (n_3851, n4493);
  and g6953 (n4494, n_3850, n_3851);
  not g6954 (n_3852, n4490);
  not g6955 (n_3853, n4494);
  and g6956 (n4495, n_3852, n_3853);
  not g6957 (n_3854, n4486);
  and g6958 (n4496, n_3854, n4495);
  not g6959 (n_3855, n4485);
  and g6960 (n4497, n_3855, n4496);
  and g6961 (n4498, n_3855, n_3854);
  not g6962 (n_3856, n4495);
  not g6963 (n_3857, n4498);
  and g6964 (n4499, n_3856, n_3857);
  not g6965 (n_3858, n4497);
  not g6966 (n_3859, n4499);
  and g6967 (n4500, n_3858, n_3859);
  and g6968 (n4501, n_3852, n4494);
  and g6969 (n4502, n4490, n_3853);
  not g6970 (n_3860, n4501);
  not g6971 (n_3861, n4502);
  and g6972 (n4503, n_3860, n_3861);
  and g6973 (n4504, n4495, n_3857);
  and g6974 (n4505, n_3845, n_3844);
  not g6975 (n_3862, n4504);
  not g6976 (n_3863, n4505);
  and g6977 (n4506, n_3862, n_3863);
  not g6978 (n_3864, n4503);
  not g6979 (n_3865, n4506);
  and g6980 (n4507, n_3864, n_3865);
  not g6981 (n_3866, n4500);
  not g6982 (n_3867, n4507);
  and g6983 (n4508, n_3866, n_3867);
  and g6984 (n4509, n_3866, n_3865);
  and g6985 (n4510, \A[976] , \A[977] );
  not g6986 (n_3870, \A[977] );
  and g6987 (n4511, \A[976] , n_3870);
  not g6988 (n_3871, \A[976] );
  and g6989 (n4512, n_3871, \A[977] );
  not g6990 (n_3872, n4511);
  not g6991 (n_3873, n4512);
  and g6992 (n4513, n_3872, n_3873);
  not g6993 (n_3875, n4513);
  and g6994 (n4514, \A[978] , n_3875);
  not g6995 (n_3876, n4510);
  not g6996 (n_3877, n4514);
  and g6997 (n4515, n_3876, n_3877);
  and g6998 (n4516, \A[973] , \A[974] );
  not g6999 (n_3880, \A[974] );
  and g7000 (n4517, \A[973] , n_3880);
  not g7001 (n_3881, \A[973] );
  and g7002 (n4518, n_3881, \A[974] );
  not g7003 (n_3882, n4517);
  not g7004 (n_3883, n4518);
  and g7005 (n4519, n_3882, n_3883);
  not g7006 (n_3885, n4519);
  and g7007 (n4520, \A[975] , n_3885);
  not g7008 (n_3886, n4516);
  not g7009 (n_3887, n4520);
  and g7010 (n4521, n_3886, n_3887);
  not g7011 (n_3888, n4515);
  and g7012 (n4522, n_3888, n4521);
  not g7013 (n_3889, n4521);
  and g7014 (n4523, n4515, n_3889);
  not g7015 (n_3890, n4522);
  not g7016 (n_3891, n4523);
  and g7017 (n4524, n_3890, n_3891);
  and g7018 (n4525, \A[975] , n_3882);
  and g7019 (n4526, n_3883, n4525);
  not g7020 (n_3892, \A[975] );
  and g7021 (n4527, n_3892, n_3885);
  not g7022 (n_3893, n4526);
  not g7023 (n_3894, n4527);
  and g7024 (n4528, n_3893, n_3894);
  and g7025 (n4529, \A[978] , n_3872);
  and g7026 (n4530, n_3873, n4529);
  not g7027 (n_3895, \A[978] );
  and g7028 (n4531, n_3895, n_3875);
  not g7029 (n_3896, n4530);
  not g7030 (n_3897, n4531);
  and g7031 (n4532, n_3896, n_3897);
  not g7032 (n_3898, n4528);
  not g7033 (n_3899, n4532);
  and g7034 (n4533, n_3898, n_3899);
  not g7035 (n_3900, n4524);
  and g7036 (n4534, n_3900, n4533);
  and g7037 (n4535, n_3888, n_3889);
  not g7038 (n_3901, n4534);
  not g7039 (n_3902, n4535);
  and g7040 (n4536, n_3901, n_3902);
  and g7041 (n4537, n_3890, n4533);
  and g7042 (n4538, n_3891, n4537);
  not g7043 (n_3903, n4533);
  and g7044 (n4539, n_3900, n_3903);
  not g7045 (n_3904, n4538);
  not g7046 (n_3905, n4539);
  and g7047 (n4540, n_3904, n_3905);
  not g7048 (n_3906, n4536);
  not g7049 (n_3907, n4540);
  and g7050 (n4541, n_3906, n_3907);
  and g7051 (n4542, n_3898, n4532);
  and g7052 (n4543, n4528, n_3899);
  not g7053 (n_3908, n4542);
  not g7054 (n_3909, n4543);
  and g7055 (n4544, n_3908, n_3909);
  not g7056 (n_3910, n4544);
  and g7057 (n4545, n_3864, n_3910);
  not g7058 (n_3911, n4541);
  and g7059 (n4546, n_3911, n4545);
  not g7060 (n_3912, n4509);
  and g7061 (n4547, n_3912, n4546);
  and g7062 (n4548, n_3906, n_3910);
  not g7063 (n_3913, n4548);
  and g7064 (n4549, n_3907, n_3913);
  not g7065 (n_3914, n4547);
  and g7066 (n4550, n_3914, n4549);
  not g7067 (n_3915, n4549);
  and g7068 (n4551, n4547, n_3915);
  not g7069 (n_3916, n4550);
  not g7070 (n_3917, n4551);
  and g7071 (n4552, n_3916, n_3917);
  not g7072 (n_3918, n4508);
  not g7073 (n_3919, n4552);
  and g7074 (n4553, n_3918, n_3919);
  and g7075 (n4554, n_3914, n_3915);
  not g7080 (n_3920, n4554);
  not g7081 (n_3921, n4558);
  and g7082 (n4559, n_3920, n_3921);
  not g7083 (n_3922, n4559);
  and g7084 (n4560, n4508, n_3922);
  not g7085 (n_3923, n4553);
  not g7086 (n_3924, n4560);
  and g7087 (n4561, n_3923, n_3924);
  and g7088 (n4562, \A[982] , \A[983] );
  not g7089 (n_3927, \A[983] );
  and g7090 (n4563, \A[982] , n_3927);
  not g7091 (n_3928, \A[982] );
  and g7092 (n4564, n_3928, \A[983] );
  not g7093 (n_3929, n4563);
  not g7094 (n_3930, n4564);
  and g7095 (n4565, n_3929, n_3930);
  not g7096 (n_3932, n4565);
  and g7097 (n4566, \A[984] , n_3932);
  not g7098 (n_3933, n4562);
  not g7099 (n_3934, n4566);
  and g7100 (n4567, n_3933, n_3934);
  and g7101 (n4568, \A[979] , \A[980] );
  not g7102 (n_3937, \A[980] );
  and g7103 (n4569, \A[979] , n_3937);
  not g7104 (n_3938, \A[979] );
  and g7105 (n4570, n_3938, \A[980] );
  not g7106 (n_3939, n4569);
  not g7107 (n_3940, n4570);
  and g7108 (n4571, n_3939, n_3940);
  not g7109 (n_3942, n4571);
  and g7110 (n4572, \A[981] , n_3942);
  not g7111 (n_3943, n4568);
  not g7112 (n_3944, n4572);
  and g7113 (n4573, n_3943, n_3944);
  not g7114 (n_3945, n4573);
  and g7115 (n4574, n4567, n_3945);
  not g7116 (n_3946, n4567);
  and g7117 (n4575, n_3946, n4573);
  and g7118 (n4576, \A[981] , n_3939);
  and g7119 (n4577, n_3940, n4576);
  not g7120 (n_3947, \A[981] );
  and g7121 (n4578, n_3947, n_3942);
  not g7122 (n_3948, n4577);
  not g7123 (n_3949, n4578);
  and g7124 (n4579, n_3948, n_3949);
  and g7125 (n4580, \A[984] , n_3929);
  and g7126 (n4581, n_3930, n4580);
  not g7127 (n_3950, \A[984] );
  and g7128 (n4582, n_3950, n_3932);
  not g7129 (n_3951, n4581);
  not g7130 (n_3952, n4582);
  and g7131 (n4583, n_3951, n_3952);
  not g7132 (n_3953, n4579);
  not g7133 (n_3954, n4583);
  and g7134 (n4584, n_3953, n_3954);
  not g7135 (n_3955, n4575);
  and g7136 (n4585, n_3955, n4584);
  not g7137 (n_3956, n4574);
  and g7138 (n4586, n_3956, n4585);
  and g7139 (n4587, n_3956, n_3955);
  not g7140 (n_3957, n4584);
  not g7141 (n_3958, n4587);
  and g7142 (n4588, n_3957, n_3958);
  not g7143 (n_3959, n4586);
  not g7144 (n_3960, n4588);
  and g7145 (n4589, n_3959, n_3960);
  and g7146 (n4590, n_3953, n4583);
  and g7147 (n4591, n4579, n_3954);
  not g7148 (n_3961, n4590);
  not g7149 (n_3962, n4591);
  and g7150 (n4592, n_3961, n_3962);
  and g7151 (n4593, n4584, n_3958);
  and g7152 (n4594, n_3946, n_3945);
  not g7153 (n_3963, n4593);
  not g7154 (n_3964, n4594);
  and g7155 (n4595, n_3963, n_3964);
  not g7156 (n_3965, n4592);
  not g7157 (n_3966, n4595);
  and g7158 (n4596, n_3965, n_3966);
  not g7159 (n_3967, n4589);
  not g7160 (n_3968, n4596);
  and g7161 (n4597, n_3967, n_3968);
  and g7162 (n4598, n_3967, n_3966);
  and g7163 (n4599, \A[988] , \A[989] );
  not g7164 (n_3971, \A[989] );
  and g7165 (n4600, \A[988] , n_3971);
  not g7166 (n_3972, \A[988] );
  and g7167 (n4601, n_3972, \A[989] );
  not g7168 (n_3973, n4600);
  not g7169 (n_3974, n4601);
  and g7170 (n4602, n_3973, n_3974);
  not g7171 (n_3976, n4602);
  and g7172 (n4603, \A[990] , n_3976);
  not g7173 (n_3977, n4599);
  not g7174 (n_3978, n4603);
  and g7175 (n4604, n_3977, n_3978);
  and g7176 (n4605, \A[985] , \A[986] );
  not g7177 (n_3981, \A[986] );
  and g7178 (n4606, \A[985] , n_3981);
  not g7179 (n_3982, \A[985] );
  and g7180 (n4607, n_3982, \A[986] );
  not g7181 (n_3983, n4606);
  not g7182 (n_3984, n4607);
  and g7183 (n4608, n_3983, n_3984);
  not g7184 (n_3986, n4608);
  and g7185 (n4609, \A[987] , n_3986);
  not g7186 (n_3987, n4605);
  not g7187 (n_3988, n4609);
  and g7188 (n4610, n_3987, n_3988);
  not g7189 (n_3989, n4604);
  and g7190 (n4611, n_3989, n4610);
  not g7191 (n_3990, n4610);
  and g7192 (n4612, n4604, n_3990);
  not g7193 (n_3991, n4611);
  not g7194 (n_3992, n4612);
  and g7195 (n4613, n_3991, n_3992);
  and g7196 (n4614, \A[987] , n_3983);
  and g7197 (n4615, n_3984, n4614);
  not g7198 (n_3993, \A[987] );
  and g7199 (n4616, n_3993, n_3986);
  not g7200 (n_3994, n4615);
  not g7201 (n_3995, n4616);
  and g7202 (n4617, n_3994, n_3995);
  and g7203 (n4618, \A[990] , n_3973);
  and g7204 (n4619, n_3974, n4618);
  not g7205 (n_3996, \A[990] );
  and g7206 (n4620, n_3996, n_3976);
  not g7207 (n_3997, n4619);
  not g7208 (n_3998, n4620);
  and g7209 (n4621, n_3997, n_3998);
  not g7210 (n_3999, n4617);
  not g7211 (n_4000, n4621);
  and g7212 (n4622, n_3999, n_4000);
  not g7213 (n_4001, n4613);
  and g7214 (n4623, n_4001, n4622);
  and g7215 (n4624, n_3989, n_3990);
  not g7216 (n_4002, n4623);
  not g7217 (n_4003, n4624);
  and g7218 (n4625, n_4002, n_4003);
  and g7219 (n4626, n_3991, n4622);
  and g7220 (n4627, n_3992, n4626);
  not g7221 (n_4004, n4622);
  and g7222 (n4628, n_4001, n_4004);
  not g7223 (n_4005, n4627);
  not g7224 (n_4006, n4628);
  and g7225 (n4629, n_4005, n_4006);
  not g7226 (n_4007, n4625);
  not g7227 (n_4008, n4629);
  and g7228 (n4630, n_4007, n_4008);
  and g7229 (n4631, n_3999, n4621);
  and g7230 (n4632, n4617, n_4000);
  not g7231 (n_4009, n4631);
  not g7232 (n_4010, n4632);
  and g7233 (n4633, n_4009, n_4010);
  not g7234 (n_4011, n4633);
  and g7235 (n4634, n_3965, n_4011);
  not g7236 (n_4012, n4630);
  and g7237 (n4635, n_4012, n4634);
  not g7238 (n_4013, n4598);
  and g7239 (n4636, n_4013, n4635);
  and g7240 (n4637, n_4007, n_4011);
  not g7241 (n_4014, n4637);
  and g7242 (n4638, n_4008, n_4014);
  not g7243 (n_4015, n4636);
  not g7244 (n_4016, n4638);
  and g7245 (n4639, n_4015, n_4016);
  not g7250 (n_4017, n4639);
  not g7251 (n_4018, n4643);
  and g7252 (n4644, n_4017, n_4018);
  not g7253 (n_4019, n4644);
  and g7254 (n4645, n4597, n_4019);
  and g7255 (n4646, n_4015, n4638);
  and g7256 (n4647, n4636, n_4016);
  not g7257 (n_4020, n4646);
  not g7258 (n_4021, n4647);
  and g7259 (n4648, n_4020, n_4021);
  not g7260 (n_4022, n4597);
  not g7261 (n_4023, n4648);
  and g7262 (n4649, n_4022, n_4023);
  and g7263 (n4650, n_4012, n_4011);
  and g7264 (n4651, n_3965, n_4013);
  not g7265 (n_4024, n4650);
  and g7266 (n4652, n_4024, n4651);
  not g7267 (n_4025, n4651);
  and g7268 (n4653, n4650, n_4025);
  not g7269 (n_4026, n4652);
  not g7270 (n_4027, n4653);
  and g7271 (n4654, n_4026, n_4027);
  and g7272 (n4655, n_3911, n_3910);
  and g7273 (n4656, n_3864, n_3912);
  not g7274 (n_4028, n4655);
  and g7275 (n4657, n_4028, n4656);
  not g7276 (n_4029, n4656);
  and g7277 (n4658, n4655, n_4029);
  not g7278 (n_4030, n4657);
  not g7279 (n_4031, n4658);
  and g7280 (n4659, n_4030, n_4031);
  not g7281 (n_4032, n4654);
  not g7282 (n_4033, n4659);
  and g7283 (n4660, n_4032, n_4033);
  not g7284 (n_4034, n4649);
  not g7285 (n_4035, n4660);
  and g7286 (n4661, n_4034, n_4035);
  not g7287 (n_4036, n4645);
  and g7288 (n4662, n_4036, n4661);
  and g7289 (n4663, n_4036, n_4034);
  not g7290 (n_4037, n4663);
  and g7291 (n4664, n4660, n_4037);
  not g7292 (n_4038, n4662);
  not g7293 (n_4039, n4664);
  and g7294 (n4665, n_4038, n_4039);
  not g7295 (n_4040, n4561);
  not g7296 (n_4041, n4665);
  and g7297 (n4666, n_4040, n_4041);
  and g7298 (n4667, n_4034, n4660);
  and g7299 (n4668, n_4036, n4667);
  and g7300 (n4669, n_4035, n_4037);
  not g7301 (n_4042, n4668);
  not g7302 (n_4043, n4669);
  and g7303 (n4670, n_4042, n_4043);
  not g7304 (n_4044, n4670);
  and g7305 (n4671, n4561, n_4044);
  and g7306 (n4672, n_4032, n4659);
  and g7307 (n4673, n4654, n_4033);
  not g7308 (n_4045, n4672);
  not g7309 (n_4046, n4673);
  and g7310 (n4674, n_4045, n_4046);
  not g7311 (n_4048, \A[961] );
  and g7312 (n4675, n_4048, \A[962] );
  not g7313 (n_4050, \A[962] );
  and g7314 (n4676, \A[961] , n_4050);
  not g7315 (n_4052, n4676);
  and g7316 (n4677, \A[963] , n_4052);
  not g7317 (n_4053, n4675);
  and g7318 (n4678, n_4053, n4677);
  and g7319 (n4679, n_4053, n_4052);
  not g7320 (n_4054, \A[963] );
  not g7321 (n_4055, n4679);
  and g7322 (n4680, n_4054, n_4055);
  not g7323 (n_4056, n4678);
  not g7324 (n_4057, n4680);
  and g7325 (n4681, n_4056, n_4057);
  not g7326 (n_4059, \A[964] );
  and g7327 (n4682, n_4059, \A[965] );
  not g7328 (n_4061, \A[965] );
  and g7329 (n4683, \A[964] , n_4061);
  not g7330 (n_4063, n4683);
  and g7331 (n4684, \A[966] , n_4063);
  not g7332 (n_4064, n4682);
  and g7333 (n4685, n_4064, n4684);
  and g7334 (n4686, n_4064, n_4063);
  not g7335 (n_4065, \A[966] );
  not g7336 (n_4066, n4686);
  and g7337 (n4687, n_4065, n_4066);
  not g7338 (n_4067, n4685);
  not g7339 (n_4068, n4687);
  and g7340 (n4688, n_4067, n_4068);
  not g7341 (n_4069, n4681);
  and g7342 (n4689, n_4069, n4688);
  not g7343 (n_4070, n4688);
  and g7344 (n4690, n4681, n_4070);
  not g7345 (n_4071, n4689);
  not g7346 (n_4072, n4690);
  and g7347 (n4691, n_4071, n_4072);
  and g7348 (n4692, \A[964] , \A[965] );
  and g7349 (n4693, \A[966] , n_4066);
  not g7350 (n_4073, n4692);
  not g7351 (n_4074, n4693);
  and g7352 (n4694, n_4073, n_4074);
  and g7353 (n4695, \A[961] , \A[962] );
  and g7354 (n4696, \A[963] , n_4055);
  not g7355 (n_4075, n4695);
  not g7356 (n_4076, n4696);
  and g7357 (n4697, n_4075, n_4076);
  not g7358 (n_4077, n4694);
  and g7359 (n4698, n_4077, n4697);
  not g7360 (n_4078, n4697);
  and g7361 (n4699, n4694, n_4078);
  not g7362 (n_4079, n4698);
  not g7363 (n_4080, n4699);
  and g7364 (n4700, n_4079, n_4080);
  and g7365 (n4701, n_4069, n_4070);
  not g7366 (n_4081, n4700);
  and g7367 (n4702, n_4081, n4701);
  and g7368 (n4703, n_4077, n_4078);
  not g7369 (n_4082, n4702);
  not g7370 (n_4083, n4703);
  and g7371 (n4704, n_4082, n_4083);
  and g7372 (n4705, n_4079, n4701);
  and g7373 (n4706, n_4080, n4705);
  not g7374 (n_4084, n4701);
  and g7375 (n4707, n_4081, n_4084);
  not g7376 (n_4085, n4706);
  not g7377 (n_4086, n4707);
  and g7378 (n4708, n_4085, n_4086);
  not g7379 (n_4087, n4704);
  not g7380 (n_4088, n4708);
  and g7381 (n4709, n_4087, n_4088);
  not g7382 (n_4089, n4691);
  not g7383 (n_4090, n4709);
  and g7384 (n4710, n_4089, n_4090);
  not g7385 (n_4092, \A[955] );
  and g7386 (n4711, n_4092, \A[956] );
  not g7387 (n_4094, \A[956] );
  and g7388 (n4712, \A[955] , n_4094);
  not g7389 (n_4096, n4712);
  and g7390 (n4713, \A[957] , n_4096);
  not g7391 (n_4097, n4711);
  and g7392 (n4714, n_4097, n4713);
  and g7393 (n4715, n_4097, n_4096);
  not g7394 (n_4098, \A[957] );
  not g7395 (n_4099, n4715);
  and g7396 (n4716, n_4098, n_4099);
  not g7397 (n_4100, n4714);
  not g7398 (n_4101, n4716);
  and g7399 (n4717, n_4100, n_4101);
  not g7400 (n_4103, \A[958] );
  and g7401 (n4718, n_4103, \A[959] );
  not g7402 (n_4105, \A[959] );
  and g7403 (n4719, \A[958] , n_4105);
  not g7404 (n_4107, n4719);
  and g7405 (n4720, \A[960] , n_4107);
  not g7406 (n_4108, n4718);
  and g7407 (n4721, n_4108, n4720);
  and g7408 (n4722, n_4108, n_4107);
  not g7409 (n_4109, \A[960] );
  not g7410 (n_4110, n4722);
  and g7411 (n4723, n_4109, n_4110);
  not g7412 (n_4111, n4721);
  not g7413 (n_4112, n4723);
  and g7414 (n4724, n_4111, n_4112);
  not g7415 (n_4113, n4717);
  and g7416 (n4725, n_4113, n4724);
  not g7417 (n_4114, n4724);
  and g7418 (n4726, n4717, n_4114);
  not g7419 (n_4115, n4725);
  not g7420 (n_4116, n4726);
  and g7421 (n4727, n_4115, n_4116);
  and g7422 (n4728, \A[958] , \A[959] );
  and g7423 (n4729, \A[960] , n_4110);
  not g7424 (n_4117, n4728);
  not g7425 (n_4118, n4729);
  and g7426 (n4730, n_4117, n_4118);
  and g7427 (n4731, \A[955] , \A[956] );
  and g7428 (n4732, \A[957] , n_4099);
  not g7429 (n_4119, n4731);
  not g7430 (n_4120, n4732);
  and g7431 (n4733, n_4119, n_4120);
  not g7432 (n_4121, n4730);
  and g7433 (n4734, n_4121, n4733);
  not g7434 (n_4122, n4733);
  and g7435 (n4735, n4730, n_4122);
  not g7436 (n_4123, n4734);
  not g7437 (n_4124, n4735);
  and g7438 (n4736, n_4123, n_4124);
  and g7439 (n4737, n_4113, n_4114);
  not g7440 (n_4125, n4736);
  and g7441 (n4738, n_4125, n4737);
  and g7442 (n4739, n_4121, n_4122);
  not g7443 (n_4126, n4738);
  not g7444 (n_4127, n4739);
  and g7445 (n4740, n_4126, n_4127);
  and g7446 (n4741, n_4123, n4737);
  and g7447 (n4742, n_4124, n4741);
  not g7448 (n_4128, n4737);
  and g7449 (n4743, n_4125, n_4128);
  not g7450 (n_4129, n4742);
  not g7451 (n_4130, n4743);
  and g7452 (n4744, n_4129, n_4130);
  not g7453 (n_4131, n4740);
  not g7454 (n_4132, n4744);
  and g7455 (n4745, n_4131, n_4132);
  not g7456 (n_4133, n4727);
  not g7457 (n_4134, n4745);
  and g7458 (n4746, n_4133, n_4134);
  not g7459 (n_4135, n4710);
  and g7460 (n4747, n_4135, n4746);
  not g7461 (n_4136, n4746);
  and g7462 (n4748, n4710, n_4136);
  not g7463 (n_4137, n4747);
  not g7464 (n_4138, n4748);
  and g7465 (n4749, n_4137, n_4138);
  not g7466 (n_4140, \A[949] );
  and g7467 (n4750, n_4140, \A[950] );
  not g7468 (n_4142, \A[950] );
  and g7469 (n4751, \A[949] , n_4142);
  not g7470 (n_4144, n4751);
  and g7471 (n4752, \A[951] , n_4144);
  not g7472 (n_4145, n4750);
  and g7473 (n4753, n_4145, n4752);
  and g7474 (n4754, n_4145, n_4144);
  not g7475 (n_4146, \A[951] );
  not g7476 (n_4147, n4754);
  and g7477 (n4755, n_4146, n_4147);
  not g7478 (n_4148, n4753);
  not g7479 (n_4149, n4755);
  and g7480 (n4756, n_4148, n_4149);
  not g7481 (n_4151, \A[952] );
  and g7482 (n4757, n_4151, \A[953] );
  not g7483 (n_4153, \A[953] );
  and g7484 (n4758, \A[952] , n_4153);
  not g7485 (n_4155, n4758);
  and g7486 (n4759, \A[954] , n_4155);
  not g7487 (n_4156, n4757);
  and g7488 (n4760, n_4156, n4759);
  and g7489 (n4761, n_4156, n_4155);
  not g7490 (n_4157, \A[954] );
  not g7491 (n_4158, n4761);
  and g7492 (n4762, n_4157, n_4158);
  not g7493 (n_4159, n4760);
  not g7494 (n_4160, n4762);
  and g7495 (n4763, n_4159, n_4160);
  not g7496 (n_4161, n4756);
  and g7497 (n4764, n_4161, n4763);
  not g7498 (n_4162, n4763);
  and g7499 (n4765, n4756, n_4162);
  not g7500 (n_4163, n4764);
  not g7501 (n_4164, n4765);
  and g7502 (n4766, n_4163, n_4164);
  and g7503 (n4767, \A[952] , \A[953] );
  and g7504 (n4768, \A[954] , n_4158);
  not g7505 (n_4165, n4767);
  not g7506 (n_4166, n4768);
  and g7507 (n4769, n_4165, n_4166);
  and g7508 (n4770, \A[949] , \A[950] );
  and g7509 (n4771, \A[951] , n_4147);
  not g7510 (n_4167, n4770);
  not g7511 (n_4168, n4771);
  and g7512 (n4772, n_4167, n_4168);
  not g7513 (n_4169, n4769);
  and g7514 (n4773, n_4169, n4772);
  not g7515 (n_4170, n4772);
  and g7516 (n4774, n4769, n_4170);
  not g7517 (n_4171, n4773);
  not g7518 (n_4172, n4774);
  and g7519 (n4775, n_4171, n_4172);
  and g7520 (n4776, n_4161, n_4162);
  not g7521 (n_4173, n4775);
  and g7522 (n4777, n_4173, n4776);
  and g7523 (n4778, n_4169, n_4170);
  not g7524 (n_4174, n4777);
  not g7525 (n_4175, n4778);
  and g7526 (n4779, n_4174, n_4175);
  and g7527 (n4780, n_4171, n4776);
  and g7528 (n4781, n_4172, n4780);
  not g7529 (n_4176, n4776);
  and g7530 (n4782, n_4173, n_4176);
  not g7531 (n_4177, n4781);
  not g7532 (n_4178, n4782);
  and g7533 (n4783, n_4177, n_4178);
  not g7534 (n_4179, n4779);
  not g7535 (n_4180, n4783);
  and g7536 (n4784, n_4179, n_4180);
  not g7537 (n_4181, n4766);
  not g7538 (n_4182, n4784);
  and g7539 (n4785, n_4181, n_4182);
  not g7540 (n_4184, \A[943] );
  and g7541 (n4786, n_4184, \A[944] );
  not g7542 (n_4186, \A[944] );
  and g7543 (n4787, \A[943] , n_4186);
  not g7544 (n_4188, n4787);
  and g7545 (n4788, \A[945] , n_4188);
  not g7546 (n_4189, n4786);
  and g7547 (n4789, n_4189, n4788);
  and g7548 (n4790, n_4189, n_4188);
  not g7549 (n_4190, \A[945] );
  not g7550 (n_4191, n4790);
  and g7551 (n4791, n_4190, n_4191);
  not g7552 (n_4192, n4789);
  not g7553 (n_4193, n4791);
  and g7554 (n4792, n_4192, n_4193);
  not g7555 (n_4195, \A[946] );
  and g7556 (n4793, n_4195, \A[947] );
  not g7557 (n_4197, \A[947] );
  and g7558 (n4794, \A[946] , n_4197);
  not g7559 (n_4199, n4794);
  and g7560 (n4795, \A[948] , n_4199);
  not g7561 (n_4200, n4793);
  and g7562 (n4796, n_4200, n4795);
  and g7563 (n4797, n_4200, n_4199);
  not g7564 (n_4201, \A[948] );
  not g7565 (n_4202, n4797);
  and g7566 (n4798, n_4201, n_4202);
  not g7567 (n_4203, n4796);
  not g7568 (n_4204, n4798);
  and g7569 (n4799, n_4203, n_4204);
  not g7570 (n_4205, n4792);
  and g7571 (n4800, n_4205, n4799);
  not g7572 (n_4206, n4799);
  and g7573 (n4801, n4792, n_4206);
  not g7574 (n_4207, n4800);
  not g7575 (n_4208, n4801);
  and g7576 (n4802, n_4207, n_4208);
  and g7577 (n4803, \A[946] , \A[947] );
  and g7578 (n4804, \A[948] , n_4202);
  not g7579 (n_4209, n4803);
  not g7580 (n_4210, n4804);
  and g7581 (n4805, n_4209, n_4210);
  and g7582 (n4806, \A[943] , \A[944] );
  and g7583 (n4807, \A[945] , n_4191);
  not g7584 (n_4211, n4806);
  not g7585 (n_4212, n4807);
  and g7586 (n4808, n_4211, n_4212);
  not g7587 (n_4213, n4805);
  and g7588 (n4809, n_4213, n4808);
  not g7589 (n_4214, n4808);
  and g7590 (n4810, n4805, n_4214);
  not g7591 (n_4215, n4809);
  not g7592 (n_4216, n4810);
  and g7593 (n4811, n_4215, n_4216);
  and g7594 (n4812, n_4205, n_4206);
  not g7595 (n_4217, n4811);
  and g7596 (n4813, n_4217, n4812);
  and g7597 (n4814, n_4213, n_4214);
  not g7598 (n_4218, n4813);
  not g7599 (n_4219, n4814);
  and g7600 (n4815, n_4218, n_4219);
  and g7601 (n4816, n_4215, n4812);
  and g7602 (n4817, n_4216, n4816);
  not g7603 (n_4220, n4812);
  and g7604 (n4818, n_4217, n_4220);
  not g7605 (n_4221, n4817);
  not g7606 (n_4222, n4818);
  and g7607 (n4819, n_4221, n_4222);
  not g7608 (n_4223, n4815);
  not g7609 (n_4224, n4819);
  and g7610 (n4820, n_4223, n_4224);
  not g7611 (n_4225, n4802);
  not g7612 (n_4226, n4820);
  and g7613 (n4821, n_4225, n_4226);
  not g7614 (n_4227, n4785);
  and g7615 (n4822, n_4227, n4821);
  not g7616 (n_4228, n4821);
  and g7617 (n4823, n4785, n_4228);
  not g7618 (n_4229, n4822);
  not g7619 (n_4230, n4823);
  and g7620 (n4824, n_4229, n_4230);
  not g7621 (n_4231, n4749);
  and g7622 (n4825, n_4231, n4824);
  not g7623 (n_4232, n4824);
  and g7624 (n4826, n4749, n_4232);
  not g7625 (n_4233, n4825);
  not g7626 (n_4234, n4826);
  and g7627 (n4827, n_4233, n_4234);
  not g7628 (n_4235, n4674);
  not g7629 (n_4236, n4827);
  and g7630 (n4828, n_4235, n_4236);
  not g7631 (n_4237, n4671);
  and g7632 (n4829, n_4237, n4828);
  not g7633 (n_4238, n4666);
  and g7634 (n4830, n_4238, n4829);
  and g7635 (n4831, n_4238, n_4237);
  not g7636 (n_4239, n4828);
  not g7637 (n_4240, n4831);
  and g7638 (n4832, n_4239, n_4240);
  not g7639 (n_4241, n4830);
  not g7640 (n_4242, n4832);
  and g7641 (n4833, n_4241, n_4242);
  and g7642 (n4834, n_4133, n_4131);
  not g7643 (n_4243, n4834);
  and g7644 (n4835, n_4132, n_4243);
  and g7645 (n4836, n_4089, n_4133);
  and g7646 (n4837, n_4090, n4836);
  and g7647 (n4838, n_4134, n4837);
  and g7648 (n4839, n_4089, n_4087);
  not g7649 (n_4244, n4839);
  and g7650 (n4840, n_4088, n_4244);
  not g7651 (n_4245, n4838);
  not g7652 (n_4246, n4840);
  and g7653 (n4841, n_4245, n_4246);
  not g7658 (n_4247, n4841);
  not g7659 (n_4248, n4845);
  and g7660 (n4846, n_4247, n_4248);
  not g7661 (n_4249, n4846);
  and g7662 (n4847, n4835, n_4249);
  and g7663 (n4848, n_4245, n4840);
  and g7664 (n4849, n4838, n_4246);
  not g7665 (n_4250, n4848);
  not g7666 (n_4251, n4849);
  and g7667 (n4850, n_4250, n_4251);
  not g7668 (n_4252, n4835);
  not g7669 (n_4253, n4850);
  and g7670 (n4851, n_4252, n_4253);
  and g7671 (n4852, n_4231, n_4232);
  not g7672 (n_4254, n4851);
  and g7673 (n4853, n_4254, n4852);
  not g7674 (n_4255, n4847);
  and g7675 (n4854, n_4255, n4853);
  and g7676 (n4855, n_4255, n_4254);
  not g7677 (n_4256, n4852);
  not g7678 (n_4257, n4855);
  and g7679 (n4856, n_4256, n_4257);
  not g7680 (n_4258, n4854);
  not g7681 (n_4259, n4856);
  and g7682 (n4857, n_4258, n_4259);
  and g7683 (n4858, n_4225, n_4223);
  not g7684 (n_4260, n4858);
  and g7685 (n4859, n_4224, n_4260);
  and g7686 (n4860, n_4181, n_4225);
  and g7687 (n4861, n_4182, n4860);
  and g7688 (n4862, n_4226, n4861);
  and g7689 (n4863, n_4181, n_4179);
  not g7690 (n_4261, n4863);
  and g7691 (n4864, n_4180, n_4261);
  not g7692 (n_4262, n4862);
  and g7693 (n4865, n_4262, n4864);
  not g7694 (n_4263, n4864);
  and g7695 (n4866, n4862, n_4263);
  not g7696 (n_4264, n4865);
  not g7697 (n_4265, n4866);
  and g7698 (n4867, n_4264, n_4265);
  not g7699 (n_4266, n4859);
  not g7700 (n_4267, n4867);
  and g7701 (n4868, n_4266, n_4267);
  and g7702 (n4869, n_4262, n_4263);
  not g7707 (n_4268, n4869);
  not g7708 (n_4269, n4873);
  and g7709 (n4874, n_4268, n_4269);
  not g7710 (n_4270, n4874);
  and g7711 (n4875, n4859, n_4270);
  not g7712 (n_4271, n4868);
  not g7713 (n_4272, n4875);
  and g7714 (n4876, n_4271, n_4272);
  not g7715 (n_4273, n4857);
  and g7716 (n4877, n_4273, n4876);
  and g7717 (n4878, n_4254, n_4256);
  and g7718 (n4879, n_4255, n4878);
  and g7719 (n4880, n4852, n_4257);
  not g7720 (n_4274, n4879);
  not g7721 (n_4275, n4880);
  and g7722 (n4881, n_4274, n_4275);
  not g7723 (n_4276, n4876);
  not g7724 (n_4277, n4881);
  and g7725 (n4882, n_4276, n_4277);
  not g7726 (n_4278, n4877);
  not g7727 (n_4279, n4882);
  and g7728 (n4883, n_4278, n_4279);
  not g7729 (n_4280, n4833);
  and g7730 (n4884, n_4280, n4883);
  and g7731 (n4885, n_4237, n_4239);
  and g7732 (n4886, n_4238, n4885);
  and g7733 (n4887, n4828, n_4240);
  not g7734 (n_4281, n4886);
  not g7735 (n_4282, n4887);
  and g7736 (n4888, n_4281, n_4282);
  not g7737 (n_4283, n4883);
  not g7738 (n_4284, n4888);
  and g7739 (n4889, n_4283, n_4284);
  not g7740 (n_4285, n4884);
  not g7741 (n_4286, n4889);
  and g7742 (n4890, n_4285, n_4286);
  and g7743 (n4891, \A[10] , \A[11] );
  not g7744 (n_4289, \A[11] );
  and g7745 (n4892, \A[10] , n_4289);
  not g7746 (n_4290, \A[10] );
  and g7747 (n4893, n_4290, \A[11] );
  not g7748 (n_4291, n4892);
  not g7749 (n_4292, n4893);
  and g7750 (n4894, n_4291, n_4292);
  not g7751 (n_4294, n4894);
  and g7752 (n4895, \A[12] , n_4294);
  not g7753 (n_4295, n4891);
  not g7754 (n_4296, n4895);
  and g7755 (n4896, n_4295, n_4296);
  and g7756 (n4897, \A[7] , \A[8] );
  not g7757 (n_4299, \A[8] );
  and g7758 (n4898, \A[7] , n_4299);
  not g7759 (n_4300, \A[7] );
  and g7760 (n4899, n_4300, \A[8] );
  not g7761 (n_4301, n4898);
  not g7762 (n_4302, n4899);
  and g7763 (n4900, n_4301, n_4302);
  not g7764 (n_4304, n4900);
  and g7765 (n4901, \A[9] , n_4304);
  not g7766 (n_4305, n4897);
  not g7767 (n_4306, n4901);
  and g7768 (n4902, n_4305, n_4306);
  not g7769 (n_4307, n4902);
  and g7770 (n4903, n4896, n_4307);
  not g7771 (n_4308, n4896);
  and g7772 (n4904, n_4308, n4902);
  and g7773 (n4905, \A[9] , n_4301);
  and g7774 (n4906, n_4302, n4905);
  not g7775 (n_4309, \A[9] );
  and g7776 (n4907, n_4309, n_4304);
  not g7777 (n_4310, n4906);
  not g7778 (n_4311, n4907);
  and g7779 (n4908, n_4310, n_4311);
  and g7780 (n4909, \A[12] , n_4291);
  and g7781 (n4910, n_4292, n4909);
  not g7782 (n_4312, \A[12] );
  and g7783 (n4911, n_4312, n_4294);
  not g7784 (n_4313, n4910);
  not g7785 (n_4314, n4911);
  and g7786 (n4912, n_4313, n_4314);
  not g7787 (n_4315, n4908);
  not g7788 (n_4316, n4912);
  and g7789 (n4913, n_4315, n_4316);
  not g7790 (n_4317, n4904);
  and g7791 (n4914, n_4317, n4913);
  not g7792 (n_4318, n4903);
  and g7793 (n4915, n_4318, n4914);
  and g7794 (n4916, n_4318, n_4317);
  not g7795 (n_4319, n4913);
  not g7796 (n_4320, n4916);
  and g7797 (n4917, n_4319, n_4320);
  not g7798 (n_4321, n4915);
  not g7799 (n_4322, n4917);
  and g7800 (n4918, n_4321, n_4322);
  and g7801 (n4919, n_4315, n4912);
  and g7802 (n4920, n4908, n_4316);
  not g7803 (n_4323, n4919);
  not g7804 (n_4324, n4920);
  and g7805 (n4921, n_4323, n_4324);
  and g7806 (n4922, n4913, n_4320);
  and g7807 (n4923, n_4308, n_4307);
  not g7808 (n_4325, n4922);
  not g7809 (n_4326, n4923);
  and g7810 (n4924, n_4325, n_4326);
  not g7811 (n_4327, n4921);
  not g7812 (n_4328, n4924);
  and g7813 (n4925, n_4327, n_4328);
  not g7814 (n_4329, n4918);
  not g7815 (n_4330, n4925);
  and g7816 (n4926, n_4329, n_4330);
  and g7817 (n4927, n_4329, n_4328);
  and g7818 (n4928, \A[16] , \A[17] );
  not g7819 (n_4333, \A[17] );
  and g7820 (n4929, \A[16] , n_4333);
  not g7821 (n_4334, \A[16] );
  and g7822 (n4930, n_4334, \A[17] );
  not g7823 (n_4335, n4929);
  not g7824 (n_4336, n4930);
  and g7825 (n4931, n_4335, n_4336);
  not g7826 (n_4338, n4931);
  and g7827 (n4932, \A[18] , n_4338);
  not g7828 (n_4339, n4928);
  not g7829 (n_4340, n4932);
  and g7830 (n4933, n_4339, n_4340);
  and g7831 (n4934, \A[13] , \A[14] );
  not g7832 (n_4343, \A[14] );
  and g7833 (n4935, \A[13] , n_4343);
  not g7834 (n_4344, \A[13] );
  and g7835 (n4936, n_4344, \A[14] );
  not g7836 (n_4345, n4935);
  not g7837 (n_4346, n4936);
  and g7838 (n4937, n_4345, n_4346);
  not g7839 (n_4348, n4937);
  and g7840 (n4938, \A[15] , n_4348);
  not g7841 (n_4349, n4934);
  not g7842 (n_4350, n4938);
  and g7843 (n4939, n_4349, n_4350);
  not g7844 (n_4351, n4933);
  and g7845 (n4940, n_4351, n4939);
  not g7846 (n_4352, n4939);
  and g7847 (n4941, n4933, n_4352);
  not g7848 (n_4353, n4940);
  not g7849 (n_4354, n4941);
  and g7850 (n4942, n_4353, n_4354);
  and g7851 (n4943, \A[15] , n_4345);
  and g7852 (n4944, n_4346, n4943);
  not g7853 (n_4355, \A[15] );
  and g7854 (n4945, n_4355, n_4348);
  not g7855 (n_4356, n4944);
  not g7856 (n_4357, n4945);
  and g7857 (n4946, n_4356, n_4357);
  and g7858 (n4947, \A[18] , n_4335);
  and g7859 (n4948, n_4336, n4947);
  not g7860 (n_4358, \A[18] );
  and g7861 (n4949, n_4358, n_4338);
  not g7862 (n_4359, n4948);
  not g7863 (n_4360, n4949);
  and g7864 (n4950, n_4359, n_4360);
  not g7865 (n_4361, n4946);
  not g7866 (n_4362, n4950);
  and g7867 (n4951, n_4361, n_4362);
  not g7868 (n_4363, n4942);
  and g7869 (n4952, n_4363, n4951);
  and g7870 (n4953, n_4351, n_4352);
  not g7871 (n_4364, n4952);
  not g7872 (n_4365, n4953);
  and g7873 (n4954, n_4364, n_4365);
  and g7874 (n4955, n_4353, n4951);
  and g7875 (n4956, n_4354, n4955);
  not g7876 (n_4366, n4951);
  and g7877 (n4957, n_4363, n_4366);
  not g7878 (n_4367, n4956);
  not g7879 (n_4368, n4957);
  and g7880 (n4958, n_4367, n_4368);
  not g7881 (n_4369, n4954);
  not g7882 (n_4370, n4958);
  and g7883 (n4959, n_4369, n_4370);
  and g7884 (n4960, n_4361, n4950);
  and g7885 (n4961, n4946, n_4362);
  not g7886 (n_4371, n4960);
  not g7887 (n_4372, n4961);
  and g7888 (n4962, n_4371, n_4372);
  not g7889 (n_4373, n4962);
  and g7890 (n4963, n_4327, n_4373);
  not g7891 (n_4374, n4959);
  and g7892 (n4964, n_4374, n4963);
  not g7893 (n_4375, n4927);
  and g7894 (n4965, n_4375, n4964);
  and g7895 (n4966, n_4369, n_4373);
  not g7896 (n_4376, n4966);
  and g7897 (n4967, n_4370, n_4376);
  not g7898 (n_4377, n4965);
  and g7899 (n4968, n_4377, n4967);
  not g7900 (n_4378, n4967);
  and g7901 (n4969, n4965, n_4378);
  not g7902 (n_4379, n4968);
  not g7903 (n_4380, n4969);
  and g7904 (n4970, n_4379, n_4380);
  not g7905 (n_4381, n4926);
  not g7906 (n_4382, n4970);
  and g7907 (n4971, n_4381, n_4382);
  and g7908 (n4972, n_4377, n_4378);
  not g7913 (n_4383, n4972);
  not g7914 (n_4384, n4976);
  and g7915 (n4977, n_4383, n_4384);
  not g7916 (n_4385, n4977);
  and g7917 (n4978, n4926, n_4385);
  not g7918 (n_4386, n4971);
  not g7919 (n_4387, n4978);
  and g7920 (n4979, n_4386, n_4387);
  and g7921 (n4980, \A[22] , \A[23] );
  not g7922 (n_4390, \A[23] );
  and g7923 (n4981, \A[22] , n_4390);
  not g7924 (n_4391, \A[22] );
  and g7925 (n4982, n_4391, \A[23] );
  not g7926 (n_4392, n4981);
  not g7927 (n_4393, n4982);
  and g7928 (n4983, n_4392, n_4393);
  not g7929 (n_4395, n4983);
  and g7930 (n4984, \A[24] , n_4395);
  not g7931 (n_4396, n4980);
  not g7932 (n_4397, n4984);
  and g7933 (n4985, n_4396, n_4397);
  and g7934 (n4986, \A[19] , \A[20] );
  not g7935 (n_4400, \A[20] );
  and g7936 (n4987, \A[19] , n_4400);
  not g7937 (n_4401, \A[19] );
  and g7938 (n4988, n_4401, \A[20] );
  not g7939 (n_4402, n4987);
  not g7940 (n_4403, n4988);
  and g7941 (n4989, n_4402, n_4403);
  not g7942 (n_4405, n4989);
  and g7943 (n4990, \A[21] , n_4405);
  not g7944 (n_4406, n4986);
  not g7945 (n_4407, n4990);
  and g7946 (n4991, n_4406, n_4407);
  not g7947 (n_4408, n4991);
  and g7948 (n4992, n4985, n_4408);
  not g7949 (n_4409, n4985);
  and g7950 (n4993, n_4409, n4991);
  and g7951 (n4994, \A[21] , n_4402);
  and g7952 (n4995, n_4403, n4994);
  not g7953 (n_4410, \A[21] );
  and g7954 (n4996, n_4410, n_4405);
  not g7955 (n_4411, n4995);
  not g7956 (n_4412, n4996);
  and g7957 (n4997, n_4411, n_4412);
  and g7958 (n4998, \A[24] , n_4392);
  and g7959 (n4999, n_4393, n4998);
  not g7960 (n_4413, \A[24] );
  and g7961 (n5000, n_4413, n_4395);
  not g7962 (n_4414, n4999);
  not g7963 (n_4415, n5000);
  and g7964 (n5001, n_4414, n_4415);
  not g7965 (n_4416, n4997);
  not g7966 (n_4417, n5001);
  and g7967 (n5002, n_4416, n_4417);
  not g7968 (n_4418, n4993);
  and g7969 (n5003, n_4418, n5002);
  not g7970 (n_4419, n4992);
  and g7971 (n5004, n_4419, n5003);
  and g7972 (n5005, n_4419, n_4418);
  not g7973 (n_4420, n5002);
  not g7974 (n_4421, n5005);
  and g7975 (n5006, n_4420, n_4421);
  not g7976 (n_4422, n5004);
  not g7977 (n_4423, n5006);
  and g7978 (n5007, n_4422, n_4423);
  and g7979 (n5008, n_4416, n5001);
  and g7980 (n5009, n4997, n_4417);
  not g7981 (n_4424, n5008);
  not g7982 (n_4425, n5009);
  and g7983 (n5010, n_4424, n_4425);
  and g7984 (n5011, n5002, n_4421);
  and g7985 (n5012, n_4409, n_4408);
  not g7986 (n_4426, n5011);
  not g7987 (n_4427, n5012);
  and g7988 (n5013, n_4426, n_4427);
  not g7989 (n_4428, n5010);
  not g7990 (n_4429, n5013);
  and g7991 (n5014, n_4428, n_4429);
  not g7992 (n_4430, n5007);
  not g7993 (n_4431, n5014);
  and g7994 (n5015, n_4430, n_4431);
  and g7995 (n5016, n_4430, n_4429);
  and g7996 (n5017, \A[28] , \A[29] );
  not g7997 (n_4434, \A[29] );
  and g7998 (n5018, \A[28] , n_4434);
  not g7999 (n_4435, \A[28] );
  and g8000 (n5019, n_4435, \A[29] );
  not g8001 (n_4436, n5018);
  not g8002 (n_4437, n5019);
  and g8003 (n5020, n_4436, n_4437);
  not g8004 (n_4439, n5020);
  and g8005 (n5021, \A[30] , n_4439);
  not g8006 (n_4440, n5017);
  not g8007 (n_4441, n5021);
  and g8008 (n5022, n_4440, n_4441);
  and g8009 (n5023, \A[25] , \A[26] );
  not g8010 (n_4444, \A[26] );
  and g8011 (n5024, \A[25] , n_4444);
  not g8012 (n_4445, \A[25] );
  and g8013 (n5025, n_4445, \A[26] );
  not g8014 (n_4446, n5024);
  not g8015 (n_4447, n5025);
  and g8016 (n5026, n_4446, n_4447);
  not g8017 (n_4449, n5026);
  and g8018 (n5027, \A[27] , n_4449);
  not g8019 (n_4450, n5023);
  not g8020 (n_4451, n5027);
  and g8021 (n5028, n_4450, n_4451);
  not g8022 (n_4452, n5022);
  and g8023 (n5029, n_4452, n5028);
  not g8024 (n_4453, n5028);
  and g8025 (n5030, n5022, n_4453);
  not g8026 (n_4454, n5029);
  not g8027 (n_4455, n5030);
  and g8028 (n5031, n_4454, n_4455);
  and g8029 (n5032, \A[27] , n_4446);
  and g8030 (n5033, n_4447, n5032);
  not g8031 (n_4456, \A[27] );
  and g8032 (n5034, n_4456, n_4449);
  not g8033 (n_4457, n5033);
  not g8034 (n_4458, n5034);
  and g8035 (n5035, n_4457, n_4458);
  and g8036 (n5036, \A[30] , n_4436);
  and g8037 (n5037, n_4437, n5036);
  not g8038 (n_4459, \A[30] );
  and g8039 (n5038, n_4459, n_4439);
  not g8040 (n_4460, n5037);
  not g8041 (n_4461, n5038);
  and g8042 (n5039, n_4460, n_4461);
  not g8043 (n_4462, n5035);
  not g8044 (n_4463, n5039);
  and g8045 (n5040, n_4462, n_4463);
  not g8046 (n_4464, n5031);
  and g8047 (n5041, n_4464, n5040);
  and g8048 (n5042, n_4452, n_4453);
  not g8049 (n_4465, n5041);
  not g8050 (n_4466, n5042);
  and g8051 (n5043, n_4465, n_4466);
  and g8052 (n5044, n_4454, n5040);
  and g8053 (n5045, n_4455, n5044);
  not g8054 (n_4467, n5040);
  and g8055 (n5046, n_4464, n_4467);
  not g8056 (n_4468, n5045);
  not g8057 (n_4469, n5046);
  and g8058 (n5047, n_4468, n_4469);
  not g8059 (n_4470, n5043);
  not g8060 (n_4471, n5047);
  and g8061 (n5048, n_4470, n_4471);
  and g8062 (n5049, n_4462, n5039);
  and g8063 (n5050, n5035, n_4463);
  not g8064 (n_4472, n5049);
  not g8065 (n_4473, n5050);
  and g8066 (n5051, n_4472, n_4473);
  not g8067 (n_4474, n5051);
  and g8068 (n5052, n_4428, n_4474);
  not g8069 (n_4475, n5048);
  and g8070 (n5053, n_4475, n5052);
  not g8071 (n_4476, n5016);
  and g8072 (n5054, n_4476, n5053);
  and g8073 (n5055, n_4470, n_4474);
  not g8074 (n_4477, n5055);
  and g8075 (n5056, n_4471, n_4477);
  not g8076 (n_4478, n5054);
  not g8077 (n_4479, n5056);
  and g8078 (n5057, n_4478, n_4479);
  not g8083 (n_4480, n5057);
  not g8084 (n_4481, n5061);
  and g8085 (n5062, n_4480, n_4481);
  not g8086 (n_4482, n5062);
  and g8087 (n5063, n5015, n_4482);
  and g8088 (n5064, n_4478, n5056);
  and g8089 (n5065, n5054, n_4479);
  not g8090 (n_4483, n5064);
  not g8091 (n_4484, n5065);
  and g8092 (n5066, n_4483, n_4484);
  not g8093 (n_4485, n5015);
  not g8094 (n_4486, n5066);
  and g8095 (n5067, n_4485, n_4486);
  and g8096 (n5068, n_4475, n_4474);
  and g8097 (n5069, n_4428, n_4476);
  not g8098 (n_4487, n5068);
  and g8099 (n5070, n_4487, n5069);
  not g8100 (n_4488, n5069);
  and g8101 (n5071, n5068, n_4488);
  not g8102 (n_4489, n5070);
  not g8103 (n_4490, n5071);
  and g8104 (n5072, n_4489, n_4490);
  and g8105 (n5073, n_4374, n_4373);
  and g8106 (n5074, n_4327, n_4375);
  not g8107 (n_4491, n5073);
  and g8108 (n5075, n_4491, n5074);
  not g8109 (n_4492, n5074);
  and g8110 (n5076, n5073, n_4492);
  not g8111 (n_4493, n5075);
  not g8112 (n_4494, n5076);
  and g8113 (n5077, n_4493, n_4494);
  not g8114 (n_4495, n5072);
  not g8115 (n_4496, n5077);
  and g8116 (n5078, n_4495, n_4496);
  not g8117 (n_4497, n5067);
  not g8118 (n_4498, n5078);
  and g8119 (n5079, n_4497, n_4498);
  not g8120 (n_4499, n5063);
  and g8121 (n5080, n_4499, n5079);
  and g8122 (n5081, n_4499, n_4497);
  not g8123 (n_4500, n5081);
  and g8124 (n5082, n5078, n_4500);
  not g8125 (n_4501, n5080);
  not g8126 (n_4502, n5082);
  and g8127 (n5083, n_4501, n_4502);
  not g8128 (n_4503, n4979);
  not g8129 (n_4504, n5083);
  and g8130 (n5084, n_4503, n_4504);
  and g8131 (n5085, n_4497, n5078);
  and g8132 (n5086, n_4499, n5085);
  and g8133 (n5087, n_4498, n_4500);
  not g8134 (n_4505, n5086);
  not g8135 (n_4506, n5087);
  and g8136 (n5088, n_4505, n_4506);
  not g8137 (n_4507, n5088);
  and g8138 (n5089, n4979, n_4507);
  and g8139 (n5090, n_4495, n5077);
  and g8140 (n5091, n5072, n_4496);
  not g8141 (n_4508, n5090);
  not g8142 (n_4509, n5091);
  and g8143 (n5092, n_4508, n_4509);
  not g8144 (n_4511, \A[991] );
  and g8145 (n5093, n_4511, \A[992] );
  not g8146 (n_4513, \A[992] );
  and g8147 (n5094, \A[991] , n_4513);
  not g8148 (n_4515, n5094);
  and g8149 (n5095, \A[993] , n_4515);
  not g8150 (n_4516, n5093);
  and g8151 (n5096, n_4516, n5095);
  and g8152 (n5097, n_4516, n_4515);
  not g8153 (n_4517, \A[993] );
  not g8154 (n_4518, n5097);
  and g8155 (n5098, n_4517, n_4518);
  not g8156 (n_4519, n5096);
  not g8157 (n_4520, n5098);
  and g8158 (n5099, n_4519, n_4520);
  not g8159 (n_4522, \A[994] );
  and g8160 (n5100, n_4522, \A[995] );
  not g8161 (n_4524, \A[995] );
  and g8162 (n5101, \A[994] , n_4524);
  not g8163 (n_4526, n5101);
  and g8164 (n5102, \A[996] , n_4526);
  not g8165 (n_4527, n5100);
  and g8166 (n5103, n_4527, n5102);
  and g8167 (n5104, n_4527, n_4526);
  not g8168 (n_4528, \A[996] );
  not g8169 (n_4529, n5104);
  and g8170 (n5105, n_4528, n_4529);
  not g8171 (n_4530, n5103);
  not g8172 (n_4531, n5105);
  and g8173 (n5106, n_4530, n_4531);
  not g8174 (n_4532, n5099);
  and g8175 (n5107, n_4532, n5106);
  not g8176 (n_4533, n5106);
  and g8177 (n5108, n5099, n_4533);
  not g8178 (n_4534, n5107);
  not g8179 (n_4535, n5108);
  and g8180 (n5109, n_4534, n_4535);
  and g8181 (n5110, \A[994] , \A[995] );
  and g8182 (n5111, \A[996] , n_4529);
  not g8183 (n_4536, n5110);
  not g8184 (n_4537, n5111);
  and g8185 (n5112, n_4536, n_4537);
  and g8186 (n5113, \A[991] , \A[992] );
  and g8187 (n5114, \A[993] , n_4518);
  not g8188 (n_4538, n5113);
  not g8189 (n_4539, n5114);
  and g8190 (n5115, n_4538, n_4539);
  not g8191 (n_4540, n5112);
  and g8192 (n5116, n_4540, n5115);
  not g8193 (n_4541, n5115);
  and g8194 (n5117, n5112, n_4541);
  not g8195 (n_4542, n5116);
  not g8196 (n_4543, n5117);
  and g8197 (n5118, n_4542, n_4543);
  and g8198 (n5119, n_4532, n_4533);
  not g8199 (n_4544, n5118);
  and g8200 (n5120, n_4544, n5119);
  and g8201 (n5121, n_4540, n_4541);
  not g8202 (n_4545, n5120);
  not g8203 (n_4546, n5121);
  and g8204 (n5122, n_4545, n_4546);
  and g8205 (n5123, n_4542, n5119);
  and g8206 (n5124, n_4543, n5123);
  not g8207 (n_4547, n5119);
  and g8208 (n5125, n_4544, n_4547);
  not g8209 (n_4548, n5124);
  not g8210 (n_4549, n5125);
  and g8211 (n5126, n_4548, n_4549);
  not g8212 (n_4550, n5122);
  not g8213 (n_4551, n5126);
  and g8214 (n5127, n_4550, n_4551);
  not g8215 (n_4552, n5109);
  not g8216 (n_4553, n5127);
  and g8217 (n5128, n_4552, n_4553);
  not g8218 (n_4556, \A[4] );
  and g8219 (n5129, \A[3] , n_4556);
  not g8220 (n_4557, \A[3] );
  and g8221 (n5130, n_4557, \A[4] );
  not g8222 (n_4559, n5130);
  and g8223 (n5131, \A[5] , n_4559);
  not g8224 (n_4560, n5129);
  and g8225 (n5132, n_4560, n5131);
  and g8226 (n5133, n_4560, n_4559);
  not g8227 (n_4561, \A[5] );
  not g8228 (n_4562, n5133);
  and g8229 (n5134, n_4561, n_4562);
  not g8230 (n_4563, n5132);
  not g8231 (n_4564, n5134);
  and g8232 (n5135, n_4563, n_4564);
  not g8233 (n_4566, \A[0] );
  and g8234 (n5136, n_4566, \A[1] );
  not g8235 (n_4568, \A[1] );
  and g8236 (n5137, \A[0] , n_4568);
  not g8237 (n_4569, n5136);
  not g8238 (n_4570, n5137);
  and g8239 (n5138, n_4569, n_4570);
  not g8240 (n_4572, \A[2] );
  not g8241 (n_4573, n5138);
  and g8242 (n5139, n_4572, n_4573);
  and g8243 (n5140, \A[2] , n_4569);
  and g8244 (n5141, n_4570, n5140);
  not g8245 (n_4575, n5141);
  and g8246 (n5142, \A[6] , n_4575);
  not g8247 (n_4576, n5139);
  and g8248 (n5143, n_4576, n5142);
  and g8249 (n5144, n_4576, n_4575);
  not g8250 (n_4577, \A[6] );
  not g8251 (n_4578, n5144);
  and g8252 (n5145, n_4577, n_4578);
  not g8253 (n_4579, n5143);
  not g8254 (n_4580, n5145);
  and g8255 (n5146, n_4579, n_4580);
  not g8256 (n_4581, n5146);
  and g8257 (n5147, n5135, n_4581);
  not g8258 (n_4582, n5135);
  and g8259 (n5148, n_4582, n_4579);
  and g8260 (n5149, n_4580, n5148);
  not g8261 (n_4584, \A[997] );
  and g8262 (n5150, n_4584, \A[998] );
  not g8263 (n_4586, \A[998] );
  and g8264 (n5151, \A[997] , n_4586);
  not g8265 (n_4588, n5151);
  and g8266 (n5152, \A[999] , n_4588);
  not g8267 (n_4589, n5150);
  and g8268 (n5153, n_4589, n5152);
  and g8269 (n5154, n_4589, n_4588);
  not g8270 (n_4590, \A[999] );
  not g8271 (n_4591, n5154);
  and g8272 (n5155, n_4590, n_4591);
  not g8273 (n_4592, n5153);
  not g8274 (n_4593, n5155);
  and g8275 (n5156, n_4592, n_4593);
  not g8276 (n_4594, n5149);
  not g8277 (n_4595, n5156);
  and g8278 (n5157, n_4594, n_4595);
  not g8279 (n_4596, n5147);
  and g8280 (n5158, n_4596, n5157);
  and g8281 (n5159, n_4596, n_4594);
  not g8282 (n_4597, n5159);
  and g8283 (n5160, n5156, n_4597);
  not g8284 (n_4598, n5158);
  not g8285 (n_4599, n5160);
  and g8286 (n5161, n_4598, n_4599);
  and g8287 (n5162, n5128, n5161);
  not g8288 (n_4600, n5128);
  not g8289 (n_4601, n5161);
  and g8290 (n5163, n_4600, n_4601);
  not g8291 (n_4602, n5162);
  not g8292 (n_4603, n5163);
  and g8293 (n5164, n_4602, n_4603);
  not g8294 (n_4604, n5092);
  not g8295 (n_4605, n5164);
  and g8296 (n5165, n_4604, n_4605);
  not g8297 (n_4606, n5089);
  and g8298 (n5166, n_4606, n5165);
  not g8299 (n_4607, n5084);
  and g8300 (n5167, n_4607, n5166);
  and g8301 (n5168, n_4607, n_4606);
  not g8302 (n_4608, n5165);
  not g8303 (n_4609, n5168);
  and g8304 (n5169, n_4608, n_4609);
  not g8305 (n_4610, n5167);
  not g8306 (n_4611, n5169);
  and g8307 (n5170, n_4610, n_4611);
  and g8308 (n5171, n_4552, n_4550);
  not g8309 (n_4612, n5171);
  and g8310 (n5172, n_4551, n_4612);
  and g8311 (n5173, n_4582, n_4581);
  and g8312 (n5174, \A[6] , n_4578);
  and g8313 (n5175, \A[3] , \A[4] );
  and g8314 (n5176, \A[5] , n_4562);
  not g8315 (n_4613, n5175);
  not g8316 (n_4614, n5176);
  and g8317 (n5177, n_4613, n_4614);
  and g8318 (n5178, \A[0] , \A[1] );
  and g8319 (n5179, \A[2] , n_4573);
  not g8320 (n_4615, n5178);
  not g8321 (n_4616, n5179);
  and g8322 (n5180, n_4615, n_4616);
  not g8323 (n_4617, n5177);
  and g8324 (n5181, n_4617, n5180);
  not g8325 (n_4618, n5180);
  and g8326 (n5182, n5177, n_4618);
  not g8327 (n_4619, n5181);
  not g8328 (n_4620, n5182);
  and g8329 (n5183, n_4619, n_4620);
  not g8330 (n_4621, n5174);
  and g8331 (n5184, n_4621, n5183);
  not g8332 (n_4622, n5173);
  and g8333 (n5185, n_4622, n5184);
  and g8334 (n5186, n_4622, n_4621);
  not g8335 (n_4623, n5183);
  not g8336 (n_4624, n5186);
  and g8337 (n5187, n_4623, n_4624);
  not g8338 (n_4625, n5185);
  not g8339 (n_4626, n5187);
  and g8340 (n5188, n_4625, n_4626);
  and g8341 (n5189, n_4595, n_4597);
  and g8342 (n5190, n5188, n5189);
  and g8343 (n5191, \A[997] , \A[998] );
  and g8344 (n5192, \A[999] , n_4591);
  not g8345 (n_4627, n5191);
  not g8346 (n_4628, n5192);
  and g8347 (n5193, n_4627, n_4628);
  not g8348 (n_4629, n5188);
  not g8349 (n_4630, n5189);
  and g8350 (n5194, n_4629, n_4630);
  not g8351 (n_4631, n5194);
  and g8352 (n5195, n5193, n_4631);
  not g8353 (n_4632, n5190);
  and g8354 (n5196, n_4632, n5195);
  and g8355 (n5197, n_4632, n_4631);
  not g8356 (n_4633, n5193);
  not g8357 (n_4634, n5197);
  and g8358 (n5198, n_4633, n_4634);
  and g8359 (n5199, n5128, n_4601);
  not g8360 (n_4635, n5198);
  and g8361 (n5200, n_4635, n5199);
  not g8362 (n_4636, n5196);
  and g8363 (n5201, n_4636, n5200);
  and g8364 (n5202, n_4636, n_4635);
  not g8365 (n_4637, n5199);
  not g8366 (n_4638, n5202);
  and g8367 (n5203, n_4637, n_4638);
  not g8368 (n_4639, n5201);
  not g8369 (n_4640, n5203);
  and g8370 (n5204, n_4639, n_4640);
  not g8371 (n_4641, n5172);
  not g8372 (n_4642, n5204);
  and g8373 (n5205, n_4641, n_4642);
  and g8374 (n5206, n_4635, n_4637);
  and g8375 (n5207, n_4636, n5206);
  and g8376 (n5208, n5199, n_4638);
  not g8377 (n_4643, n5207);
  not g8378 (n_4644, n5208);
  and g8379 (n5209, n_4643, n_4644);
  not g8380 (n_4645, n5209);
  and g8381 (n5210, n5172, n_4645);
  not g8382 (n_4646, n5205);
  not g8383 (n_4647, n5210);
  and g8384 (n5211, n_4646, n_4647);
  not g8385 (n_4648, n5170);
  and g8386 (n5212, n_4648, n5211);
  and g8387 (n5213, n_4606, n_4608);
  and g8388 (n5214, n_4607, n5213);
  and g8389 (n5215, n5165, n_4609);
  not g8390 (n_4649, n5214);
  not g8391 (n_4650, n5215);
  and g8392 (n5216, n_4649, n_4650);
  not g8393 (n_4651, n5211);
  not g8394 (n_4652, n5216);
  and g8395 (n5217, n_4651, n_4652);
  not g8396 (n_4653, n5212);
  not g8397 (n_4654, n5217);
  and g8398 (n5218, n_4653, n_4654);
  and g8399 (n5219, \A[46] , \A[47] );
  not g8400 (n_4657, \A[47] );
  and g8401 (n5220, \A[46] , n_4657);
  not g8402 (n_4658, \A[46] );
  and g8403 (n5221, n_4658, \A[47] );
  not g8404 (n_4659, n5220);
  not g8405 (n_4660, n5221);
  and g8406 (n5222, n_4659, n_4660);
  not g8407 (n_4662, n5222);
  and g8408 (n5223, \A[48] , n_4662);
  not g8409 (n_4663, n5219);
  not g8410 (n_4664, n5223);
  and g8411 (n5224, n_4663, n_4664);
  and g8412 (n5225, \A[43] , \A[44] );
  not g8413 (n_4667, \A[44] );
  and g8414 (n5226, \A[43] , n_4667);
  not g8415 (n_4668, \A[43] );
  and g8416 (n5227, n_4668, \A[44] );
  not g8417 (n_4669, n5226);
  not g8418 (n_4670, n5227);
  and g8419 (n5228, n_4669, n_4670);
  not g8420 (n_4672, n5228);
  and g8421 (n5229, \A[45] , n_4672);
  not g8422 (n_4673, n5225);
  not g8423 (n_4674, n5229);
  and g8424 (n5230, n_4673, n_4674);
  not g8425 (n_4675, n5230);
  and g8426 (n5231, n5224, n_4675);
  not g8427 (n_4676, n5224);
  and g8428 (n5232, n_4676, n5230);
  and g8429 (n5233, \A[45] , n_4669);
  and g8430 (n5234, n_4670, n5233);
  not g8431 (n_4677, \A[45] );
  and g8432 (n5235, n_4677, n_4672);
  not g8433 (n_4678, n5234);
  not g8434 (n_4679, n5235);
  and g8435 (n5236, n_4678, n_4679);
  and g8436 (n5237, \A[48] , n_4659);
  and g8437 (n5238, n_4660, n5237);
  not g8438 (n_4680, \A[48] );
  and g8439 (n5239, n_4680, n_4662);
  not g8440 (n_4681, n5238);
  not g8441 (n_4682, n5239);
  and g8442 (n5240, n_4681, n_4682);
  not g8443 (n_4683, n5236);
  not g8444 (n_4684, n5240);
  and g8445 (n5241, n_4683, n_4684);
  not g8446 (n_4685, n5232);
  and g8447 (n5242, n_4685, n5241);
  not g8448 (n_4686, n5231);
  and g8449 (n5243, n_4686, n5242);
  and g8450 (n5244, n_4686, n_4685);
  not g8451 (n_4687, n5241);
  not g8452 (n_4688, n5244);
  and g8453 (n5245, n_4687, n_4688);
  not g8454 (n_4689, n5243);
  not g8455 (n_4690, n5245);
  and g8456 (n5246, n_4689, n_4690);
  and g8457 (n5247, n_4683, n5240);
  and g8458 (n5248, n5236, n_4684);
  not g8459 (n_4691, n5247);
  not g8460 (n_4692, n5248);
  and g8461 (n5249, n_4691, n_4692);
  and g8462 (n5250, n5241, n_4688);
  and g8463 (n5251, n_4676, n_4675);
  not g8464 (n_4693, n5250);
  not g8465 (n_4694, n5251);
  and g8466 (n5252, n_4693, n_4694);
  not g8467 (n_4695, n5249);
  not g8468 (n_4696, n5252);
  and g8469 (n5253, n_4695, n_4696);
  not g8470 (n_4697, n5246);
  not g8471 (n_4698, n5253);
  and g8472 (n5254, n_4697, n_4698);
  and g8473 (n5255, n_4697, n_4696);
  and g8474 (n5256, \A[52] , \A[53] );
  not g8475 (n_4701, \A[53] );
  and g8476 (n5257, \A[52] , n_4701);
  not g8477 (n_4702, \A[52] );
  and g8478 (n5258, n_4702, \A[53] );
  not g8479 (n_4703, n5257);
  not g8480 (n_4704, n5258);
  and g8481 (n5259, n_4703, n_4704);
  not g8482 (n_4706, n5259);
  and g8483 (n5260, \A[54] , n_4706);
  not g8484 (n_4707, n5256);
  not g8485 (n_4708, n5260);
  and g8486 (n5261, n_4707, n_4708);
  and g8487 (n5262, \A[49] , \A[50] );
  not g8488 (n_4711, \A[50] );
  and g8489 (n5263, \A[49] , n_4711);
  not g8490 (n_4712, \A[49] );
  and g8491 (n5264, n_4712, \A[50] );
  not g8492 (n_4713, n5263);
  not g8493 (n_4714, n5264);
  and g8494 (n5265, n_4713, n_4714);
  not g8495 (n_4716, n5265);
  and g8496 (n5266, \A[51] , n_4716);
  not g8497 (n_4717, n5262);
  not g8498 (n_4718, n5266);
  and g8499 (n5267, n_4717, n_4718);
  not g8500 (n_4719, n5261);
  and g8501 (n5268, n_4719, n5267);
  not g8502 (n_4720, n5267);
  and g8503 (n5269, n5261, n_4720);
  not g8504 (n_4721, n5268);
  not g8505 (n_4722, n5269);
  and g8506 (n5270, n_4721, n_4722);
  and g8507 (n5271, \A[51] , n_4713);
  and g8508 (n5272, n_4714, n5271);
  not g8509 (n_4723, \A[51] );
  and g8510 (n5273, n_4723, n_4716);
  not g8511 (n_4724, n5272);
  not g8512 (n_4725, n5273);
  and g8513 (n5274, n_4724, n_4725);
  and g8514 (n5275, \A[54] , n_4703);
  and g8515 (n5276, n_4704, n5275);
  not g8516 (n_4726, \A[54] );
  and g8517 (n5277, n_4726, n_4706);
  not g8518 (n_4727, n5276);
  not g8519 (n_4728, n5277);
  and g8520 (n5278, n_4727, n_4728);
  not g8521 (n_4729, n5274);
  not g8522 (n_4730, n5278);
  and g8523 (n5279, n_4729, n_4730);
  not g8524 (n_4731, n5270);
  and g8525 (n5280, n_4731, n5279);
  and g8526 (n5281, n_4719, n_4720);
  not g8527 (n_4732, n5280);
  not g8528 (n_4733, n5281);
  and g8529 (n5282, n_4732, n_4733);
  and g8530 (n5283, n_4721, n5279);
  and g8531 (n5284, n_4722, n5283);
  not g8532 (n_4734, n5279);
  and g8533 (n5285, n_4731, n_4734);
  not g8534 (n_4735, n5284);
  not g8535 (n_4736, n5285);
  and g8536 (n5286, n_4735, n_4736);
  not g8537 (n_4737, n5282);
  not g8538 (n_4738, n5286);
  and g8539 (n5287, n_4737, n_4738);
  and g8540 (n5288, n_4729, n5278);
  and g8541 (n5289, n5274, n_4730);
  not g8542 (n_4739, n5288);
  not g8543 (n_4740, n5289);
  and g8544 (n5290, n_4739, n_4740);
  not g8545 (n_4741, n5290);
  and g8546 (n5291, n_4695, n_4741);
  not g8547 (n_4742, n5287);
  and g8548 (n5292, n_4742, n5291);
  not g8549 (n_4743, n5255);
  and g8550 (n5293, n_4743, n5292);
  and g8551 (n5294, n_4737, n_4741);
  not g8552 (n_4744, n5294);
  and g8553 (n5295, n_4738, n_4744);
  not g8554 (n_4745, n5293);
  not g8555 (n_4746, n5295);
  and g8556 (n5296, n_4745, n_4746);
  not g8561 (n_4747, n5296);
  not g8562 (n_4748, n5300);
  and g8563 (n5301, n_4747, n_4748);
  not g8564 (n_4749, n5301);
  and g8565 (n5302, n5254, n_4749);
  and g8566 (n5303, n_4745, n5295);
  and g8567 (n5304, n5293, n_4746);
  not g8568 (n_4750, n5303);
  not g8569 (n_4751, n5304);
  and g8570 (n5305, n_4750, n_4751);
  not g8571 (n_4752, n5254);
  not g8572 (n_4753, n5305);
  and g8573 (n5306, n_4752, n_4753);
  and g8574 (n5307, n_4742, n_4741);
  and g8575 (n5308, n_4695, n_4743);
  not g8576 (n_4754, n5307);
  and g8577 (n5309, n_4754, n5308);
  not g8578 (n_4755, n5308);
  and g8579 (n5310, n5307, n_4755);
  not g8580 (n_4756, n5309);
  not g8581 (n_4757, n5310);
  and g8582 (n5311, n_4756, n_4757);
  not g8583 (n_4759, \A[37] );
  and g8584 (n5312, n_4759, \A[38] );
  not g8585 (n_4761, \A[38] );
  and g8586 (n5313, \A[37] , n_4761);
  not g8587 (n_4763, n5313);
  and g8588 (n5314, \A[39] , n_4763);
  not g8589 (n_4764, n5312);
  and g8590 (n5315, n_4764, n5314);
  and g8591 (n5316, n_4764, n_4763);
  not g8592 (n_4765, \A[39] );
  not g8593 (n_4766, n5316);
  and g8594 (n5317, n_4765, n_4766);
  not g8595 (n_4767, n5315);
  not g8596 (n_4768, n5317);
  and g8597 (n5318, n_4767, n_4768);
  not g8598 (n_4770, \A[40] );
  and g8599 (n5319, n_4770, \A[41] );
  not g8600 (n_4772, \A[41] );
  and g8601 (n5320, \A[40] , n_4772);
  not g8602 (n_4774, n5320);
  and g8603 (n5321, \A[42] , n_4774);
  not g8604 (n_4775, n5319);
  and g8605 (n5322, n_4775, n5321);
  and g8606 (n5323, n_4775, n_4774);
  not g8607 (n_4776, \A[42] );
  not g8608 (n_4777, n5323);
  and g8609 (n5324, n_4776, n_4777);
  not g8610 (n_4778, n5322);
  not g8611 (n_4779, n5324);
  and g8612 (n5325, n_4778, n_4779);
  not g8613 (n_4780, n5318);
  and g8614 (n5326, n_4780, n5325);
  not g8615 (n_4781, n5325);
  and g8616 (n5327, n5318, n_4781);
  not g8617 (n_4782, n5326);
  not g8618 (n_4783, n5327);
  and g8619 (n5328, n_4782, n_4783);
  and g8620 (n5329, \A[40] , \A[41] );
  and g8621 (n5330, \A[42] , n_4777);
  not g8622 (n_4784, n5329);
  not g8623 (n_4785, n5330);
  and g8624 (n5331, n_4784, n_4785);
  and g8625 (n5332, \A[37] , \A[38] );
  and g8626 (n5333, \A[39] , n_4766);
  not g8627 (n_4786, n5332);
  not g8628 (n_4787, n5333);
  and g8629 (n5334, n_4786, n_4787);
  not g8630 (n_4788, n5331);
  and g8631 (n5335, n_4788, n5334);
  not g8632 (n_4789, n5334);
  and g8633 (n5336, n5331, n_4789);
  not g8634 (n_4790, n5335);
  not g8635 (n_4791, n5336);
  and g8636 (n5337, n_4790, n_4791);
  and g8637 (n5338, n_4780, n_4781);
  not g8638 (n_4792, n5337);
  and g8639 (n5339, n_4792, n5338);
  and g8640 (n5340, n_4788, n_4789);
  not g8641 (n_4793, n5339);
  not g8642 (n_4794, n5340);
  and g8643 (n5341, n_4793, n_4794);
  and g8644 (n5342, n_4790, n5338);
  and g8645 (n5343, n_4791, n5342);
  not g8646 (n_4795, n5338);
  and g8647 (n5344, n_4792, n_4795);
  not g8648 (n_4796, n5343);
  not g8649 (n_4797, n5344);
  and g8650 (n5345, n_4796, n_4797);
  not g8651 (n_4798, n5341);
  not g8652 (n_4799, n5345);
  and g8653 (n5346, n_4798, n_4799);
  not g8654 (n_4800, n5328);
  not g8655 (n_4801, n5346);
  and g8656 (n5347, n_4800, n_4801);
  not g8657 (n_4803, \A[31] );
  and g8658 (n5348, n_4803, \A[32] );
  not g8659 (n_4805, \A[32] );
  and g8660 (n5349, \A[31] , n_4805);
  not g8661 (n_4807, n5349);
  and g8662 (n5350, \A[33] , n_4807);
  not g8663 (n_4808, n5348);
  and g8664 (n5351, n_4808, n5350);
  and g8665 (n5352, n_4808, n_4807);
  not g8666 (n_4809, \A[33] );
  not g8667 (n_4810, n5352);
  and g8668 (n5353, n_4809, n_4810);
  not g8669 (n_4811, n5351);
  not g8670 (n_4812, n5353);
  and g8671 (n5354, n_4811, n_4812);
  not g8672 (n_4814, \A[34] );
  and g8673 (n5355, n_4814, \A[35] );
  not g8674 (n_4816, \A[35] );
  and g8675 (n5356, \A[34] , n_4816);
  not g8676 (n_4818, n5356);
  and g8677 (n5357, \A[36] , n_4818);
  not g8678 (n_4819, n5355);
  and g8679 (n5358, n_4819, n5357);
  and g8680 (n5359, n_4819, n_4818);
  not g8681 (n_4820, \A[36] );
  not g8682 (n_4821, n5359);
  and g8683 (n5360, n_4820, n_4821);
  not g8684 (n_4822, n5358);
  not g8685 (n_4823, n5360);
  and g8686 (n5361, n_4822, n_4823);
  not g8687 (n_4824, n5354);
  and g8688 (n5362, n_4824, n5361);
  not g8689 (n_4825, n5361);
  and g8690 (n5363, n5354, n_4825);
  not g8691 (n_4826, n5362);
  not g8692 (n_4827, n5363);
  and g8693 (n5364, n_4826, n_4827);
  and g8694 (n5365, \A[34] , \A[35] );
  and g8695 (n5366, \A[36] , n_4821);
  not g8696 (n_4828, n5365);
  not g8697 (n_4829, n5366);
  and g8698 (n5367, n_4828, n_4829);
  and g8699 (n5368, \A[31] , \A[32] );
  and g8700 (n5369, \A[33] , n_4810);
  not g8701 (n_4830, n5368);
  not g8702 (n_4831, n5369);
  and g8703 (n5370, n_4830, n_4831);
  not g8704 (n_4832, n5367);
  and g8705 (n5371, n_4832, n5370);
  not g8706 (n_4833, n5370);
  and g8707 (n5372, n5367, n_4833);
  not g8708 (n_4834, n5371);
  not g8709 (n_4835, n5372);
  and g8710 (n5373, n_4834, n_4835);
  and g8711 (n5374, n_4824, n_4825);
  not g8712 (n_4836, n5373);
  and g8713 (n5375, n_4836, n5374);
  and g8714 (n5376, n_4832, n_4833);
  not g8715 (n_4837, n5375);
  not g8716 (n_4838, n5376);
  and g8717 (n5377, n_4837, n_4838);
  and g8718 (n5378, n_4834, n5374);
  and g8719 (n5379, n_4835, n5378);
  not g8720 (n_4839, n5374);
  and g8721 (n5380, n_4836, n_4839);
  not g8722 (n_4840, n5379);
  not g8723 (n_4841, n5380);
  and g8724 (n5381, n_4840, n_4841);
  not g8725 (n_4842, n5377);
  not g8726 (n_4843, n5381);
  and g8727 (n5382, n_4842, n_4843);
  not g8728 (n_4844, n5364);
  not g8729 (n_4845, n5382);
  and g8730 (n5383, n_4844, n_4845);
  not g8731 (n_4846, n5347);
  and g8732 (n5384, n_4846, n5383);
  not g8733 (n_4847, n5383);
  and g8734 (n5385, n5347, n_4847);
  not g8735 (n_4848, n5384);
  not g8736 (n_4849, n5385);
  and g8737 (n5386, n_4848, n_4849);
  not g8738 (n_4850, n5311);
  not g8739 (n_4851, n5386);
  and g8740 (n5387, n_4850, n_4851);
  not g8741 (n_4852, n5306);
  and g8742 (n5388, n_4852, n5387);
  not g8743 (n_4853, n5302);
  and g8744 (n5389, n_4853, n5388);
  and g8745 (n5390, n_4853, n_4852);
  not g8746 (n_4854, n5387);
  not g8747 (n_4855, n5390);
  and g8748 (n5391, n_4854, n_4855);
  not g8749 (n_4856, n5389);
  not g8750 (n_4857, n5391);
  and g8751 (n5392, n_4856, n_4857);
  and g8752 (n5393, n_4844, n_4842);
  not g8753 (n_4858, n5393);
  and g8754 (n5394, n_4843, n_4858);
  and g8755 (n5395, n_4800, n_4844);
  and g8756 (n5396, n_4801, n5395);
  and g8757 (n5397, n_4845, n5396);
  and g8758 (n5398, n_4800, n_4798);
  not g8759 (n_4859, n5398);
  and g8760 (n5399, n_4799, n_4859);
  not g8761 (n_4860, n5397);
  and g8762 (n5400, n_4860, n5399);
  not g8763 (n_4861, n5399);
  and g8764 (n5401, n5397, n_4861);
  not g8765 (n_4862, n5400);
  not g8766 (n_4863, n5401);
  and g8767 (n5402, n_4862, n_4863);
  not g8768 (n_4864, n5394);
  not g8769 (n_4865, n5402);
  and g8770 (n5403, n_4864, n_4865);
  and g8771 (n5404, n_4860, n_4861);
  not g8776 (n_4866, n5404);
  not g8777 (n_4867, n5408);
  and g8778 (n5409, n_4866, n_4867);
  not g8779 (n_4868, n5409);
  and g8780 (n5410, n5394, n_4868);
  not g8781 (n_4869, n5403);
  not g8782 (n_4870, n5410);
  and g8783 (n5411, n_4869, n_4870);
  not g8784 (n_4871, n5392);
  and g8785 (n5412, n_4871, n5411);
  and g8786 (n5413, n_4852, n_4854);
  and g8787 (n5414, n_4853, n5413);
  and g8788 (n5415, n5387, n_4855);
  not g8789 (n_4872, n5414);
  not g8790 (n_4873, n5415);
  and g8791 (n5416, n_4872, n_4873);
  not g8792 (n_4874, n5411);
  not g8793 (n_4875, n5416);
  and g8794 (n5417, n_4874, n_4875);
  not g8795 (n_4876, n5412);
  not g8796 (n_4877, n5417);
  and g8797 (n5418, n_4876, n_4877);
  and g8798 (n5419, \A[58] , \A[59] );
  not g8799 (n_4880, \A[59] );
  and g8800 (n5420, \A[58] , n_4880);
  not g8801 (n_4881, \A[58] );
  and g8802 (n5421, n_4881, \A[59] );
  not g8803 (n_4882, n5420);
  not g8804 (n_4883, n5421);
  and g8805 (n5422, n_4882, n_4883);
  not g8806 (n_4885, n5422);
  and g8807 (n5423, \A[60] , n_4885);
  not g8808 (n_4886, n5419);
  not g8809 (n_4887, n5423);
  and g8810 (n5424, n_4886, n_4887);
  and g8811 (n5425, \A[55] , \A[56] );
  not g8812 (n_4890, \A[56] );
  and g8813 (n5426, \A[55] , n_4890);
  not g8814 (n_4891, \A[55] );
  and g8815 (n5427, n_4891, \A[56] );
  not g8816 (n_4892, n5426);
  not g8817 (n_4893, n5427);
  and g8818 (n5428, n_4892, n_4893);
  not g8819 (n_4895, n5428);
  and g8820 (n5429, \A[57] , n_4895);
  not g8821 (n_4896, n5425);
  not g8822 (n_4897, n5429);
  and g8823 (n5430, n_4896, n_4897);
  not g8824 (n_4898, n5430);
  and g8825 (n5431, n5424, n_4898);
  not g8826 (n_4899, n5424);
  and g8827 (n5432, n_4899, n5430);
  and g8828 (n5433, \A[57] , n_4892);
  and g8829 (n5434, n_4893, n5433);
  not g8830 (n_4900, \A[57] );
  and g8831 (n5435, n_4900, n_4895);
  not g8832 (n_4901, n5434);
  not g8833 (n_4902, n5435);
  and g8834 (n5436, n_4901, n_4902);
  and g8835 (n5437, \A[60] , n_4882);
  and g8836 (n5438, n_4883, n5437);
  not g8837 (n_4903, \A[60] );
  and g8838 (n5439, n_4903, n_4885);
  not g8839 (n_4904, n5438);
  not g8840 (n_4905, n5439);
  and g8841 (n5440, n_4904, n_4905);
  not g8842 (n_4906, n5436);
  not g8843 (n_4907, n5440);
  and g8844 (n5441, n_4906, n_4907);
  not g8845 (n_4908, n5432);
  and g8846 (n5442, n_4908, n5441);
  not g8847 (n_4909, n5431);
  and g8848 (n5443, n_4909, n5442);
  and g8849 (n5444, n_4909, n_4908);
  not g8850 (n_4910, n5441);
  not g8851 (n_4911, n5444);
  and g8852 (n5445, n_4910, n_4911);
  not g8853 (n_4912, n5443);
  not g8854 (n_4913, n5445);
  and g8855 (n5446, n_4912, n_4913);
  and g8856 (n5447, n_4906, n5440);
  and g8857 (n5448, n5436, n_4907);
  not g8858 (n_4914, n5447);
  not g8859 (n_4915, n5448);
  and g8860 (n5449, n_4914, n_4915);
  and g8861 (n5450, n5441, n_4911);
  and g8862 (n5451, n_4899, n_4898);
  not g8863 (n_4916, n5450);
  not g8864 (n_4917, n5451);
  and g8865 (n5452, n_4916, n_4917);
  not g8866 (n_4918, n5449);
  not g8867 (n_4919, n5452);
  and g8868 (n5453, n_4918, n_4919);
  not g8869 (n_4920, n5446);
  not g8870 (n_4921, n5453);
  and g8871 (n5454, n_4920, n_4921);
  and g8872 (n5455, n_4920, n_4919);
  and g8873 (n5456, \A[64] , \A[65] );
  not g8874 (n_4924, \A[65] );
  and g8875 (n5457, \A[64] , n_4924);
  not g8876 (n_4925, \A[64] );
  and g8877 (n5458, n_4925, \A[65] );
  not g8878 (n_4926, n5457);
  not g8879 (n_4927, n5458);
  and g8880 (n5459, n_4926, n_4927);
  not g8881 (n_4929, n5459);
  and g8882 (n5460, \A[66] , n_4929);
  not g8883 (n_4930, n5456);
  not g8884 (n_4931, n5460);
  and g8885 (n5461, n_4930, n_4931);
  and g8886 (n5462, \A[61] , \A[62] );
  not g8887 (n_4934, \A[62] );
  and g8888 (n5463, \A[61] , n_4934);
  not g8889 (n_4935, \A[61] );
  and g8890 (n5464, n_4935, \A[62] );
  not g8891 (n_4936, n5463);
  not g8892 (n_4937, n5464);
  and g8893 (n5465, n_4936, n_4937);
  not g8894 (n_4939, n5465);
  and g8895 (n5466, \A[63] , n_4939);
  not g8896 (n_4940, n5462);
  not g8897 (n_4941, n5466);
  and g8898 (n5467, n_4940, n_4941);
  not g8899 (n_4942, n5461);
  and g8900 (n5468, n_4942, n5467);
  not g8901 (n_4943, n5467);
  and g8902 (n5469, n5461, n_4943);
  not g8903 (n_4944, n5468);
  not g8904 (n_4945, n5469);
  and g8905 (n5470, n_4944, n_4945);
  and g8906 (n5471, \A[63] , n_4936);
  and g8907 (n5472, n_4937, n5471);
  not g8908 (n_4946, \A[63] );
  and g8909 (n5473, n_4946, n_4939);
  not g8910 (n_4947, n5472);
  not g8911 (n_4948, n5473);
  and g8912 (n5474, n_4947, n_4948);
  and g8913 (n5475, \A[66] , n_4926);
  and g8914 (n5476, n_4927, n5475);
  not g8915 (n_4949, \A[66] );
  and g8916 (n5477, n_4949, n_4929);
  not g8917 (n_4950, n5476);
  not g8918 (n_4951, n5477);
  and g8919 (n5478, n_4950, n_4951);
  not g8920 (n_4952, n5474);
  not g8921 (n_4953, n5478);
  and g8922 (n5479, n_4952, n_4953);
  not g8923 (n_4954, n5470);
  and g8924 (n5480, n_4954, n5479);
  and g8925 (n5481, n_4942, n_4943);
  not g8926 (n_4955, n5480);
  not g8927 (n_4956, n5481);
  and g8928 (n5482, n_4955, n_4956);
  and g8929 (n5483, n_4944, n5479);
  and g8930 (n5484, n_4945, n5483);
  not g8931 (n_4957, n5479);
  and g8932 (n5485, n_4954, n_4957);
  not g8933 (n_4958, n5484);
  not g8934 (n_4959, n5485);
  and g8935 (n5486, n_4958, n_4959);
  not g8936 (n_4960, n5482);
  not g8937 (n_4961, n5486);
  and g8938 (n5487, n_4960, n_4961);
  and g8939 (n5488, n_4952, n5478);
  and g8940 (n5489, n5474, n_4953);
  not g8941 (n_4962, n5488);
  not g8942 (n_4963, n5489);
  and g8943 (n5490, n_4962, n_4963);
  not g8944 (n_4964, n5490);
  and g8945 (n5491, n_4918, n_4964);
  not g8946 (n_4965, n5487);
  and g8947 (n5492, n_4965, n5491);
  not g8948 (n_4966, n5455);
  and g8949 (n5493, n_4966, n5492);
  and g8950 (n5494, n_4960, n_4964);
  not g8951 (n_4967, n5494);
  and g8952 (n5495, n_4961, n_4967);
  not g8953 (n_4968, n5493);
  and g8954 (n5496, n_4968, n5495);
  not g8955 (n_4969, n5495);
  and g8956 (n5497, n5493, n_4969);
  not g8957 (n_4970, n5496);
  not g8958 (n_4971, n5497);
  and g8959 (n5498, n_4970, n_4971);
  not g8960 (n_4972, n5454);
  not g8961 (n_4973, n5498);
  and g8962 (n5499, n_4972, n_4973);
  and g8963 (n5500, n_4968, n_4969);
  not g8968 (n_4974, n5500);
  not g8969 (n_4975, n5504);
  and g8970 (n5505, n_4974, n_4975);
  not g8971 (n_4976, n5505);
  and g8972 (n5506, n5454, n_4976);
  not g8973 (n_4977, n5499);
  not g8974 (n_4978, n5506);
  and g8975 (n5507, n_4977, n_4978);
  and g8976 (n5508, \A[70] , \A[71] );
  not g8977 (n_4981, \A[71] );
  and g8978 (n5509, \A[70] , n_4981);
  not g8979 (n_4982, \A[70] );
  and g8980 (n5510, n_4982, \A[71] );
  not g8981 (n_4983, n5509);
  not g8982 (n_4984, n5510);
  and g8983 (n5511, n_4983, n_4984);
  not g8984 (n_4986, n5511);
  and g8985 (n5512, \A[72] , n_4986);
  not g8986 (n_4987, n5508);
  not g8987 (n_4988, n5512);
  and g8988 (n5513, n_4987, n_4988);
  and g8989 (n5514, \A[67] , \A[68] );
  not g8990 (n_4991, \A[68] );
  and g8991 (n5515, \A[67] , n_4991);
  not g8992 (n_4992, \A[67] );
  and g8993 (n5516, n_4992, \A[68] );
  not g8994 (n_4993, n5515);
  not g8995 (n_4994, n5516);
  and g8996 (n5517, n_4993, n_4994);
  not g8997 (n_4996, n5517);
  and g8998 (n5518, \A[69] , n_4996);
  not g8999 (n_4997, n5514);
  not g9000 (n_4998, n5518);
  and g9001 (n5519, n_4997, n_4998);
  not g9002 (n_4999, n5519);
  and g9003 (n5520, n5513, n_4999);
  not g9004 (n_5000, n5513);
  and g9005 (n5521, n_5000, n5519);
  and g9006 (n5522, \A[69] , n_4993);
  and g9007 (n5523, n_4994, n5522);
  not g9008 (n_5001, \A[69] );
  and g9009 (n5524, n_5001, n_4996);
  not g9010 (n_5002, n5523);
  not g9011 (n_5003, n5524);
  and g9012 (n5525, n_5002, n_5003);
  and g9013 (n5526, \A[72] , n_4983);
  and g9014 (n5527, n_4984, n5526);
  not g9015 (n_5004, \A[72] );
  and g9016 (n5528, n_5004, n_4986);
  not g9017 (n_5005, n5527);
  not g9018 (n_5006, n5528);
  and g9019 (n5529, n_5005, n_5006);
  not g9020 (n_5007, n5525);
  not g9021 (n_5008, n5529);
  and g9022 (n5530, n_5007, n_5008);
  not g9023 (n_5009, n5521);
  and g9024 (n5531, n_5009, n5530);
  not g9025 (n_5010, n5520);
  and g9026 (n5532, n_5010, n5531);
  and g9027 (n5533, n_5010, n_5009);
  not g9028 (n_5011, n5530);
  not g9029 (n_5012, n5533);
  and g9030 (n5534, n_5011, n_5012);
  not g9031 (n_5013, n5532);
  not g9032 (n_5014, n5534);
  and g9033 (n5535, n_5013, n_5014);
  and g9034 (n5536, n_5007, n5529);
  and g9035 (n5537, n5525, n_5008);
  not g9036 (n_5015, n5536);
  not g9037 (n_5016, n5537);
  and g9038 (n5538, n_5015, n_5016);
  and g9039 (n5539, n5530, n_5012);
  and g9040 (n5540, n_5000, n_4999);
  not g9041 (n_5017, n5539);
  not g9042 (n_5018, n5540);
  and g9043 (n5541, n_5017, n_5018);
  not g9044 (n_5019, n5538);
  not g9045 (n_5020, n5541);
  and g9046 (n5542, n_5019, n_5020);
  not g9047 (n_5021, n5535);
  not g9048 (n_5022, n5542);
  and g9049 (n5543, n_5021, n_5022);
  and g9050 (n5544, n_5021, n_5020);
  and g9051 (n5545, \A[76] , \A[77] );
  not g9052 (n_5025, \A[77] );
  and g9053 (n5546, \A[76] , n_5025);
  not g9054 (n_5026, \A[76] );
  and g9055 (n5547, n_5026, \A[77] );
  not g9056 (n_5027, n5546);
  not g9057 (n_5028, n5547);
  and g9058 (n5548, n_5027, n_5028);
  not g9059 (n_5030, n5548);
  and g9060 (n5549, \A[78] , n_5030);
  not g9061 (n_5031, n5545);
  not g9062 (n_5032, n5549);
  and g9063 (n5550, n_5031, n_5032);
  and g9064 (n5551, \A[73] , \A[74] );
  not g9065 (n_5035, \A[74] );
  and g9066 (n5552, \A[73] , n_5035);
  not g9067 (n_5036, \A[73] );
  and g9068 (n5553, n_5036, \A[74] );
  not g9069 (n_5037, n5552);
  not g9070 (n_5038, n5553);
  and g9071 (n5554, n_5037, n_5038);
  not g9072 (n_5040, n5554);
  and g9073 (n5555, \A[75] , n_5040);
  not g9074 (n_5041, n5551);
  not g9075 (n_5042, n5555);
  and g9076 (n5556, n_5041, n_5042);
  not g9077 (n_5043, n5550);
  and g9078 (n5557, n_5043, n5556);
  not g9079 (n_5044, n5556);
  and g9080 (n5558, n5550, n_5044);
  not g9081 (n_5045, n5557);
  not g9082 (n_5046, n5558);
  and g9083 (n5559, n_5045, n_5046);
  and g9084 (n5560, \A[75] , n_5037);
  and g9085 (n5561, n_5038, n5560);
  not g9086 (n_5047, \A[75] );
  and g9087 (n5562, n_5047, n_5040);
  not g9088 (n_5048, n5561);
  not g9089 (n_5049, n5562);
  and g9090 (n5563, n_5048, n_5049);
  and g9091 (n5564, \A[78] , n_5027);
  and g9092 (n5565, n_5028, n5564);
  not g9093 (n_5050, \A[78] );
  and g9094 (n5566, n_5050, n_5030);
  not g9095 (n_5051, n5565);
  not g9096 (n_5052, n5566);
  and g9097 (n5567, n_5051, n_5052);
  not g9098 (n_5053, n5563);
  not g9099 (n_5054, n5567);
  and g9100 (n5568, n_5053, n_5054);
  not g9101 (n_5055, n5559);
  and g9102 (n5569, n_5055, n5568);
  and g9103 (n5570, n_5043, n_5044);
  not g9104 (n_5056, n5569);
  not g9105 (n_5057, n5570);
  and g9106 (n5571, n_5056, n_5057);
  and g9107 (n5572, n_5045, n5568);
  and g9108 (n5573, n_5046, n5572);
  not g9109 (n_5058, n5568);
  and g9110 (n5574, n_5055, n_5058);
  not g9111 (n_5059, n5573);
  not g9112 (n_5060, n5574);
  and g9113 (n5575, n_5059, n_5060);
  not g9114 (n_5061, n5571);
  not g9115 (n_5062, n5575);
  and g9116 (n5576, n_5061, n_5062);
  and g9117 (n5577, n_5053, n5567);
  and g9118 (n5578, n5563, n_5054);
  not g9119 (n_5063, n5577);
  not g9120 (n_5064, n5578);
  and g9121 (n5579, n_5063, n_5064);
  not g9122 (n_5065, n5579);
  and g9123 (n5580, n_5019, n_5065);
  not g9124 (n_5066, n5576);
  and g9125 (n5581, n_5066, n5580);
  not g9126 (n_5067, n5544);
  and g9127 (n5582, n_5067, n5581);
  and g9128 (n5583, n_5061, n_5065);
  not g9129 (n_5068, n5583);
  and g9130 (n5584, n_5062, n_5068);
  not g9131 (n_5069, n5582);
  not g9132 (n_5070, n5584);
  and g9133 (n5585, n_5069, n_5070);
  not g9138 (n_5071, n5585);
  not g9139 (n_5072, n5589);
  and g9140 (n5590, n_5071, n_5072);
  not g9141 (n_5073, n5590);
  and g9142 (n5591, n5543, n_5073);
  and g9143 (n5592, n_5069, n5584);
  and g9144 (n5593, n5582, n_5070);
  not g9145 (n_5074, n5592);
  not g9146 (n_5075, n5593);
  and g9147 (n5594, n_5074, n_5075);
  not g9148 (n_5076, n5543);
  not g9149 (n_5077, n5594);
  and g9150 (n5595, n_5076, n_5077);
  and g9151 (n5596, n_5066, n_5065);
  and g9152 (n5597, n_5019, n_5067);
  not g9153 (n_5078, n5596);
  and g9154 (n5598, n_5078, n5597);
  not g9155 (n_5079, n5597);
  and g9156 (n5599, n5596, n_5079);
  not g9157 (n_5080, n5598);
  not g9158 (n_5081, n5599);
  and g9159 (n5600, n_5080, n_5081);
  and g9160 (n5601, n_4965, n_4964);
  and g9161 (n5602, n_4918, n_4966);
  not g9162 (n_5082, n5601);
  and g9163 (n5603, n_5082, n5602);
  not g9164 (n_5083, n5602);
  and g9165 (n5604, n5601, n_5083);
  not g9166 (n_5084, n5603);
  not g9167 (n_5085, n5604);
  and g9168 (n5605, n_5084, n_5085);
  not g9169 (n_5086, n5600);
  not g9170 (n_5087, n5605);
  and g9171 (n5606, n_5086, n_5087);
  not g9172 (n_5088, n5595);
  not g9173 (n_5089, n5606);
  and g9174 (n5607, n_5088, n_5089);
  not g9175 (n_5090, n5591);
  and g9176 (n5608, n_5090, n5607);
  and g9177 (n5609, n_5090, n_5088);
  not g9178 (n_5091, n5609);
  and g9179 (n5610, n5606, n_5091);
  not g9180 (n_5092, n5608);
  not g9181 (n_5093, n5610);
  and g9182 (n5611, n_5092, n_5093);
  not g9183 (n_5094, n5507);
  not g9184 (n_5095, n5611);
  and g9185 (n5612, n_5094, n_5095);
  and g9186 (n5613, n_5088, n5606);
  and g9187 (n5614, n_5090, n5613);
  and g9188 (n5615, n_5089, n_5091);
  not g9189 (n_5096, n5614);
  not g9190 (n_5097, n5615);
  and g9191 (n5616, n_5096, n_5097);
  not g9192 (n_5098, n5616);
  and g9193 (n5617, n5507, n_5098);
  and g9194 (n5618, n_5086, n5605);
  and g9195 (n5619, n5600, n_5087);
  not g9196 (n_5099, n5618);
  not g9197 (n_5100, n5619);
  and g9198 (n5620, n_5099, n_5100);
  and g9199 (n5621, n_4850, n5386);
  and g9200 (n5622, n5311, n_4851);
  not g9201 (n_5101, n5621);
  not g9202 (n_5102, n5622);
  and g9203 (n5623, n_5101, n_5102);
  not g9204 (n_5103, n5620);
  not g9205 (n_5104, n5623);
  and g9206 (n5624, n_5103, n_5104);
  not g9207 (n_5105, n5617);
  not g9208 (n_5106, n5624);
  and g9209 (n5625, n_5105, n_5106);
  not g9210 (n_5107, n5612);
  and g9211 (n5626, n_5107, n5625);
  and g9212 (n5627, n_5107, n_5105);
  not g9213 (n_5108, n5627);
  and g9214 (n5628, n5624, n_5108);
  not g9215 (n_5109, n5626);
  not g9216 (n_5110, n5628);
  and g9217 (n5629, n_5109, n_5110);
  not g9218 (n_5111, n5418);
  not g9219 (n_5112, n5629);
  and g9220 (n5630, n_5111, n_5112);
  and g9221 (n5631, n_5105, n5624);
  and g9222 (n5632, n_5107, n5631);
  and g9223 (n5633, n_5106, n_5108);
  not g9224 (n_5113, n5632);
  not g9225 (n_5114, n5633);
  and g9226 (n5634, n_5113, n_5114);
  not g9227 (n_5115, n5634);
  and g9228 (n5635, n5418, n_5115);
  and g9229 (n5636, n_5103, n5623);
  and g9230 (n5637, n5620, n_5104);
  not g9231 (n_5116, n5636);
  not g9232 (n_5117, n5637);
  and g9233 (n5638, n_5116, n_5117);
  and g9234 (n5639, n_4604, n5164);
  and g9235 (n5640, n_4508, n_4605);
  and g9236 (n5641, n_4509, n5640);
  not g9237 (n_5118, n5639);
  not g9238 (n_5119, n5641);
  and g9239 (n5642, n_5118, n_5119);
  not g9240 (n_5120, n5638);
  not g9241 (n_5121, n5642);
  and g9242 (n5643, n_5120, n_5121);
  not g9243 (n_5122, n5635);
  not g9244 (n_5123, n5643);
  and g9245 (n5644, n_5122, n_5123);
  not g9246 (n_5124, n5630);
  and g9247 (n5645, n_5124, n5644);
  and g9248 (n5646, n_5124, n_5122);
  not g9249 (n_5125, n5646);
  and g9250 (n5647, n5643, n_5125);
  not g9251 (n_5126, n5645);
  not g9252 (n_5127, n5647);
  and g9253 (n5648, n_5126, n_5127);
  not g9254 (n_5128, n5218);
  not g9255 (n_5129, n5648);
  and g9256 (n5649, n_5128, n_5129);
  and g9257 (n5650, n_5122, n5643);
  and g9258 (n5651, n_5124, n5650);
  and g9259 (n5652, n_5123, n_5125);
  not g9260 (n_5130, n5651);
  not g9261 (n_5131, n5652);
  and g9262 (n5653, n_5130, n_5131);
  not g9263 (n_5132, n5653);
  and g9264 (n5654, n5218, n_5132);
  and g9265 (n5655, n_5120, n5642);
  and g9266 (n5656, n5638, n_5121);
  not g9267 (n_5133, n5655);
  not g9268 (n_5134, n5656);
  and g9269 (n5657, n_5133, n_5134);
  and g9270 (n5658, n_4235, n4827);
  and g9271 (n5659, n4674, n_4236);
  not g9272 (n_5135, n5658);
  not g9273 (n_5136, n5659);
  and g9274 (n5660, n_5135, n_5136);
  not g9275 (n_5137, n5657);
  not g9276 (n_5138, n5660);
  and g9277 (n5661, n_5137, n_5138);
  not g9278 (n_5139, n5654);
  not g9279 (n_5140, n5661);
  and g9280 (n5662, n_5139, n_5140);
  not g9281 (n_5141, n5649);
  and g9282 (n5663, n_5141, n5662);
  and g9283 (n5664, n_5141, n_5139);
  not g9284 (n_5142, n5664);
  and g9285 (n5665, n5661, n_5142);
  not g9286 (n_5143, n5663);
  not g9287 (n_5144, n5665);
  and g9288 (n5666, n_5143, n_5144);
  not g9289 (n_5145, n4890);
  not g9290 (n_5146, n5666);
  and g9291 (n5667, n_5145, n_5146);
  and g9292 (n5668, n_5139, n5661);
  and g9293 (n5669, n_5141, n5668);
  and g9294 (n5670, n_5140, n_5142);
  not g9295 (n_5147, n5669);
  not g9296 (n_5148, n5670);
  and g9297 (n5671, n_5147, n_5148);
  not g9298 (n_5149, n5671);
  and g9299 (n5672, n4890, n_5149);
  and g9300 (n5673, n_5137, n5660);
  and g9301 (n5674, n_5133, n_5138);
  and g9302 (n5675, n_5134, n5674);
  not g9303 (n_5150, n5673);
  not g9304 (n_5151, n5675);
  and g9305 (n5676, n_5150, n_5151);
  not g9306 (n_5153, \A[937] );
  and g9307 (n5677, n_5153, \A[938] );
  not g9308 (n_5155, \A[938] );
  and g9309 (n5678, \A[937] , n_5155);
  not g9310 (n_5157, n5678);
  and g9311 (n5679, \A[939] , n_5157);
  not g9312 (n_5158, n5677);
  and g9313 (n5680, n_5158, n5679);
  and g9314 (n5681, n_5158, n_5157);
  not g9315 (n_5159, \A[939] );
  not g9316 (n_5160, n5681);
  and g9317 (n5682, n_5159, n_5160);
  not g9318 (n_5161, n5680);
  not g9319 (n_5162, n5682);
  and g9320 (n5683, n_5161, n_5162);
  not g9321 (n_5164, \A[940] );
  and g9322 (n5684, n_5164, \A[941] );
  not g9323 (n_5166, \A[941] );
  and g9324 (n5685, \A[940] , n_5166);
  not g9325 (n_5168, n5685);
  and g9326 (n5686, \A[942] , n_5168);
  not g9327 (n_5169, n5684);
  and g9328 (n5687, n_5169, n5686);
  and g9329 (n5688, n_5169, n_5168);
  not g9330 (n_5170, \A[942] );
  not g9331 (n_5171, n5688);
  and g9332 (n5689, n_5170, n_5171);
  not g9333 (n_5172, n5687);
  not g9334 (n_5173, n5689);
  and g9335 (n5690, n_5172, n_5173);
  not g9336 (n_5174, n5683);
  and g9337 (n5691, n_5174, n5690);
  not g9338 (n_5175, n5690);
  and g9339 (n5692, n5683, n_5175);
  not g9340 (n_5176, n5691);
  not g9341 (n_5177, n5692);
  and g9342 (n5693, n_5176, n_5177);
  and g9343 (n5694, \A[940] , \A[941] );
  and g9344 (n5695, \A[942] , n_5171);
  not g9345 (n_5178, n5694);
  not g9346 (n_5179, n5695);
  and g9347 (n5696, n_5178, n_5179);
  and g9348 (n5697, \A[937] , \A[938] );
  and g9349 (n5698, \A[939] , n_5160);
  not g9350 (n_5180, n5697);
  not g9351 (n_5181, n5698);
  and g9352 (n5699, n_5180, n_5181);
  not g9353 (n_5182, n5696);
  and g9354 (n5700, n_5182, n5699);
  not g9355 (n_5183, n5699);
  and g9356 (n5701, n5696, n_5183);
  not g9357 (n_5184, n5700);
  not g9358 (n_5185, n5701);
  and g9359 (n5702, n_5184, n_5185);
  and g9360 (n5703, n_5174, n_5175);
  not g9361 (n_5186, n5702);
  and g9362 (n5704, n_5186, n5703);
  and g9363 (n5705, n_5182, n_5183);
  not g9364 (n_5187, n5704);
  not g9365 (n_5188, n5705);
  and g9366 (n5706, n_5187, n_5188);
  and g9367 (n5707, n_5184, n5703);
  and g9368 (n5708, n_5185, n5707);
  not g9369 (n_5189, n5703);
  and g9370 (n5709, n_5186, n_5189);
  not g9371 (n_5190, n5708);
  not g9372 (n_5191, n5709);
  and g9373 (n5710, n_5190, n_5191);
  not g9374 (n_5192, n5706);
  not g9375 (n_5193, n5710);
  and g9376 (n5711, n_5192, n_5193);
  not g9377 (n_5194, n5693);
  not g9378 (n_5195, n5711);
  and g9379 (n5712, n_5194, n_5195);
  not g9380 (n_5197, \A[931] );
  and g9381 (n5713, n_5197, \A[932] );
  not g9382 (n_5199, \A[932] );
  and g9383 (n5714, \A[931] , n_5199);
  not g9384 (n_5201, n5714);
  and g9385 (n5715, \A[933] , n_5201);
  not g9386 (n_5202, n5713);
  and g9387 (n5716, n_5202, n5715);
  and g9388 (n5717, n_5202, n_5201);
  not g9389 (n_5203, \A[933] );
  not g9390 (n_5204, n5717);
  and g9391 (n5718, n_5203, n_5204);
  not g9392 (n_5205, n5716);
  not g9393 (n_5206, n5718);
  and g9394 (n5719, n_5205, n_5206);
  not g9395 (n_5208, \A[934] );
  and g9396 (n5720, n_5208, \A[935] );
  not g9397 (n_5210, \A[935] );
  and g9398 (n5721, \A[934] , n_5210);
  not g9399 (n_5212, n5721);
  and g9400 (n5722, \A[936] , n_5212);
  not g9401 (n_5213, n5720);
  and g9402 (n5723, n_5213, n5722);
  and g9403 (n5724, n_5213, n_5212);
  not g9404 (n_5214, \A[936] );
  not g9405 (n_5215, n5724);
  and g9406 (n5725, n_5214, n_5215);
  not g9407 (n_5216, n5723);
  not g9408 (n_5217, n5725);
  and g9409 (n5726, n_5216, n_5217);
  not g9410 (n_5218, n5719);
  and g9411 (n5727, n_5218, n5726);
  not g9412 (n_5219, n5726);
  and g9413 (n5728, n5719, n_5219);
  not g9414 (n_5220, n5727);
  not g9415 (n_5221, n5728);
  and g9416 (n5729, n_5220, n_5221);
  and g9417 (n5730, \A[934] , \A[935] );
  and g9418 (n5731, \A[936] , n_5215);
  not g9419 (n_5222, n5730);
  not g9420 (n_5223, n5731);
  and g9421 (n5732, n_5222, n_5223);
  and g9422 (n5733, \A[931] , \A[932] );
  and g9423 (n5734, \A[933] , n_5204);
  not g9424 (n_5224, n5733);
  not g9425 (n_5225, n5734);
  and g9426 (n5735, n_5224, n_5225);
  not g9427 (n_5226, n5732);
  and g9428 (n5736, n_5226, n5735);
  not g9429 (n_5227, n5735);
  and g9430 (n5737, n5732, n_5227);
  not g9431 (n_5228, n5736);
  not g9432 (n_5229, n5737);
  and g9433 (n5738, n_5228, n_5229);
  and g9434 (n5739, n_5218, n_5219);
  not g9435 (n_5230, n5738);
  and g9436 (n5740, n_5230, n5739);
  and g9437 (n5741, n_5226, n_5227);
  not g9438 (n_5231, n5740);
  not g9439 (n_5232, n5741);
  and g9440 (n5742, n_5231, n_5232);
  and g9441 (n5743, n_5228, n5739);
  and g9442 (n5744, n_5229, n5743);
  not g9443 (n_5233, n5739);
  and g9444 (n5745, n_5230, n_5233);
  not g9445 (n_5234, n5744);
  not g9446 (n_5235, n5745);
  and g9447 (n5746, n_5234, n_5235);
  not g9448 (n_5236, n5742);
  not g9449 (n_5237, n5746);
  and g9450 (n5747, n_5236, n_5237);
  not g9451 (n_5238, n5729);
  not g9452 (n_5239, n5747);
  and g9453 (n5748, n_5238, n_5239);
  not g9454 (n_5240, n5712);
  and g9455 (n5749, n_5240, n5748);
  not g9456 (n_5241, n5748);
  and g9457 (n5750, n5712, n_5241);
  not g9458 (n_5242, n5749);
  not g9459 (n_5243, n5750);
  and g9460 (n5751, n_5242, n_5243);
  not g9461 (n_5245, \A[925] );
  and g9462 (n5752, n_5245, \A[926] );
  not g9463 (n_5247, \A[926] );
  and g9464 (n5753, \A[925] , n_5247);
  not g9465 (n_5249, n5753);
  and g9466 (n5754, \A[927] , n_5249);
  not g9467 (n_5250, n5752);
  and g9468 (n5755, n_5250, n5754);
  and g9469 (n5756, n_5250, n_5249);
  not g9470 (n_5251, \A[927] );
  not g9471 (n_5252, n5756);
  and g9472 (n5757, n_5251, n_5252);
  not g9473 (n_5253, n5755);
  not g9474 (n_5254, n5757);
  and g9475 (n5758, n_5253, n_5254);
  not g9476 (n_5256, \A[928] );
  and g9477 (n5759, n_5256, \A[929] );
  not g9478 (n_5258, \A[929] );
  and g9479 (n5760, \A[928] , n_5258);
  not g9480 (n_5260, n5760);
  and g9481 (n5761, \A[930] , n_5260);
  not g9482 (n_5261, n5759);
  and g9483 (n5762, n_5261, n5761);
  and g9484 (n5763, n_5261, n_5260);
  not g9485 (n_5262, \A[930] );
  not g9486 (n_5263, n5763);
  and g9487 (n5764, n_5262, n_5263);
  not g9488 (n_5264, n5762);
  not g9489 (n_5265, n5764);
  and g9490 (n5765, n_5264, n_5265);
  not g9491 (n_5266, n5758);
  and g9492 (n5766, n_5266, n5765);
  not g9493 (n_5267, n5765);
  and g9494 (n5767, n5758, n_5267);
  not g9495 (n_5268, n5766);
  not g9496 (n_5269, n5767);
  and g9497 (n5768, n_5268, n_5269);
  and g9498 (n5769, \A[928] , \A[929] );
  and g9499 (n5770, \A[930] , n_5263);
  not g9500 (n_5270, n5769);
  not g9501 (n_5271, n5770);
  and g9502 (n5771, n_5270, n_5271);
  and g9503 (n5772, \A[925] , \A[926] );
  and g9504 (n5773, \A[927] , n_5252);
  not g9505 (n_5272, n5772);
  not g9506 (n_5273, n5773);
  and g9507 (n5774, n_5272, n_5273);
  not g9508 (n_5274, n5771);
  and g9509 (n5775, n_5274, n5774);
  not g9510 (n_5275, n5774);
  and g9511 (n5776, n5771, n_5275);
  not g9512 (n_5276, n5775);
  not g9513 (n_5277, n5776);
  and g9514 (n5777, n_5276, n_5277);
  and g9515 (n5778, n_5266, n_5267);
  not g9516 (n_5278, n5777);
  and g9517 (n5779, n_5278, n5778);
  and g9518 (n5780, n_5274, n_5275);
  not g9519 (n_5279, n5779);
  not g9520 (n_5280, n5780);
  and g9521 (n5781, n_5279, n_5280);
  and g9522 (n5782, n_5276, n5778);
  and g9523 (n5783, n_5277, n5782);
  not g9524 (n_5281, n5778);
  and g9525 (n5784, n_5278, n_5281);
  not g9526 (n_5282, n5783);
  not g9527 (n_5283, n5784);
  and g9528 (n5785, n_5282, n_5283);
  not g9529 (n_5284, n5781);
  not g9530 (n_5285, n5785);
  and g9531 (n5786, n_5284, n_5285);
  not g9532 (n_5286, n5768);
  not g9533 (n_5287, n5786);
  and g9534 (n5787, n_5286, n_5287);
  not g9535 (n_5289, \A[919] );
  and g9536 (n5788, n_5289, \A[920] );
  not g9537 (n_5291, \A[920] );
  and g9538 (n5789, \A[919] , n_5291);
  not g9539 (n_5293, n5789);
  and g9540 (n5790, \A[921] , n_5293);
  not g9541 (n_5294, n5788);
  and g9542 (n5791, n_5294, n5790);
  and g9543 (n5792, n_5294, n_5293);
  not g9544 (n_5295, \A[921] );
  not g9545 (n_5296, n5792);
  and g9546 (n5793, n_5295, n_5296);
  not g9547 (n_5297, n5791);
  not g9548 (n_5298, n5793);
  and g9549 (n5794, n_5297, n_5298);
  not g9550 (n_5300, \A[922] );
  and g9551 (n5795, n_5300, \A[923] );
  not g9552 (n_5302, \A[923] );
  and g9553 (n5796, \A[922] , n_5302);
  not g9554 (n_5304, n5796);
  and g9555 (n5797, \A[924] , n_5304);
  not g9556 (n_5305, n5795);
  and g9557 (n5798, n_5305, n5797);
  and g9558 (n5799, n_5305, n_5304);
  not g9559 (n_5306, \A[924] );
  not g9560 (n_5307, n5799);
  and g9561 (n5800, n_5306, n_5307);
  not g9562 (n_5308, n5798);
  not g9563 (n_5309, n5800);
  and g9564 (n5801, n_5308, n_5309);
  not g9565 (n_5310, n5794);
  and g9566 (n5802, n_5310, n5801);
  not g9567 (n_5311, n5801);
  and g9568 (n5803, n5794, n_5311);
  not g9569 (n_5312, n5802);
  not g9570 (n_5313, n5803);
  and g9571 (n5804, n_5312, n_5313);
  and g9572 (n5805, \A[922] , \A[923] );
  and g9573 (n5806, \A[924] , n_5307);
  not g9574 (n_5314, n5805);
  not g9575 (n_5315, n5806);
  and g9576 (n5807, n_5314, n_5315);
  and g9577 (n5808, \A[919] , \A[920] );
  and g9578 (n5809, \A[921] , n_5296);
  not g9579 (n_5316, n5808);
  not g9580 (n_5317, n5809);
  and g9581 (n5810, n_5316, n_5317);
  not g9582 (n_5318, n5807);
  and g9583 (n5811, n_5318, n5810);
  not g9584 (n_5319, n5810);
  and g9585 (n5812, n5807, n_5319);
  not g9586 (n_5320, n5811);
  not g9587 (n_5321, n5812);
  and g9588 (n5813, n_5320, n_5321);
  and g9589 (n5814, n_5310, n_5311);
  not g9590 (n_5322, n5813);
  and g9591 (n5815, n_5322, n5814);
  and g9592 (n5816, n_5318, n_5319);
  not g9593 (n_5323, n5815);
  not g9594 (n_5324, n5816);
  and g9595 (n5817, n_5323, n_5324);
  and g9596 (n5818, n_5320, n5814);
  and g9597 (n5819, n_5321, n5818);
  not g9598 (n_5325, n5814);
  and g9599 (n5820, n_5322, n_5325);
  not g9600 (n_5326, n5819);
  not g9601 (n_5327, n5820);
  and g9602 (n5821, n_5326, n_5327);
  not g9603 (n_5328, n5817);
  not g9604 (n_5329, n5821);
  and g9605 (n5822, n_5328, n_5329);
  not g9606 (n_5330, n5804);
  not g9607 (n_5331, n5822);
  and g9608 (n5823, n_5330, n_5331);
  not g9609 (n_5332, n5787);
  and g9610 (n5824, n_5332, n5823);
  not g9611 (n_5333, n5823);
  and g9612 (n5825, n5787, n_5333);
  not g9613 (n_5334, n5824);
  not g9614 (n_5335, n5825);
  and g9615 (n5826, n_5334, n_5335);
  not g9616 (n_5336, n5751);
  and g9617 (n5827, n_5336, n5826);
  not g9618 (n_5337, n5826);
  and g9619 (n5828, n5751, n_5337);
  not g9620 (n_5338, n5827);
  not g9621 (n_5339, n5828);
  and g9622 (n5829, n_5338, n_5339);
  not g9623 (n_5341, \A[913] );
  and g9624 (n5830, n_5341, \A[914] );
  not g9625 (n_5343, \A[914] );
  and g9626 (n5831, \A[913] , n_5343);
  not g9627 (n_5345, n5831);
  and g9628 (n5832, \A[915] , n_5345);
  not g9629 (n_5346, n5830);
  and g9630 (n5833, n_5346, n5832);
  and g9631 (n5834, n_5346, n_5345);
  not g9632 (n_5347, \A[915] );
  not g9633 (n_5348, n5834);
  and g9634 (n5835, n_5347, n_5348);
  not g9635 (n_5349, n5833);
  not g9636 (n_5350, n5835);
  and g9637 (n5836, n_5349, n_5350);
  not g9638 (n_5352, \A[916] );
  and g9639 (n5837, n_5352, \A[917] );
  not g9640 (n_5354, \A[917] );
  and g9641 (n5838, \A[916] , n_5354);
  not g9642 (n_5356, n5838);
  and g9643 (n5839, \A[918] , n_5356);
  not g9644 (n_5357, n5837);
  and g9645 (n5840, n_5357, n5839);
  and g9646 (n5841, n_5357, n_5356);
  not g9647 (n_5358, \A[918] );
  not g9648 (n_5359, n5841);
  and g9649 (n5842, n_5358, n_5359);
  not g9650 (n_5360, n5840);
  not g9651 (n_5361, n5842);
  and g9652 (n5843, n_5360, n_5361);
  not g9653 (n_5362, n5836);
  and g9654 (n5844, n_5362, n5843);
  not g9655 (n_5363, n5843);
  and g9656 (n5845, n5836, n_5363);
  not g9657 (n_5364, n5844);
  not g9658 (n_5365, n5845);
  and g9659 (n5846, n_5364, n_5365);
  and g9660 (n5847, \A[916] , \A[917] );
  and g9661 (n5848, \A[918] , n_5359);
  not g9662 (n_5366, n5847);
  not g9663 (n_5367, n5848);
  and g9664 (n5849, n_5366, n_5367);
  and g9665 (n5850, \A[913] , \A[914] );
  and g9666 (n5851, \A[915] , n_5348);
  not g9667 (n_5368, n5850);
  not g9668 (n_5369, n5851);
  and g9669 (n5852, n_5368, n_5369);
  not g9670 (n_5370, n5849);
  and g9671 (n5853, n_5370, n5852);
  not g9672 (n_5371, n5852);
  and g9673 (n5854, n5849, n_5371);
  not g9674 (n_5372, n5853);
  not g9675 (n_5373, n5854);
  and g9676 (n5855, n_5372, n_5373);
  and g9677 (n5856, n_5362, n_5363);
  not g9678 (n_5374, n5855);
  and g9679 (n5857, n_5374, n5856);
  and g9680 (n5858, n_5370, n_5371);
  not g9681 (n_5375, n5857);
  not g9682 (n_5376, n5858);
  and g9683 (n5859, n_5375, n_5376);
  and g9684 (n5860, n_5372, n5856);
  and g9685 (n5861, n_5373, n5860);
  not g9686 (n_5377, n5856);
  and g9687 (n5862, n_5374, n_5377);
  not g9688 (n_5378, n5861);
  not g9689 (n_5379, n5862);
  and g9690 (n5863, n_5378, n_5379);
  not g9691 (n_5380, n5859);
  not g9692 (n_5381, n5863);
  and g9693 (n5864, n_5380, n_5381);
  not g9694 (n_5382, n5846);
  not g9695 (n_5383, n5864);
  and g9696 (n5865, n_5382, n_5383);
  not g9697 (n_5385, \A[907] );
  and g9698 (n5866, n_5385, \A[908] );
  not g9699 (n_5387, \A[908] );
  and g9700 (n5867, \A[907] , n_5387);
  not g9701 (n_5389, n5867);
  and g9702 (n5868, \A[909] , n_5389);
  not g9703 (n_5390, n5866);
  and g9704 (n5869, n_5390, n5868);
  and g9705 (n5870, n_5390, n_5389);
  not g9706 (n_5391, \A[909] );
  not g9707 (n_5392, n5870);
  and g9708 (n5871, n_5391, n_5392);
  not g9709 (n_5393, n5869);
  not g9710 (n_5394, n5871);
  and g9711 (n5872, n_5393, n_5394);
  not g9712 (n_5396, \A[910] );
  and g9713 (n5873, n_5396, \A[911] );
  not g9714 (n_5398, \A[911] );
  and g9715 (n5874, \A[910] , n_5398);
  not g9716 (n_5400, n5874);
  and g9717 (n5875, \A[912] , n_5400);
  not g9718 (n_5401, n5873);
  and g9719 (n5876, n_5401, n5875);
  and g9720 (n5877, n_5401, n_5400);
  not g9721 (n_5402, \A[912] );
  not g9722 (n_5403, n5877);
  and g9723 (n5878, n_5402, n_5403);
  not g9724 (n_5404, n5876);
  not g9725 (n_5405, n5878);
  and g9726 (n5879, n_5404, n_5405);
  not g9727 (n_5406, n5872);
  and g9728 (n5880, n_5406, n5879);
  not g9729 (n_5407, n5879);
  and g9730 (n5881, n5872, n_5407);
  not g9731 (n_5408, n5880);
  not g9732 (n_5409, n5881);
  and g9733 (n5882, n_5408, n_5409);
  and g9734 (n5883, \A[910] , \A[911] );
  and g9735 (n5884, \A[912] , n_5403);
  not g9736 (n_5410, n5883);
  not g9737 (n_5411, n5884);
  and g9738 (n5885, n_5410, n_5411);
  and g9739 (n5886, \A[907] , \A[908] );
  and g9740 (n5887, \A[909] , n_5392);
  not g9741 (n_5412, n5886);
  not g9742 (n_5413, n5887);
  and g9743 (n5888, n_5412, n_5413);
  not g9744 (n_5414, n5885);
  and g9745 (n5889, n_5414, n5888);
  not g9746 (n_5415, n5888);
  and g9747 (n5890, n5885, n_5415);
  not g9748 (n_5416, n5889);
  not g9749 (n_5417, n5890);
  and g9750 (n5891, n_5416, n_5417);
  and g9751 (n5892, n_5406, n_5407);
  not g9752 (n_5418, n5891);
  and g9753 (n5893, n_5418, n5892);
  and g9754 (n5894, n_5414, n_5415);
  not g9755 (n_5419, n5893);
  not g9756 (n_5420, n5894);
  and g9757 (n5895, n_5419, n_5420);
  and g9758 (n5896, n_5416, n5892);
  and g9759 (n5897, n_5417, n5896);
  not g9760 (n_5421, n5892);
  and g9761 (n5898, n_5418, n_5421);
  not g9762 (n_5422, n5897);
  not g9763 (n_5423, n5898);
  and g9764 (n5899, n_5422, n_5423);
  not g9765 (n_5424, n5895);
  not g9766 (n_5425, n5899);
  and g9767 (n5900, n_5424, n_5425);
  not g9768 (n_5426, n5882);
  not g9769 (n_5427, n5900);
  and g9770 (n5901, n_5426, n_5427);
  not g9771 (n_5428, n5865);
  and g9772 (n5902, n_5428, n5901);
  not g9773 (n_5429, n5901);
  and g9774 (n5903, n5865, n_5429);
  not g9775 (n_5430, n5902);
  not g9776 (n_5431, n5903);
  and g9777 (n5904, n_5430, n_5431);
  not g9778 (n_5433, \A[901] );
  and g9779 (n5905, n_5433, \A[902] );
  not g9780 (n_5435, \A[902] );
  and g9781 (n5906, \A[901] , n_5435);
  not g9782 (n_5437, n5906);
  and g9783 (n5907, \A[903] , n_5437);
  not g9784 (n_5438, n5905);
  and g9785 (n5908, n_5438, n5907);
  and g9786 (n5909, n_5438, n_5437);
  not g9787 (n_5439, \A[903] );
  not g9788 (n_5440, n5909);
  and g9789 (n5910, n_5439, n_5440);
  not g9790 (n_5441, n5908);
  not g9791 (n_5442, n5910);
  and g9792 (n5911, n_5441, n_5442);
  not g9793 (n_5444, \A[904] );
  and g9794 (n5912, n_5444, \A[905] );
  not g9795 (n_5446, \A[905] );
  and g9796 (n5913, \A[904] , n_5446);
  not g9797 (n_5448, n5913);
  and g9798 (n5914, \A[906] , n_5448);
  not g9799 (n_5449, n5912);
  and g9800 (n5915, n_5449, n5914);
  and g9801 (n5916, n_5449, n_5448);
  not g9802 (n_5450, \A[906] );
  not g9803 (n_5451, n5916);
  and g9804 (n5917, n_5450, n_5451);
  not g9805 (n_5452, n5915);
  not g9806 (n_5453, n5917);
  and g9807 (n5918, n_5452, n_5453);
  not g9808 (n_5454, n5911);
  and g9809 (n5919, n_5454, n5918);
  not g9810 (n_5455, n5918);
  and g9811 (n5920, n5911, n_5455);
  not g9812 (n_5456, n5919);
  not g9813 (n_5457, n5920);
  and g9814 (n5921, n_5456, n_5457);
  and g9815 (n5922, \A[904] , \A[905] );
  and g9816 (n5923, \A[906] , n_5451);
  not g9817 (n_5458, n5922);
  not g9818 (n_5459, n5923);
  and g9819 (n5924, n_5458, n_5459);
  and g9820 (n5925, \A[901] , \A[902] );
  and g9821 (n5926, \A[903] , n_5440);
  not g9822 (n_5460, n5925);
  not g9823 (n_5461, n5926);
  and g9824 (n5927, n_5460, n_5461);
  not g9825 (n_5462, n5924);
  and g9826 (n5928, n_5462, n5927);
  not g9827 (n_5463, n5927);
  and g9828 (n5929, n5924, n_5463);
  not g9829 (n_5464, n5928);
  not g9830 (n_5465, n5929);
  and g9831 (n5930, n_5464, n_5465);
  and g9832 (n5931, n_5454, n_5455);
  not g9833 (n_5466, n5930);
  and g9834 (n5932, n_5466, n5931);
  and g9835 (n5933, n_5462, n_5463);
  not g9836 (n_5467, n5932);
  not g9837 (n_5468, n5933);
  and g9838 (n5934, n_5467, n_5468);
  and g9839 (n5935, n_5464, n5931);
  and g9840 (n5936, n_5465, n5935);
  not g9841 (n_5469, n5931);
  and g9842 (n5937, n_5466, n_5469);
  not g9843 (n_5470, n5936);
  not g9844 (n_5471, n5937);
  and g9845 (n5938, n_5470, n_5471);
  not g9846 (n_5472, n5934);
  not g9847 (n_5473, n5938);
  and g9848 (n5939, n_5472, n_5473);
  not g9849 (n_5474, n5921);
  not g9850 (n_5475, n5939);
  and g9851 (n5940, n_5474, n_5475);
  not g9852 (n_5477, \A[895] );
  and g9853 (n5941, n_5477, \A[896] );
  not g9854 (n_5479, \A[896] );
  and g9855 (n5942, \A[895] , n_5479);
  not g9856 (n_5481, n5942);
  and g9857 (n5943, \A[897] , n_5481);
  not g9858 (n_5482, n5941);
  and g9859 (n5944, n_5482, n5943);
  and g9860 (n5945, n_5482, n_5481);
  not g9861 (n_5483, \A[897] );
  not g9862 (n_5484, n5945);
  and g9863 (n5946, n_5483, n_5484);
  not g9864 (n_5485, n5944);
  not g9865 (n_5486, n5946);
  and g9866 (n5947, n_5485, n_5486);
  not g9867 (n_5488, \A[898] );
  and g9868 (n5948, n_5488, \A[899] );
  not g9869 (n_5490, \A[899] );
  and g9870 (n5949, \A[898] , n_5490);
  not g9871 (n_5492, n5949);
  and g9872 (n5950, \A[900] , n_5492);
  not g9873 (n_5493, n5948);
  and g9874 (n5951, n_5493, n5950);
  and g9875 (n5952, n_5493, n_5492);
  not g9876 (n_5494, \A[900] );
  not g9877 (n_5495, n5952);
  and g9878 (n5953, n_5494, n_5495);
  not g9879 (n_5496, n5951);
  not g9880 (n_5497, n5953);
  and g9881 (n5954, n_5496, n_5497);
  not g9882 (n_5498, n5947);
  and g9883 (n5955, n_5498, n5954);
  not g9884 (n_5499, n5954);
  and g9885 (n5956, n5947, n_5499);
  not g9886 (n_5500, n5955);
  not g9887 (n_5501, n5956);
  and g9888 (n5957, n_5500, n_5501);
  and g9889 (n5958, \A[898] , \A[899] );
  and g9890 (n5959, \A[900] , n_5495);
  not g9891 (n_5502, n5958);
  not g9892 (n_5503, n5959);
  and g9893 (n5960, n_5502, n_5503);
  and g9894 (n5961, \A[895] , \A[896] );
  and g9895 (n5962, \A[897] , n_5484);
  not g9896 (n_5504, n5961);
  not g9897 (n_5505, n5962);
  and g9898 (n5963, n_5504, n_5505);
  not g9899 (n_5506, n5960);
  and g9900 (n5964, n_5506, n5963);
  not g9901 (n_5507, n5963);
  and g9902 (n5965, n5960, n_5507);
  not g9903 (n_5508, n5964);
  not g9904 (n_5509, n5965);
  and g9905 (n5966, n_5508, n_5509);
  and g9906 (n5967, n_5498, n_5499);
  not g9907 (n_5510, n5966);
  and g9908 (n5968, n_5510, n5967);
  and g9909 (n5969, n_5506, n_5507);
  not g9910 (n_5511, n5968);
  not g9911 (n_5512, n5969);
  and g9912 (n5970, n_5511, n_5512);
  and g9913 (n5971, n_5508, n5967);
  and g9914 (n5972, n_5509, n5971);
  not g9915 (n_5513, n5967);
  and g9916 (n5973, n_5510, n_5513);
  not g9917 (n_5514, n5972);
  not g9918 (n_5515, n5973);
  and g9919 (n5974, n_5514, n_5515);
  not g9920 (n_5516, n5970);
  not g9921 (n_5517, n5974);
  and g9922 (n5975, n_5516, n_5517);
  not g9923 (n_5518, n5957);
  not g9924 (n_5519, n5975);
  and g9925 (n5976, n_5518, n_5519);
  not g9926 (n_5520, n5940);
  and g9927 (n5977, n_5520, n5976);
  not g9928 (n_5521, n5976);
  and g9929 (n5978, n5940, n_5521);
  not g9930 (n_5522, n5977);
  not g9931 (n_5523, n5978);
  and g9932 (n5979, n_5522, n_5523);
  not g9933 (n_5524, n5904);
  and g9934 (n5980, n_5524, n5979);
  not g9935 (n_5525, n5979);
  and g9936 (n5981, n5904, n_5525);
  not g9937 (n_5526, n5980);
  not g9938 (n_5527, n5981);
  and g9939 (n5982, n_5526, n_5527);
  not g9940 (n_5528, n5829);
  and g9941 (n5983, n_5528, n5982);
  not g9942 (n_5529, n5982);
  and g9943 (n5984, n5829, n_5529);
  not g9944 (n_5530, n5983);
  not g9945 (n_5531, n5984);
  and g9946 (n5985, n_5530, n_5531);
  not g9947 (n_5533, \A[889] );
  and g9948 (n5986, n_5533, \A[890] );
  not g9949 (n_5535, \A[890] );
  and g9950 (n5987, \A[889] , n_5535);
  not g9951 (n_5537, n5987);
  and g9952 (n5988, \A[891] , n_5537);
  not g9953 (n_5538, n5986);
  and g9954 (n5989, n_5538, n5988);
  and g9955 (n5990, n_5538, n_5537);
  not g9956 (n_5539, \A[891] );
  not g9957 (n_5540, n5990);
  and g9958 (n5991, n_5539, n_5540);
  not g9959 (n_5541, n5989);
  not g9960 (n_5542, n5991);
  and g9961 (n5992, n_5541, n_5542);
  not g9962 (n_5544, \A[892] );
  and g9963 (n5993, n_5544, \A[893] );
  not g9964 (n_5546, \A[893] );
  and g9965 (n5994, \A[892] , n_5546);
  not g9966 (n_5548, n5994);
  and g9967 (n5995, \A[894] , n_5548);
  not g9968 (n_5549, n5993);
  and g9969 (n5996, n_5549, n5995);
  and g9970 (n5997, n_5549, n_5548);
  not g9971 (n_5550, \A[894] );
  not g9972 (n_5551, n5997);
  and g9973 (n5998, n_5550, n_5551);
  not g9974 (n_5552, n5996);
  not g9975 (n_5553, n5998);
  and g9976 (n5999, n_5552, n_5553);
  not g9977 (n_5554, n5992);
  and g9978 (n6000, n_5554, n5999);
  not g9979 (n_5555, n5999);
  and g9980 (n6001, n5992, n_5555);
  not g9981 (n_5556, n6000);
  not g9982 (n_5557, n6001);
  and g9983 (n6002, n_5556, n_5557);
  and g9984 (n6003, \A[892] , \A[893] );
  and g9985 (n6004, \A[894] , n_5551);
  not g9986 (n_5558, n6003);
  not g9987 (n_5559, n6004);
  and g9988 (n6005, n_5558, n_5559);
  and g9989 (n6006, \A[889] , \A[890] );
  and g9990 (n6007, \A[891] , n_5540);
  not g9991 (n_5560, n6006);
  not g9992 (n_5561, n6007);
  and g9993 (n6008, n_5560, n_5561);
  not g9994 (n_5562, n6005);
  and g9995 (n6009, n_5562, n6008);
  not g9996 (n_5563, n6008);
  and g9997 (n6010, n6005, n_5563);
  not g9998 (n_5564, n6009);
  not g9999 (n_5565, n6010);
  and g10000 (n6011, n_5564, n_5565);
  and g10001 (n6012, n_5554, n_5555);
  not g10002 (n_5566, n6011);
  and g10003 (n6013, n_5566, n6012);
  and g10004 (n6014, n_5562, n_5563);
  not g10005 (n_5567, n6013);
  not g10006 (n_5568, n6014);
  and g10007 (n6015, n_5567, n_5568);
  and g10008 (n6016, n_5564, n6012);
  and g10009 (n6017, n_5565, n6016);
  not g10010 (n_5569, n6012);
  and g10011 (n6018, n_5566, n_5569);
  not g10012 (n_5570, n6017);
  not g10013 (n_5571, n6018);
  and g10014 (n6019, n_5570, n_5571);
  not g10015 (n_5572, n6015);
  not g10016 (n_5573, n6019);
  and g10017 (n6020, n_5572, n_5573);
  not g10018 (n_5574, n6002);
  not g10019 (n_5575, n6020);
  and g10020 (n6021, n_5574, n_5575);
  not g10021 (n_5577, \A[883] );
  and g10022 (n6022, n_5577, \A[884] );
  not g10023 (n_5579, \A[884] );
  and g10024 (n6023, \A[883] , n_5579);
  not g10025 (n_5581, n6023);
  and g10026 (n6024, \A[885] , n_5581);
  not g10027 (n_5582, n6022);
  and g10028 (n6025, n_5582, n6024);
  and g10029 (n6026, n_5582, n_5581);
  not g10030 (n_5583, \A[885] );
  not g10031 (n_5584, n6026);
  and g10032 (n6027, n_5583, n_5584);
  not g10033 (n_5585, n6025);
  not g10034 (n_5586, n6027);
  and g10035 (n6028, n_5585, n_5586);
  not g10036 (n_5588, \A[886] );
  and g10037 (n6029, n_5588, \A[887] );
  not g10038 (n_5590, \A[887] );
  and g10039 (n6030, \A[886] , n_5590);
  not g10040 (n_5592, n6030);
  and g10041 (n6031, \A[888] , n_5592);
  not g10042 (n_5593, n6029);
  and g10043 (n6032, n_5593, n6031);
  and g10044 (n6033, n_5593, n_5592);
  not g10045 (n_5594, \A[888] );
  not g10046 (n_5595, n6033);
  and g10047 (n6034, n_5594, n_5595);
  not g10048 (n_5596, n6032);
  not g10049 (n_5597, n6034);
  and g10050 (n6035, n_5596, n_5597);
  not g10051 (n_5598, n6028);
  and g10052 (n6036, n_5598, n6035);
  not g10053 (n_5599, n6035);
  and g10054 (n6037, n6028, n_5599);
  not g10055 (n_5600, n6036);
  not g10056 (n_5601, n6037);
  and g10057 (n6038, n_5600, n_5601);
  and g10058 (n6039, \A[886] , \A[887] );
  and g10059 (n6040, \A[888] , n_5595);
  not g10060 (n_5602, n6039);
  not g10061 (n_5603, n6040);
  and g10062 (n6041, n_5602, n_5603);
  and g10063 (n6042, \A[883] , \A[884] );
  and g10064 (n6043, \A[885] , n_5584);
  not g10065 (n_5604, n6042);
  not g10066 (n_5605, n6043);
  and g10067 (n6044, n_5604, n_5605);
  not g10068 (n_5606, n6041);
  and g10069 (n6045, n_5606, n6044);
  not g10070 (n_5607, n6044);
  and g10071 (n6046, n6041, n_5607);
  not g10072 (n_5608, n6045);
  not g10073 (n_5609, n6046);
  and g10074 (n6047, n_5608, n_5609);
  and g10075 (n6048, n_5598, n_5599);
  not g10076 (n_5610, n6047);
  and g10077 (n6049, n_5610, n6048);
  and g10078 (n6050, n_5606, n_5607);
  not g10079 (n_5611, n6049);
  not g10080 (n_5612, n6050);
  and g10081 (n6051, n_5611, n_5612);
  and g10082 (n6052, n_5608, n6048);
  and g10083 (n6053, n_5609, n6052);
  not g10084 (n_5613, n6048);
  and g10085 (n6054, n_5610, n_5613);
  not g10086 (n_5614, n6053);
  not g10087 (n_5615, n6054);
  and g10088 (n6055, n_5614, n_5615);
  not g10089 (n_5616, n6051);
  not g10090 (n_5617, n6055);
  and g10091 (n6056, n_5616, n_5617);
  not g10092 (n_5618, n6038);
  not g10093 (n_5619, n6056);
  and g10094 (n6057, n_5618, n_5619);
  not g10095 (n_5620, n6021);
  and g10096 (n6058, n_5620, n6057);
  not g10097 (n_5621, n6057);
  and g10098 (n6059, n6021, n_5621);
  not g10099 (n_5622, n6058);
  not g10100 (n_5623, n6059);
  and g10101 (n6060, n_5622, n_5623);
  not g10102 (n_5625, \A[877] );
  and g10103 (n6061, n_5625, \A[878] );
  not g10104 (n_5627, \A[878] );
  and g10105 (n6062, \A[877] , n_5627);
  not g10106 (n_5629, n6062);
  and g10107 (n6063, \A[879] , n_5629);
  not g10108 (n_5630, n6061);
  and g10109 (n6064, n_5630, n6063);
  and g10110 (n6065, n_5630, n_5629);
  not g10111 (n_5631, \A[879] );
  not g10112 (n_5632, n6065);
  and g10113 (n6066, n_5631, n_5632);
  not g10114 (n_5633, n6064);
  not g10115 (n_5634, n6066);
  and g10116 (n6067, n_5633, n_5634);
  not g10117 (n_5636, \A[880] );
  and g10118 (n6068, n_5636, \A[881] );
  not g10119 (n_5638, \A[881] );
  and g10120 (n6069, \A[880] , n_5638);
  not g10121 (n_5640, n6069);
  and g10122 (n6070, \A[882] , n_5640);
  not g10123 (n_5641, n6068);
  and g10124 (n6071, n_5641, n6070);
  and g10125 (n6072, n_5641, n_5640);
  not g10126 (n_5642, \A[882] );
  not g10127 (n_5643, n6072);
  and g10128 (n6073, n_5642, n_5643);
  not g10129 (n_5644, n6071);
  not g10130 (n_5645, n6073);
  and g10131 (n6074, n_5644, n_5645);
  not g10132 (n_5646, n6067);
  and g10133 (n6075, n_5646, n6074);
  not g10134 (n_5647, n6074);
  and g10135 (n6076, n6067, n_5647);
  not g10136 (n_5648, n6075);
  not g10137 (n_5649, n6076);
  and g10138 (n6077, n_5648, n_5649);
  and g10139 (n6078, \A[880] , \A[881] );
  and g10140 (n6079, \A[882] , n_5643);
  not g10141 (n_5650, n6078);
  not g10142 (n_5651, n6079);
  and g10143 (n6080, n_5650, n_5651);
  and g10144 (n6081, \A[877] , \A[878] );
  and g10145 (n6082, \A[879] , n_5632);
  not g10146 (n_5652, n6081);
  not g10147 (n_5653, n6082);
  and g10148 (n6083, n_5652, n_5653);
  not g10149 (n_5654, n6080);
  and g10150 (n6084, n_5654, n6083);
  not g10151 (n_5655, n6083);
  and g10152 (n6085, n6080, n_5655);
  not g10153 (n_5656, n6084);
  not g10154 (n_5657, n6085);
  and g10155 (n6086, n_5656, n_5657);
  and g10156 (n6087, n_5646, n_5647);
  not g10157 (n_5658, n6086);
  and g10158 (n6088, n_5658, n6087);
  and g10159 (n6089, n_5654, n_5655);
  not g10160 (n_5659, n6088);
  not g10161 (n_5660, n6089);
  and g10162 (n6090, n_5659, n_5660);
  and g10163 (n6091, n_5656, n6087);
  and g10164 (n6092, n_5657, n6091);
  not g10165 (n_5661, n6087);
  and g10166 (n6093, n_5658, n_5661);
  not g10167 (n_5662, n6092);
  not g10168 (n_5663, n6093);
  and g10169 (n6094, n_5662, n_5663);
  not g10170 (n_5664, n6090);
  not g10171 (n_5665, n6094);
  and g10172 (n6095, n_5664, n_5665);
  not g10173 (n_5666, n6077);
  not g10174 (n_5667, n6095);
  and g10175 (n6096, n_5666, n_5667);
  not g10176 (n_5669, \A[871] );
  and g10177 (n6097, n_5669, \A[872] );
  not g10178 (n_5671, \A[872] );
  and g10179 (n6098, \A[871] , n_5671);
  not g10180 (n_5673, n6098);
  and g10181 (n6099, \A[873] , n_5673);
  not g10182 (n_5674, n6097);
  and g10183 (n6100, n_5674, n6099);
  and g10184 (n6101, n_5674, n_5673);
  not g10185 (n_5675, \A[873] );
  not g10186 (n_5676, n6101);
  and g10187 (n6102, n_5675, n_5676);
  not g10188 (n_5677, n6100);
  not g10189 (n_5678, n6102);
  and g10190 (n6103, n_5677, n_5678);
  not g10191 (n_5680, \A[874] );
  and g10192 (n6104, n_5680, \A[875] );
  not g10193 (n_5682, \A[875] );
  and g10194 (n6105, \A[874] , n_5682);
  not g10195 (n_5684, n6105);
  and g10196 (n6106, \A[876] , n_5684);
  not g10197 (n_5685, n6104);
  and g10198 (n6107, n_5685, n6106);
  and g10199 (n6108, n_5685, n_5684);
  not g10200 (n_5686, \A[876] );
  not g10201 (n_5687, n6108);
  and g10202 (n6109, n_5686, n_5687);
  not g10203 (n_5688, n6107);
  not g10204 (n_5689, n6109);
  and g10205 (n6110, n_5688, n_5689);
  not g10206 (n_5690, n6103);
  and g10207 (n6111, n_5690, n6110);
  not g10208 (n_5691, n6110);
  and g10209 (n6112, n6103, n_5691);
  not g10210 (n_5692, n6111);
  not g10211 (n_5693, n6112);
  and g10212 (n6113, n_5692, n_5693);
  and g10213 (n6114, \A[874] , \A[875] );
  and g10214 (n6115, \A[876] , n_5687);
  not g10215 (n_5694, n6114);
  not g10216 (n_5695, n6115);
  and g10217 (n6116, n_5694, n_5695);
  and g10218 (n6117, \A[871] , \A[872] );
  and g10219 (n6118, \A[873] , n_5676);
  not g10220 (n_5696, n6117);
  not g10221 (n_5697, n6118);
  and g10222 (n6119, n_5696, n_5697);
  not g10223 (n_5698, n6116);
  and g10224 (n6120, n_5698, n6119);
  not g10225 (n_5699, n6119);
  and g10226 (n6121, n6116, n_5699);
  not g10227 (n_5700, n6120);
  not g10228 (n_5701, n6121);
  and g10229 (n6122, n_5700, n_5701);
  and g10230 (n6123, n_5690, n_5691);
  not g10231 (n_5702, n6122);
  and g10232 (n6124, n_5702, n6123);
  and g10233 (n6125, n_5698, n_5699);
  not g10234 (n_5703, n6124);
  not g10235 (n_5704, n6125);
  and g10236 (n6126, n_5703, n_5704);
  and g10237 (n6127, n_5700, n6123);
  and g10238 (n6128, n_5701, n6127);
  not g10239 (n_5705, n6123);
  and g10240 (n6129, n_5702, n_5705);
  not g10241 (n_5706, n6128);
  not g10242 (n_5707, n6129);
  and g10243 (n6130, n_5706, n_5707);
  not g10244 (n_5708, n6126);
  not g10245 (n_5709, n6130);
  and g10246 (n6131, n_5708, n_5709);
  not g10247 (n_5710, n6113);
  not g10248 (n_5711, n6131);
  and g10249 (n6132, n_5710, n_5711);
  not g10250 (n_5712, n6096);
  and g10251 (n6133, n_5712, n6132);
  not g10252 (n_5713, n6132);
  and g10253 (n6134, n6096, n_5713);
  not g10254 (n_5714, n6133);
  not g10255 (n_5715, n6134);
  and g10256 (n6135, n_5714, n_5715);
  not g10257 (n_5716, n6060);
  and g10258 (n6136, n_5716, n6135);
  not g10259 (n_5717, n6135);
  and g10260 (n6137, n6060, n_5717);
  not g10261 (n_5718, n6136);
  not g10262 (n_5719, n6137);
  and g10263 (n6138, n_5718, n_5719);
  not g10264 (n_5721, \A[865] );
  and g10265 (n6139, n_5721, \A[866] );
  not g10266 (n_5723, \A[866] );
  and g10267 (n6140, \A[865] , n_5723);
  not g10268 (n_5725, n6140);
  and g10269 (n6141, \A[867] , n_5725);
  not g10270 (n_5726, n6139);
  and g10271 (n6142, n_5726, n6141);
  and g10272 (n6143, n_5726, n_5725);
  not g10273 (n_5727, \A[867] );
  not g10274 (n_5728, n6143);
  and g10275 (n6144, n_5727, n_5728);
  not g10276 (n_5729, n6142);
  not g10277 (n_5730, n6144);
  and g10278 (n6145, n_5729, n_5730);
  not g10279 (n_5732, \A[868] );
  and g10280 (n6146, n_5732, \A[869] );
  not g10281 (n_5734, \A[869] );
  and g10282 (n6147, \A[868] , n_5734);
  not g10283 (n_5736, n6147);
  and g10284 (n6148, \A[870] , n_5736);
  not g10285 (n_5737, n6146);
  and g10286 (n6149, n_5737, n6148);
  and g10287 (n6150, n_5737, n_5736);
  not g10288 (n_5738, \A[870] );
  not g10289 (n_5739, n6150);
  and g10290 (n6151, n_5738, n_5739);
  not g10291 (n_5740, n6149);
  not g10292 (n_5741, n6151);
  and g10293 (n6152, n_5740, n_5741);
  not g10294 (n_5742, n6145);
  and g10295 (n6153, n_5742, n6152);
  not g10296 (n_5743, n6152);
  and g10297 (n6154, n6145, n_5743);
  not g10298 (n_5744, n6153);
  not g10299 (n_5745, n6154);
  and g10300 (n6155, n_5744, n_5745);
  and g10301 (n6156, \A[868] , \A[869] );
  and g10302 (n6157, \A[870] , n_5739);
  not g10303 (n_5746, n6156);
  not g10304 (n_5747, n6157);
  and g10305 (n6158, n_5746, n_5747);
  and g10306 (n6159, \A[865] , \A[866] );
  and g10307 (n6160, \A[867] , n_5728);
  not g10308 (n_5748, n6159);
  not g10309 (n_5749, n6160);
  and g10310 (n6161, n_5748, n_5749);
  not g10311 (n_5750, n6158);
  and g10312 (n6162, n_5750, n6161);
  not g10313 (n_5751, n6161);
  and g10314 (n6163, n6158, n_5751);
  not g10315 (n_5752, n6162);
  not g10316 (n_5753, n6163);
  and g10317 (n6164, n_5752, n_5753);
  and g10318 (n6165, n_5742, n_5743);
  not g10319 (n_5754, n6164);
  and g10320 (n6166, n_5754, n6165);
  and g10321 (n6167, n_5750, n_5751);
  not g10322 (n_5755, n6166);
  not g10323 (n_5756, n6167);
  and g10324 (n6168, n_5755, n_5756);
  and g10325 (n6169, n_5752, n6165);
  and g10326 (n6170, n_5753, n6169);
  not g10327 (n_5757, n6165);
  and g10328 (n6171, n_5754, n_5757);
  not g10329 (n_5758, n6170);
  not g10330 (n_5759, n6171);
  and g10331 (n6172, n_5758, n_5759);
  not g10332 (n_5760, n6168);
  not g10333 (n_5761, n6172);
  and g10334 (n6173, n_5760, n_5761);
  not g10335 (n_5762, n6155);
  not g10336 (n_5763, n6173);
  and g10337 (n6174, n_5762, n_5763);
  not g10338 (n_5765, \A[859] );
  and g10339 (n6175, n_5765, \A[860] );
  not g10340 (n_5767, \A[860] );
  and g10341 (n6176, \A[859] , n_5767);
  not g10342 (n_5769, n6176);
  and g10343 (n6177, \A[861] , n_5769);
  not g10344 (n_5770, n6175);
  and g10345 (n6178, n_5770, n6177);
  and g10346 (n6179, n_5770, n_5769);
  not g10347 (n_5771, \A[861] );
  not g10348 (n_5772, n6179);
  and g10349 (n6180, n_5771, n_5772);
  not g10350 (n_5773, n6178);
  not g10351 (n_5774, n6180);
  and g10352 (n6181, n_5773, n_5774);
  not g10353 (n_5776, \A[862] );
  and g10354 (n6182, n_5776, \A[863] );
  not g10355 (n_5778, \A[863] );
  and g10356 (n6183, \A[862] , n_5778);
  not g10357 (n_5780, n6183);
  and g10358 (n6184, \A[864] , n_5780);
  not g10359 (n_5781, n6182);
  and g10360 (n6185, n_5781, n6184);
  and g10361 (n6186, n_5781, n_5780);
  not g10362 (n_5782, \A[864] );
  not g10363 (n_5783, n6186);
  and g10364 (n6187, n_5782, n_5783);
  not g10365 (n_5784, n6185);
  not g10366 (n_5785, n6187);
  and g10367 (n6188, n_5784, n_5785);
  not g10368 (n_5786, n6181);
  and g10369 (n6189, n_5786, n6188);
  not g10370 (n_5787, n6188);
  and g10371 (n6190, n6181, n_5787);
  not g10372 (n_5788, n6189);
  not g10373 (n_5789, n6190);
  and g10374 (n6191, n_5788, n_5789);
  and g10375 (n6192, \A[862] , \A[863] );
  and g10376 (n6193, \A[864] , n_5783);
  not g10377 (n_5790, n6192);
  not g10378 (n_5791, n6193);
  and g10379 (n6194, n_5790, n_5791);
  and g10380 (n6195, \A[859] , \A[860] );
  and g10381 (n6196, \A[861] , n_5772);
  not g10382 (n_5792, n6195);
  not g10383 (n_5793, n6196);
  and g10384 (n6197, n_5792, n_5793);
  not g10385 (n_5794, n6194);
  and g10386 (n6198, n_5794, n6197);
  not g10387 (n_5795, n6197);
  and g10388 (n6199, n6194, n_5795);
  not g10389 (n_5796, n6198);
  not g10390 (n_5797, n6199);
  and g10391 (n6200, n_5796, n_5797);
  and g10392 (n6201, n_5786, n_5787);
  not g10393 (n_5798, n6200);
  and g10394 (n6202, n_5798, n6201);
  and g10395 (n6203, n_5794, n_5795);
  not g10396 (n_5799, n6202);
  not g10397 (n_5800, n6203);
  and g10398 (n6204, n_5799, n_5800);
  and g10399 (n6205, n_5796, n6201);
  and g10400 (n6206, n_5797, n6205);
  not g10401 (n_5801, n6201);
  and g10402 (n6207, n_5798, n_5801);
  not g10403 (n_5802, n6206);
  not g10404 (n_5803, n6207);
  and g10405 (n6208, n_5802, n_5803);
  not g10406 (n_5804, n6204);
  not g10407 (n_5805, n6208);
  and g10408 (n6209, n_5804, n_5805);
  not g10409 (n_5806, n6191);
  not g10410 (n_5807, n6209);
  and g10411 (n6210, n_5806, n_5807);
  not g10412 (n_5808, n6174);
  and g10413 (n6211, n_5808, n6210);
  not g10414 (n_5809, n6210);
  and g10415 (n6212, n6174, n_5809);
  not g10416 (n_5810, n6211);
  not g10417 (n_5811, n6212);
  and g10418 (n6213, n_5810, n_5811);
  not g10419 (n_5813, \A[853] );
  and g10420 (n6214, n_5813, \A[854] );
  not g10421 (n_5815, \A[854] );
  and g10422 (n6215, \A[853] , n_5815);
  not g10423 (n_5817, n6215);
  and g10424 (n6216, \A[855] , n_5817);
  not g10425 (n_5818, n6214);
  and g10426 (n6217, n_5818, n6216);
  and g10427 (n6218, n_5818, n_5817);
  not g10428 (n_5819, \A[855] );
  not g10429 (n_5820, n6218);
  and g10430 (n6219, n_5819, n_5820);
  not g10431 (n_5821, n6217);
  not g10432 (n_5822, n6219);
  and g10433 (n6220, n_5821, n_5822);
  not g10434 (n_5824, \A[856] );
  and g10435 (n6221, n_5824, \A[857] );
  not g10436 (n_5826, \A[857] );
  and g10437 (n6222, \A[856] , n_5826);
  not g10438 (n_5828, n6222);
  and g10439 (n6223, \A[858] , n_5828);
  not g10440 (n_5829, n6221);
  and g10441 (n6224, n_5829, n6223);
  and g10442 (n6225, n_5829, n_5828);
  not g10443 (n_5830, \A[858] );
  not g10444 (n_5831, n6225);
  and g10445 (n6226, n_5830, n_5831);
  not g10446 (n_5832, n6224);
  not g10447 (n_5833, n6226);
  and g10448 (n6227, n_5832, n_5833);
  not g10449 (n_5834, n6220);
  and g10450 (n6228, n_5834, n6227);
  not g10451 (n_5835, n6227);
  and g10452 (n6229, n6220, n_5835);
  not g10453 (n_5836, n6228);
  not g10454 (n_5837, n6229);
  and g10455 (n6230, n_5836, n_5837);
  and g10456 (n6231, \A[856] , \A[857] );
  and g10457 (n6232, \A[858] , n_5831);
  not g10458 (n_5838, n6231);
  not g10459 (n_5839, n6232);
  and g10460 (n6233, n_5838, n_5839);
  and g10461 (n6234, \A[853] , \A[854] );
  and g10462 (n6235, \A[855] , n_5820);
  not g10463 (n_5840, n6234);
  not g10464 (n_5841, n6235);
  and g10465 (n6236, n_5840, n_5841);
  not g10466 (n_5842, n6233);
  and g10467 (n6237, n_5842, n6236);
  not g10468 (n_5843, n6236);
  and g10469 (n6238, n6233, n_5843);
  not g10470 (n_5844, n6237);
  not g10471 (n_5845, n6238);
  and g10472 (n6239, n_5844, n_5845);
  and g10473 (n6240, n_5834, n_5835);
  not g10474 (n_5846, n6239);
  and g10475 (n6241, n_5846, n6240);
  and g10476 (n6242, n_5842, n_5843);
  not g10477 (n_5847, n6241);
  not g10478 (n_5848, n6242);
  and g10479 (n6243, n_5847, n_5848);
  and g10480 (n6244, n_5844, n6240);
  and g10481 (n6245, n_5845, n6244);
  not g10482 (n_5849, n6240);
  and g10483 (n6246, n_5846, n_5849);
  not g10484 (n_5850, n6245);
  not g10485 (n_5851, n6246);
  and g10486 (n6247, n_5850, n_5851);
  not g10487 (n_5852, n6243);
  not g10488 (n_5853, n6247);
  and g10489 (n6248, n_5852, n_5853);
  not g10490 (n_5854, n6230);
  not g10491 (n_5855, n6248);
  and g10492 (n6249, n_5854, n_5855);
  not g10493 (n_5857, \A[847] );
  and g10494 (n6250, n_5857, \A[848] );
  not g10495 (n_5859, \A[848] );
  and g10496 (n6251, \A[847] , n_5859);
  not g10497 (n_5861, n6251);
  and g10498 (n6252, \A[849] , n_5861);
  not g10499 (n_5862, n6250);
  and g10500 (n6253, n_5862, n6252);
  and g10501 (n6254, n_5862, n_5861);
  not g10502 (n_5863, \A[849] );
  not g10503 (n_5864, n6254);
  and g10504 (n6255, n_5863, n_5864);
  not g10505 (n_5865, n6253);
  not g10506 (n_5866, n6255);
  and g10507 (n6256, n_5865, n_5866);
  not g10508 (n_5868, \A[850] );
  and g10509 (n6257, n_5868, \A[851] );
  not g10510 (n_5870, \A[851] );
  and g10511 (n6258, \A[850] , n_5870);
  not g10512 (n_5872, n6258);
  and g10513 (n6259, \A[852] , n_5872);
  not g10514 (n_5873, n6257);
  and g10515 (n6260, n_5873, n6259);
  and g10516 (n6261, n_5873, n_5872);
  not g10517 (n_5874, \A[852] );
  not g10518 (n_5875, n6261);
  and g10519 (n6262, n_5874, n_5875);
  not g10520 (n_5876, n6260);
  not g10521 (n_5877, n6262);
  and g10522 (n6263, n_5876, n_5877);
  not g10523 (n_5878, n6256);
  and g10524 (n6264, n_5878, n6263);
  not g10525 (n_5879, n6263);
  and g10526 (n6265, n6256, n_5879);
  not g10527 (n_5880, n6264);
  not g10528 (n_5881, n6265);
  and g10529 (n6266, n_5880, n_5881);
  and g10530 (n6267, \A[850] , \A[851] );
  and g10531 (n6268, \A[852] , n_5875);
  not g10532 (n_5882, n6267);
  not g10533 (n_5883, n6268);
  and g10534 (n6269, n_5882, n_5883);
  and g10535 (n6270, \A[847] , \A[848] );
  and g10536 (n6271, \A[849] , n_5864);
  not g10537 (n_5884, n6270);
  not g10538 (n_5885, n6271);
  and g10539 (n6272, n_5884, n_5885);
  not g10540 (n_5886, n6269);
  and g10541 (n6273, n_5886, n6272);
  not g10542 (n_5887, n6272);
  and g10543 (n6274, n6269, n_5887);
  not g10544 (n_5888, n6273);
  not g10545 (n_5889, n6274);
  and g10546 (n6275, n_5888, n_5889);
  and g10547 (n6276, n_5878, n_5879);
  not g10548 (n_5890, n6275);
  and g10549 (n6277, n_5890, n6276);
  and g10550 (n6278, n_5886, n_5887);
  not g10551 (n_5891, n6277);
  not g10552 (n_5892, n6278);
  and g10553 (n6279, n_5891, n_5892);
  and g10554 (n6280, n_5888, n6276);
  and g10555 (n6281, n_5889, n6280);
  not g10556 (n_5893, n6276);
  and g10557 (n6282, n_5890, n_5893);
  not g10558 (n_5894, n6281);
  not g10559 (n_5895, n6282);
  and g10560 (n6283, n_5894, n_5895);
  not g10561 (n_5896, n6279);
  not g10562 (n_5897, n6283);
  and g10563 (n6284, n_5896, n_5897);
  not g10564 (n_5898, n6266);
  not g10565 (n_5899, n6284);
  and g10566 (n6285, n_5898, n_5899);
  not g10567 (n_5900, n6249);
  and g10568 (n6286, n_5900, n6285);
  not g10569 (n_5901, n6285);
  and g10570 (n6287, n6249, n_5901);
  not g10571 (n_5902, n6286);
  not g10572 (n_5903, n6287);
  and g10573 (n6288, n_5902, n_5903);
  not g10574 (n_5904, n6213);
  and g10575 (n6289, n_5904, n6288);
  not g10576 (n_5905, n6288);
  and g10577 (n6290, n6213, n_5905);
  not g10578 (n_5906, n6289);
  not g10579 (n_5907, n6290);
  and g10580 (n6291, n_5906, n_5907);
  not g10581 (n_5908, n6138);
  and g10582 (n6292, n_5908, n6291);
  not g10583 (n_5909, n6291);
  and g10584 (n6293, n6138, n_5909);
  not g10585 (n_5910, n6292);
  not g10586 (n_5911, n6293);
  and g10587 (n6294, n_5910, n_5911);
  not g10588 (n_5912, n5985);
  and g10589 (n6295, n_5912, n6294);
  not g10590 (n_5913, n6294);
  and g10591 (n6296, n5985, n_5913);
  not g10592 (n_5914, n6295);
  not g10593 (n_5915, n6296);
  and g10594 (n6297, n_5914, n_5915);
  not g10595 (n_5916, n5676);
  not g10596 (n_5917, n6297);
  and g10597 (n6298, n_5916, n_5917);
  not g10598 (n_5918, n5672);
  and g10599 (n6299, n_5918, n6298);
  not g10600 (n_5919, n5667);
  and g10601 (n6300, n_5919, n6299);
  and g10602 (n6301, n_5919, n_5918);
  not g10603 (n_5920, n6298);
  not g10604 (n_5921, n6301);
  and g10605 (n6302, n_5920, n_5921);
  not g10606 (n_5922, n6300);
  not g10607 (n_5923, n6302);
  and g10608 (n6303, n_5922, n_5923);
  and g10609 (n6304, n_5426, n_5424);
  not g10610 (n_5924, n6304);
  and g10611 (n6305, n_5425, n_5924);
  and g10612 (n6306, n_5382, n_5426);
  and g10613 (n6307, n_5383, n6306);
  and g10614 (n6308, n_5427, n6307);
  and g10615 (n6309, n_5382, n_5380);
  not g10616 (n_5925, n6309);
  and g10617 (n6310, n_5381, n_5925);
  not g10618 (n_5926, n6308);
  not g10619 (n_5927, n6310);
  and g10620 (n6311, n_5926, n_5927);
  not g10625 (n_5928, n6311);
  not g10626 (n_5929, n6315);
  and g10627 (n6316, n_5928, n_5929);
  not g10628 (n_5930, n6316);
  and g10629 (n6317, n6305, n_5930);
  and g10630 (n6318, n_5926, n6310);
  and g10631 (n6319, n6308, n_5927);
  not g10632 (n_5931, n6318);
  not g10633 (n_5932, n6319);
  and g10634 (n6320, n_5931, n_5932);
  not g10635 (n_5933, n6305);
  not g10636 (n_5934, n6320);
  and g10637 (n6321, n_5933, n_5934);
  and g10638 (n6322, n_5524, n_5525);
  not g10639 (n_5935, n6321);
  and g10640 (n6323, n_5935, n6322);
  not g10641 (n_5936, n6317);
  and g10642 (n6324, n_5936, n6323);
  and g10643 (n6325, n_5936, n_5935);
  not g10644 (n_5937, n6322);
  not g10645 (n_5938, n6325);
  and g10646 (n6326, n_5937, n_5938);
  not g10647 (n_5939, n6324);
  not g10648 (n_5940, n6326);
  and g10649 (n6327, n_5939, n_5940);
  and g10650 (n6328, n_5518, n_5516);
  not g10651 (n_5941, n6328);
  and g10652 (n6329, n_5517, n_5941);
  and g10653 (n6330, n_5474, n_5518);
  and g10654 (n6331, n_5475, n6330);
  and g10655 (n6332, n_5519, n6331);
  and g10656 (n6333, n_5474, n_5472);
  not g10657 (n_5942, n6333);
  and g10658 (n6334, n_5473, n_5942);
  not g10659 (n_5943, n6332);
  and g10660 (n6335, n_5943, n6334);
  not g10661 (n_5944, n6334);
  and g10662 (n6336, n6332, n_5944);
  not g10663 (n_5945, n6335);
  not g10664 (n_5946, n6336);
  and g10665 (n6337, n_5945, n_5946);
  not g10666 (n_5947, n6329);
  not g10667 (n_5948, n6337);
  and g10668 (n6338, n_5947, n_5948);
  and g10669 (n6339, n_5943, n_5944);
  not g10674 (n_5949, n6339);
  not g10675 (n_5950, n6343);
  and g10676 (n6344, n_5949, n_5950);
  not g10677 (n_5951, n6344);
  and g10678 (n6345, n6329, n_5951);
  not g10679 (n_5952, n6338);
  not g10680 (n_5953, n6345);
  and g10681 (n6346, n_5952, n_5953);
  not g10682 (n_5954, n6327);
  and g10683 (n6347, n_5954, n6346);
  and g10684 (n6348, n_5935, n_5937);
  and g10685 (n6349, n_5936, n6348);
  and g10686 (n6350, n6322, n_5938);
  not g10687 (n_5955, n6349);
  not g10688 (n_5956, n6350);
  and g10689 (n6351, n_5955, n_5956);
  not g10690 (n_5957, n6346);
  not g10691 (n_5958, n6351);
  and g10692 (n6352, n_5957, n_5958);
  not g10693 (n_5959, n6347);
  not g10694 (n_5960, n6352);
  and g10695 (n6353, n_5959, n_5960);
  and g10696 (n6354, n_5330, n_5328);
  not g10697 (n_5961, n6354);
  and g10698 (n6355, n_5329, n_5961);
  and g10699 (n6356, n_5286, n_5330);
  and g10700 (n6357, n_5287, n6356);
  and g10701 (n6358, n_5331, n6357);
  and g10702 (n6359, n_5286, n_5284);
  not g10703 (n_5962, n6359);
  and g10704 (n6360, n_5285, n_5962);
  not g10705 (n_5963, n6358);
  and g10706 (n6361, n_5963, n6360);
  not g10707 (n_5964, n6360);
  and g10708 (n6362, n6358, n_5964);
  not g10709 (n_5965, n6361);
  not g10710 (n_5966, n6362);
  and g10711 (n6363, n_5965, n_5966);
  not g10712 (n_5967, n6355);
  not g10713 (n_5968, n6363);
  and g10714 (n6364, n_5967, n_5968);
  and g10715 (n6365, n_5963, n_5964);
  not g10720 (n_5969, n6365);
  not g10721 (n_5970, n6369);
  and g10722 (n6370, n_5969, n_5970);
  not g10723 (n_5971, n6370);
  and g10724 (n6371, n6355, n_5971);
  not g10725 (n_5972, n6364);
  not g10726 (n_5973, n6371);
  and g10727 (n6372, n_5972, n_5973);
  and g10728 (n6373, n_5238, n_5236);
  not g10729 (n_5974, n6373);
  and g10730 (n6374, n_5237, n_5974);
  and g10731 (n6375, n_5194, n_5238);
  and g10732 (n6376, n_5195, n6375);
  and g10733 (n6377, n_5239, n6376);
  and g10734 (n6378, n_5194, n_5192);
  not g10735 (n_5975, n6378);
  and g10736 (n6379, n_5193, n_5975);
  not g10737 (n_5976, n6377);
  not g10738 (n_5977, n6379);
  and g10739 (n6380, n_5976, n_5977);
  not g10744 (n_5978, n6380);
  not g10745 (n_5979, n6384);
  and g10746 (n6385, n_5978, n_5979);
  not g10747 (n_5980, n6385);
  and g10748 (n6386, n6374, n_5980);
  and g10749 (n6387, n_5976, n6379);
  and g10750 (n6388, n6377, n_5977);
  not g10751 (n_5981, n6387);
  not g10752 (n_5982, n6388);
  and g10753 (n6389, n_5981, n_5982);
  not g10754 (n_5983, n6374);
  not g10755 (n_5984, n6389);
  and g10756 (n6390, n_5983, n_5984);
  and g10757 (n6391, n_5336, n_5337);
  not g10758 (n_5985, n6390);
  not g10759 (n_5986, n6391);
  and g10760 (n6392, n_5985, n_5986);
  not g10761 (n_5987, n6386);
  and g10762 (n6393, n_5987, n6392);
  and g10763 (n6394, n_5987, n_5985);
  not g10764 (n_5988, n6394);
  and g10765 (n6395, n6391, n_5988);
  not g10766 (n_5989, n6393);
  not g10767 (n_5990, n6395);
  and g10768 (n6396, n_5989, n_5990);
  not g10769 (n_5991, n6372);
  not g10770 (n_5992, n6396);
  and g10771 (n6397, n_5991, n_5992);
  and g10772 (n6398, n_5985, n6391);
  and g10773 (n6399, n_5987, n6398);
  and g10774 (n6400, n_5986, n_5988);
  not g10775 (n_5993, n6399);
  not g10776 (n_5994, n6400);
  and g10777 (n6401, n_5993, n_5994);
  not g10778 (n_5995, n6401);
  and g10779 (n6402, n6372, n_5995);
  and g10780 (n6403, n_5528, n_5529);
  not g10781 (n_5996, n6402);
  not g10782 (n_5997, n6403);
  and g10783 (n6404, n_5996, n_5997);
  not g10784 (n_5998, n6397);
  and g10785 (n6405, n_5998, n6404);
  and g10786 (n6406, n_5998, n_5996);
  not g10787 (n_5999, n6406);
  and g10788 (n6407, n6403, n_5999);
  not g10789 (n_6000, n6405);
  not g10790 (n_6001, n6407);
  and g10791 (n6408, n_6000, n_6001);
  not g10792 (n_6002, n6353);
  not g10793 (n_6003, n6408);
  and g10794 (n6409, n_6002, n_6003);
  and g10795 (n6410, n_5996, n6403);
  and g10796 (n6411, n_5998, n6410);
  and g10797 (n6412, n_5997, n_5999);
  not g10798 (n_6004, n6411);
  not g10799 (n_6005, n6412);
  and g10800 (n6413, n_6004, n_6005);
  not g10801 (n_6006, n6413);
  and g10802 (n6414, n6353, n_6006);
  and g10803 (n6415, n_5912, n_5913);
  not g10804 (n_6007, n6414);
  and g10805 (n6416, n_6007, n6415);
  not g10806 (n_6008, n6409);
  and g10807 (n6417, n_6008, n6416);
  and g10808 (n6418, n_6008, n_6007);
  not g10809 (n_6009, n6415);
  not g10810 (n_6010, n6418);
  and g10811 (n6419, n_6009, n_6010);
  not g10812 (n_6011, n6417);
  not g10813 (n_6012, n6419);
  and g10814 (n6420, n_6011, n_6012);
  and g10815 (n6421, n_5710, n_5708);
  not g10816 (n_6013, n6421);
  and g10817 (n6422, n_5709, n_6013);
  and g10818 (n6423, n_5666, n_5710);
  and g10819 (n6424, n_5667, n6423);
  and g10820 (n6425, n_5711, n6424);
  and g10821 (n6426, n_5666, n_5664);
  not g10822 (n_6014, n6426);
  and g10823 (n6427, n_5665, n_6014);
  not g10824 (n_6015, n6425);
  and g10825 (n6428, n_6015, n6427);
  not g10826 (n_6016, n6427);
  and g10827 (n6429, n6425, n_6016);
  not g10828 (n_6017, n6428);
  not g10829 (n_6018, n6429);
  and g10830 (n6430, n_6017, n_6018);
  not g10831 (n_6019, n6422);
  not g10832 (n_6020, n6430);
  and g10833 (n6431, n_6019, n_6020);
  and g10834 (n6432, n_6015, n_6016);
  not g10839 (n_6021, n6432);
  not g10840 (n_6022, n6436);
  and g10841 (n6437, n_6021, n_6022);
  not g10842 (n_6023, n6437);
  and g10843 (n6438, n6422, n_6023);
  not g10844 (n_6024, n6431);
  not g10845 (n_6025, n6438);
  and g10846 (n6439, n_6024, n_6025);
  and g10847 (n6440, n_5618, n_5616);
  not g10848 (n_6026, n6440);
  and g10849 (n6441, n_5617, n_6026);
  and g10850 (n6442, n_5574, n_5618);
  and g10851 (n6443, n_5575, n6442);
  and g10852 (n6444, n_5619, n6443);
  and g10853 (n6445, n_5574, n_5572);
  not g10854 (n_6027, n6445);
  and g10855 (n6446, n_5573, n_6027);
  not g10856 (n_6028, n6444);
  not g10857 (n_6029, n6446);
  and g10858 (n6447, n_6028, n_6029);
  not g10863 (n_6030, n6447);
  not g10864 (n_6031, n6451);
  and g10865 (n6452, n_6030, n_6031);
  not g10866 (n_6032, n6452);
  and g10867 (n6453, n6441, n_6032);
  and g10868 (n6454, n_6028, n6446);
  and g10869 (n6455, n6444, n_6029);
  not g10870 (n_6033, n6454);
  not g10871 (n_6034, n6455);
  and g10872 (n6456, n_6033, n_6034);
  not g10873 (n_6035, n6441);
  not g10874 (n_6036, n6456);
  and g10875 (n6457, n_6035, n_6036);
  and g10876 (n6458, n_5716, n_5717);
  not g10877 (n_6037, n6457);
  not g10878 (n_6038, n6458);
  and g10879 (n6459, n_6037, n_6038);
  not g10880 (n_6039, n6453);
  and g10881 (n6460, n_6039, n6459);
  and g10882 (n6461, n_6039, n_6037);
  not g10883 (n_6040, n6461);
  and g10884 (n6462, n6458, n_6040);
  not g10885 (n_6041, n6460);
  not g10886 (n_6042, n6462);
  and g10887 (n6463, n_6041, n_6042);
  not g10888 (n_6043, n6439);
  not g10889 (n_6044, n6463);
  and g10890 (n6464, n_6043, n_6044);
  and g10891 (n6465, n_6037, n6458);
  and g10892 (n6466, n_6039, n6465);
  and g10893 (n6467, n_6038, n_6040);
  not g10894 (n_6045, n6466);
  not g10895 (n_6046, n6467);
  and g10896 (n6468, n_6045, n_6046);
  not g10897 (n_6047, n6468);
  and g10898 (n6469, n6439, n_6047);
  and g10899 (n6470, n_5908, n_5909);
  not g10900 (n_6048, n6469);
  and g10901 (n6471, n_6048, n6470);
  not g10902 (n_6049, n6464);
  and g10903 (n6472, n_6049, n6471);
  and g10904 (n6473, n_6049, n_6048);
  not g10905 (n_6050, n6470);
  not g10906 (n_6051, n6473);
  and g10907 (n6474, n_6050, n_6051);
  not g10908 (n_6052, n6472);
  not g10909 (n_6053, n6474);
  and g10910 (n6475, n_6052, n_6053);
  and g10911 (n6476, n_5806, n_5804);
  not g10912 (n_6054, n6476);
  and g10913 (n6477, n_5805, n_6054);
  and g10914 (n6478, n_5762, n_5806);
  and g10915 (n6479, n_5763, n6478);
  and g10916 (n6480, n_5807, n6479);
  and g10917 (n6481, n_5762, n_5760);
  not g10918 (n_6055, n6481);
  and g10919 (n6482, n_5761, n_6055);
  not g10920 (n_6056, n6480);
  not g10921 (n_6057, n6482);
  and g10922 (n6483, n_6056, n_6057);
  not g10927 (n_6058, n6483);
  not g10928 (n_6059, n6487);
  and g10929 (n6488, n_6058, n_6059);
  not g10930 (n_6060, n6488);
  and g10931 (n6489, n6477, n_6060);
  and g10932 (n6490, n_6056, n6482);
  and g10933 (n6491, n6480, n_6057);
  not g10934 (n_6061, n6490);
  not g10935 (n_6062, n6491);
  and g10936 (n6492, n_6061, n_6062);
  not g10937 (n_6063, n6477);
  not g10938 (n_6064, n6492);
  and g10939 (n6493, n_6063, n_6064);
  and g10940 (n6494, n_5904, n_5905);
  not g10941 (n_6065, n6493);
  and g10942 (n6495, n_6065, n6494);
  not g10943 (n_6066, n6489);
  and g10944 (n6496, n_6066, n6495);
  and g10945 (n6497, n_6066, n_6065);
  not g10946 (n_6067, n6494);
  not g10947 (n_6068, n6497);
  and g10948 (n6498, n_6067, n_6068);
  not g10949 (n_6069, n6496);
  not g10950 (n_6070, n6498);
  and g10951 (n6499, n_6069, n_6070);
  and g10952 (n6500, n_5898, n_5896);
  not g10953 (n_6071, n6500);
  and g10954 (n6501, n_5897, n_6071);
  and g10955 (n6502, n_5854, n_5898);
  and g10956 (n6503, n_5855, n6502);
  and g10957 (n6504, n_5899, n6503);
  and g10958 (n6505, n_5854, n_5852);
  not g10959 (n_6072, n6505);
  and g10960 (n6506, n_5853, n_6072);
  not g10961 (n_6073, n6504);
  and g10962 (n6507, n_6073, n6506);
  not g10963 (n_6074, n6506);
  and g10964 (n6508, n6504, n_6074);
  not g10965 (n_6075, n6507);
  not g10966 (n_6076, n6508);
  and g10967 (n6509, n_6075, n_6076);
  not g10968 (n_6077, n6501);
  not g10969 (n_6078, n6509);
  and g10970 (n6510, n_6077, n_6078);
  and g10971 (n6511, n_6073, n_6074);
  not g10976 (n_6079, n6511);
  not g10977 (n_6080, n6515);
  and g10978 (n6516, n_6079, n_6080);
  not g10979 (n_6081, n6516);
  and g10980 (n6517, n6501, n_6081);
  not g10981 (n_6082, n6510);
  not g10982 (n_6083, n6517);
  and g10983 (n6518, n_6082, n_6083);
  not g10984 (n_6084, n6499);
  and g10985 (n6519, n_6084, n6518);
  and g10986 (n6520, n_6065, n_6067);
  and g10987 (n6521, n_6066, n6520);
  and g10988 (n6522, n6494, n_6068);
  not g10989 (n_6085, n6521);
  not g10990 (n_6086, n6522);
  and g10991 (n6523, n_6085, n_6086);
  not g10992 (n_6087, n6518);
  not g10993 (n_6088, n6523);
  and g10994 (n6524, n_6087, n_6088);
  not g10995 (n_6089, n6519);
  not g10996 (n_6090, n6524);
  and g10997 (n6525, n_6089, n_6090);
  not g10998 (n_6091, n6475);
  and g10999 (n6526, n_6091, n6525);
  and g11000 (n6527, n_6048, n_6050);
  and g11001 (n6528, n_6049, n6527);
  and g11002 (n6529, n6470, n_6051);
  not g11003 (n_6092, n6528);
  not g11004 (n_6093, n6529);
  and g11005 (n6530, n_6092, n_6093);
  not g11006 (n_6094, n6525);
  not g11007 (n_6095, n6530);
  and g11008 (n6531, n_6094, n_6095);
  not g11009 (n_6096, n6526);
  not g11010 (n_6097, n6531);
  and g11011 (n6532, n_6096, n_6097);
  not g11012 (n_6098, n6420);
  and g11013 (n6533, n_6098, n6532);
  and g11014 (n6534, n_6007, n_6009);
  and g11015 (n6535, n_6008, n6534);
  and g11016 (n6536, n6415, n_6010);
  not g11017 (n_6099, n6535);
  not g11018 (n_6100, n6536);
  and g11019 (n6537, n_6099, n_6100);
  not g11020 (n_6101, n6532);
  not g11021 (n_6102, n6537);
  and g11022 (n6538, n_6101, n_6102);
  not g11023 (n_6103, n6533);
  not g11024 (n_6104, n6538);
  and g11025 (n6539, n_6103, n_6104);
  not g11026 (n_6105, n6303);
  and g11027 (n6540, n_6105, n6539);
  and g11028 (n6541, n_5918, n_5920);
  and g11029 (n6542, n_5919, n6541);
  and g11030 (n6543, n6298, n_5921);
  not g11031 (n_6106, n6542);
  not g11032 (n_6107, n6543);
  and g11033 (n6544, n_6106, n_6107);
  not g11034 (n_6108, n6539);
  not g11035 (n_6109, n6544);
  and g11036 (n6545, n_6108, n_6109);
  not g11037 (n_6110, n6540);
  not g11038 (n_6111, n6545);
  and g11039 (n6546, n_6110, n_6111);
  and g11040 (n6547, \A[202] , \A[203] );
  not g11041 (n_6114, \A[203] );
  and g11042 (n6548, \A[202] , n_6114);
  not g11043 (n_6115, \A[202] );
  and g11044 (n6549, n_6115, \A[203] );
  not g11045 (n_6116, n6548);
  not g11046 (n_6117, n6549);
  and g11047 (n6550, n_6116, n_6117);
  not g11048 (n_6119, n6550);
  and g11049 (n6551, \A[204] , n_6119);
  not g11050 (n_6120, n6547);
  not g11051 (n_6121, n6551);
  and g11052 (n6552, n_6120, n_6121);
  and g11053 (n6553, \A[199] , \A[200] );
  not g11054 (n_6124, \A[200] );
  and g11055 (n6554, \A[199] , n_6124);
  not g11056 (n_6125, \A[199] );
  and g11057 (n6555, n_6125, \A[200] );
  not g11058 (n_6126, n6554);
  not g11059 (n_6127, n6555);
  and g11060 (n6556, n_6126, n_6127);
  not g11061 (n_6129, n6556);
  and g11062 (n6557, \A[201] , n_6129);
  not g11063 (n_6130, n6553);
  not g11064 (n_6131, n6557);
  and g11065 (n6558, n_6130, n_6131);
  not g11066 (n_6132, n6558);
  and g11067 (n6559, n6552, n_6132);
  not g11068 (n_6133, n6552);
  and g11069 (n6560, n_6133, n6558);
  and g11070 (n6561, \A[201] , n_6126);
  and g11071 (n6562, n_6127, n6561);
  not g11072 (n_6134, \A[201] );
  and g11073 (n6563, n_6134, n_6129);
  not g11074 (n_6135, n6562);
  not g11075 (n_6136, n6563);
  and g11076 (n6564, n_6135, n_6136);
  and g11077 (n6565, \A[204] , n_6116);
  and g11078 (n6566, n_6117, n6565);
  not g11079 (n_6137, \A[204] );
  and g11080 (n6567, n_6137, n_6119);
  not g11081 (n_6138, n6566);
  not g11082 (n_6139, n6567);
  and g11083 (n6568, n_6138, n_6139);
  not g11084 (n_6140, n6564);
  not g11085 (n_6141, n6568);
  and g11086 (n6569, n_6140, n_6141);
  not g11087 (n_6142, n6560);
  and g11088 (n6570, n_6142, n6569);
  not g11089 (n_6143, n6559);
  and g11090 (n6571, n_6143, n6570);
  and g11091 (n6572, n_6143, n_6142);
  not g11092 (n_6144, n6569);
  not g11093 (n_6145, n6572);
  and g11094 (n6573, n_6144, n_6145);
  not g11095 (n_6146, n6571);
  not g11096 (n_6147, n6573);
  and g11097 (n6574, n_6146, n_6147);
  and g11098 (n6575, n_6140, n6568);
  and g11099 (n6576, n6564, n_6141);
  not g11100 (n_6148, n6575);
  not g11101 (n_6149, n6576);
  and g11102 (n6577, n_6148, n_6149);
  and g11103 (n6578, n6569, n_6145);
  and g11104 (n6579, n_6133, n_6132);
  not g11105 (n_6150, n6578);
  not g11106 (n_6151, n6579);
  and g11107 (n6580, n_6150, n_6151);
  not g11108 (n_6152, n6577);
  not g11109 (n_6153, n6580);
  and g11110 (n6581, n_6152, n_6153);
  not g11111 (n_6154, n6574);
  not g11112 (n_6155, n6581);
  and g11113 (n6582, n_6154, n_6155);
  and g11114 (n6583, n_6154, n_6153);
  and g11115 (n6584, \A[208] , \A[209] );
  not g11116 (n_6158, \A[209] );
  and g11117 (n6585, \A[208] , n_6158);
  not g11118 (n_6159, \A[208] );
  and g11119 (n6586, n_6159, \A[209] );
  not g11120 (n_6160, n6585);
  not g11121 (n_6161, n6586);
  and g11122 (n6587, n_6160, n_6161);
  not g11123 (n_6163, n6587);
  and g11124 (n6588, \A[210] , n_6163);
  not g11125 (n_6164, n6584);
  not g11126 (n_6165, n6588);
  and g11127 (n6589, n_6164, n_6165);
  and g11128 (n6590, \A[205] , \A[206] );
  not g11129 (n_6168, \A[206] );
  and g11130 (n6591, \A[205] , n_6168);
  not g11131 (n_6169, \A[205] );
  and g11132 (n6592, n_6169, \A[206] );
  not g11133 (n_6170, n6591);
  not g11134 (n_6171, n6592);
  and g11135 (n6593, n_6170, n_6171);
  not g11136 (n_6173, n6593);
  and g11137 (n6594, \A[207] , n_6173);
  not g11138 (n_6174, n6590);
  not g11139 (n_6175, n6594);
  and g11140 (n6595, n_6174, n_6175);
  not g11141 (n_6176, n6589);
  and g11142 (n6596, n_6176, n6595);
  not g11143 (n_6177, n6595);
  and g11144 (n6597, n6589, n_6177);
  not g11145 (n_6178, n6596);
  not g11146 (n_6179, n6597);
  and g11147 (n6598, n_6178, n_6179);
  and g11148 (n6599, \A[207] , n_6170);
  and g11149 (n6600, n_6171, n6599);
  not g11150 (n_6180, \A[207] );
  and g11151 (n6601, n_6180, n_6173);
  not g11152 (n_6181, n6600);
  not g11153 (n_6182, n6601);
  and g11154 (n6602, n_6181, n_6182);
  and g11155 (n6603, \A[210] , n_6160);
  and g11156 (n6604, n_6161, n6603);
  not g11157 (n_6183, \A[210] );
  and g11158 (n6605, n_6183, n_6163);
  not g11159 (n_6184, n6604);
  not g11160 (n_6185, n6605);
  and g11161 (n6606, n_6184, n_6185);
  not g11162 (n_6186, n6602);
  not g11163 (n_6187, n6606);
  and g11164 (n6607, n_6186, n_6187);
  not g11165 (n_6188, n6598);
  and g11166 (n6608, n_6188, n6607);
  and g11167 (n6609, n_6176, n_6177);
  not g11168 (n_6189, n6608);
  not g11169 (n_6190, n6609);
  and g11170 (n6610, n_6189, n_6190);
  and g11171 (n6611, n_6178, n6607);
  and g11172 (n6612, n_6179, n6611);
  not g11173 (n_6191, n6607);
  and g11174 (n6613, n_6188, n_6191);
  not g11175 (n_6192, n6612);
  not g11176 (n_6193, n6613);
  and g11177 (n6614, n_6192, n_6193);
  not g11178 (n_6194, n6610);
  not g11179 (n_6195, n6614);
  and g11180 (n6615, n_6194, n_6195);
  and g11181 (n6616, n_6186, n6606);
  and g11182 (n6617, n6602, n_6187);
  not g11183 (n_6196, n6616);
  not g11184 (n_6197, n6617);
  and g11185 (n6618, n_6196, n_6197);
  not g11186 (n_6198, n6618);
  and g11187 (n6619, n_6152, n_6198);
  not g11188 (n_6199, n6615);
  and g11189 (n6620, n_6199, n6619);
  not g11190 (n_6200, n6583);
  and g11191 (n6621, n_6200, n6620);
  and g11192 (n6622, n_6194, n_6198);
  not g11193 (n_6201, n6622);
  and g11194 (n6623, n_6195, n_6201);
  not g11195 (n_6202, n6621);
  and g11196 (n6624, n_6202, n6623);
  not g11197 (n_6203, n6623);
  and g11198 (n6625, n6621, n_6203);
  not g11199 (n_6204, n6624);
  not g11200 (n_6205, n6625);
  and g11201 (n6626, n_6204, n_6205);
  not g11202 (n_6206, n6582);
  not g11203 (n_6207, n6626);
  and g11204 (n6627, n_6206, n_6207);
  and g11205 (n6628, n_6202, n_6203);
  not g11210 (n_6208, n6628);
  not g11211 (n_6209, n6632);
  and g11212 (n6633, n_6208, n_6209);
  not g11213 (n_6210, n6633);
  and g11214 (n6634, n6582, n_6210);
  not g11215 (n_6211, n6627);
  not g11216 (n_6212, n6634);
  and g11217 (n6635, n_6211, n_6212);
  and g11218 (n6636, \A[214] , \A[215] );
  not g11219 (n_6215, \A[215] );
  and g11220 (n6637, \A[214] , n_6215);
  not g11221 (n_6216, \A[214] );
  and g11222 (n6638, n_6216, \A[215] );
  not g11223 (n_6217, n6637);
  not g11224 (n_6218, n6638);
  and g11225 (n6639, n_6217, n_6218);
  not g11226 (n_6220, n6639);
  and g11227 (n6640, \A[216] , n_6220);
  not g11228 (n_6221, n6636);
  not g11229 (n_6222, n6640);
  and g11230 (n6641, n_6221, n_6222);
  and g11231 (n6642, \A[211] , \A[212] );
  not g11232 (n_6225, \A[212] );
  and g11233 (n6643, \A[211] , n_6225);
  not g11234 (n_6226, \A[211] );
  and g11235 (n6644, n_6226, \A[212] );
  not g11236 (n_6227, n6643);
  not g11237 (n_6228, n6644);
  and g11238 (n6645, n_6227, n_6228);
  not g11239 (n_6230, n6645);
  and g11240 (n6646, \A[213] , n_6230);
  not g11241 (n_6231, n6642);
  not g11242 (n_6232, n6646);
  and g11243 (n6647, n_6231, n_6232);
  not g11244 (n_6233, n6647);
  and g11245 (n6648, n6641, n_6233);
  not g11246 (n_6234, n6641);
  and g11247 (n6649, n_6234, n6647);
  and g11248 (n6650, \A[213] , n_6227);
  and g11249 (n6651, n_6228, n6650);
  not g11250 (n_6235, \A[213] );
  and g11251 (n6652, n_6235, n_6230);
  not g11252 (n_6236, n6651);
  not g11253 (n_6237, n6652);
  and g11254 (n6653, n_6236, n_6237);
  and g11255 (n6654, \A[216] , n_6217);
  and g11256 (n6655, n_6218, n6654);
  not g11257 (n_6238, \A[216] );
  and g11258 (n6656, n_6238, n_6220);
  not g11259 (n_6239, n6655);
  not g11260 (n_6240, n6656);
  and g11261 (n6657, n_6239, n_6240);
  not g11262 (n_6241, n6653);
  not g11263 (n_6242, n6657);
  and g11264 (n6658, n_6241, n_6242);
  not g11265 (n_6243, n6649);
  and g11266 (n6659, n_6243, n6658);
  not g11267 (n_6244, n6648);
  and g11268 (n6660, n_6244, n6659);
  and g11269 (n6661, n_6244, n_6243);
  not g11270 (n_6245, n6658);
  not g11271 (n_6246, n6661);
  and g11272 (n6662, n_6245, n_6246);
  not g11273 (n_6247, n6660);
  not g11274 (n_6248, n6662);
  and g11275 (n6663, n_6247, n_6248);
  and g11276 (n6664, n_6241, n6657);
  and g11277 (n6665, n6653, n_6242);
  not g11278 (n_6249, n6664);
  not g11279 (n_6250, n6665);
  and g11280 (n6666, n_6249, n_6250);
  and g11281 (n6667, n6658, n_6246);
  and g11282 (n6668, n_6234, n_6233);
  not g11283 (n_6251, n6667);
  not g11284 (n_6252, n6668);
  and g11285 (n6669, n_6251, n_6252);
  not g11286 (n_6253, n6666);
  not g11287 (n_6254, n6669);
  and g11288 (n6670, n_6253, n_6254);
  not g11289 (n_6255, n6663);
  not g11290 (n_6256, n6670);
  and g11291 (n6671, n_6255, n_6256);
  and g11292 (n6672, n_6255, n_6254);
  and g11293 (n6673, \A[220] , \A[221] );
  not g11294 (n_6259, \A[221] );
  and g11295 (n6674, \A[220] , n_6259);
  not g11296 (n_6260, \A[220] );
  and g11297 (n6675, n_6260, \A[221] );
  not g11298 (n_6261, n6674);
  not g11299 (n_6262, n6675);
  and g11300 (n6676, n_6261, n_6262);
  not g11301 (n_6264, n6676);
  and g11302 (n6677, \A[222] , n_6264);
  not g11303 (n_6265, n6673);
  not g11304 (n_6266, n6677);
  and g11305 (n6678, n_6265, n_6266);
  and g11306 (n6679, \A[217] , \A[218] );
  not g11307 (n_6269, \A[218] );
  and g11308 (n6680, \A[217] , n_6269);
  not g11309 (n_6270, \A[217] );
  and g11310 (n6681, n_6270, \A[218] );
  not g11311 (n_6271, n6680);
  not g11312 (n_6272, n6681);
  and g11313 (n6682, n_6271, n_6272);
  not g11314 (n_6274, n6682);
  and g11315 (n6683, \A[219] , n_6274);
  not g11316 (n_6275, n6679);
  not g11317 (n_6276, n6683);
  and g11318 (n6684, n_6275, n_6276);
  not g11319 (n_6277, n6678);
  and g11320 (n6685, n_6277, n6684);
  not g11321 (n_6278, n6684);
  and g11322 (n6686, n6678, n_6278);
  not g11323 (n_6279, n6685);
  not g11324 (n_6280, n6686);
  and g11325 (n6687, n_6279, n_6280);
  and g11326 (n6688, \A[219] , n_6271);
  and g11327 (n6689, n_6272, n6688);
  not g11328 (n_6281, \A[219] );
  and g11329 (n6690, n_6281, n_6274);
  not g11330 (n_6282, n6689);
  not g11331 (n_6283, n6690);
  and g11332 (n6691, n_6282, n_6283);
  and g11333 (n6692, \A[222] , n_6261);
  and g11334 (n6693, n_6262, n6692);
  not g11335 (n_6284, \A[222] );
  and g11336 (n6694, n_6284, n_6264);
  not g11337 (n_6285, n6693);
  not g11338 (n_6286, n6694);
  and g11339 (n6695, n_6285, n_6286);
  not g11340 (n_6287, n6691);
  not g11341 (n_6288, n6695);
  and g11342 (n6696, n_6287, n_6288);
  not g11343 (n_6289, n6687);
  and g11344 (n6697, n_6289, n6696);
  and g11345 (n6698, n_6277, n_6278);
  not g11346 (n_6290, n6697);
  not g11347 (n_6291, n6698);
  and g11348 (n6699, n_6290, n_6291);
  and g11349 (n6700, n_6279, n6696);
  and g11350 (n6701, n_6280, n6700);
  not g11351 (n_6292, n6696);
  and g11352 (n6702, n_6289, n_6292);
  not g11353 (n_6293, n6701);
  not g11354 (n_6294, n6702);
  and g11355 (n6703, n_6293, n_6294);
  not g11356 (n_6295, n6699);
  not g11357 (n_6296, n6703);
  and g11358 (n6704, n_6295, n_6296);
  and g11359 (n6705, n_6287, n6695);
  and g11360 (n6706, n6691, n_6288);
  not g11361 (n_6297, n6705);
  not g11362 (n_6298, n6706);
  and g11363 (n6707, n_6297, n_6298);
  not g11364 (n_6299, n6707);
  and g11365 (n6708, n_6253, n_6299);
  not g11366 (n_6300, n6704);
  and g11367 (n6709, n_6300, n6708);
  not g11368 (n_6301, n6672);
  and g11369 (n6710, n_6301, n6709);
  and g11370 (n6711, n_6295, n_6299);
  not g11371 (n_6302, n6711);
  and g11372 (n6712, n_6296, n_6302);
  not g11373 (n_6303, n6710);
  not g11374 (n_6304, n6712);
  and g11375 (n6713, n_6303, n_6304);
  not g11380 (n_6305, n6713);
  not g11381 (n_6306, n6717);
  and g11382 (n6718, n_6305, n_6306);
  not g11383 (n_6307, n6718);
  and g11384 (n6719, n6671, n_6307);
  and g11385 (n6720, n_6303, n6712);
  and g11386 (n6721, n6710, n_6304);
  not g11387 (n_6308, n6720);
  not g11388 (n_6309, n6721);
  and g11389 (n6722, n_6308, n_6309);
  not g11390 (n_6310, n6671);
  not g11391 (n_6311, n6722);
  and g11392 (n6723, n_6310, n_6311);
  and g11393 (n6724, n_6300, n_6299);
  and g11394 (n6725, n_6253, n_6301);
  not g11395 (n_6312, n6724);
  and g11396 (n6726, n_6312, n6725);
  not g11397 (n_6313, n6725);
  and g11398 (n6727, n6724, n_6313);
  not g11399 (n_6314, n6726);
  not g11400 (n_6315, n6727);
  and g11401 (n6728, n_6314, n_6315);
  and g11402 (n6729, n_6199, n_6198);
  and g11403 (n6730, n_6152, n_6200);
  not g11404 (n_6316, n6729);
  and g11405 (n6731, n_6316, n6730);
  not g11406 (n_6317, n6730);
  and g11407 (n6732, n6729, n_6317);
  not g11408 (n_6318, n6731);
  not g11409 (n_6319, n6732);
  and g11410 (n6733, n_6318, n_6319);
  not g11411 (n_6320, n6728);
  not g11412 (n_6321, n6733);
  and g11413 (n6734, n_6320, n_6321);
  not g11414 (n_6322, n6723);
  not g11415 (n_6323, n6734);
  and g11416 (n6735, n_6322, n_6323);
  not g11417 (n_6324, n6719);
  and g11418 (n6736, n_6324, n6735);
  and g11419 (n6737, n_6324, n_6322);
  not g11420 (n_6325, n6737);
  and g11421 (n6738, n6734, n_6325);
  not g11422 (n_6326, n6736);
  not g11423 (n_6327, n6738);
  and g11424 (n6739, n_6326, n_6327);
  not g11425 (n_6328, n6635);
  not g11426 (n_6329, n6739);
  and g11427 (n6740, n_6328, n_6329);
  and g11428 (n6741, n_6322, n6734);
  and g11429 (n6742, n_6324, n6741);
  and g11430 (n6743, n_6323, n_6325);
  not g11431 (n_6330, n6742);
  not g11432 (n_6331, n6743);
  and g11433 (n6744, n_6330, n_6331);
  not g11434 (n_6332, n6744);
  and g11435 (n6745, n6635, n_6332);
  and g11436 (n6746, n_6320, n6733);
  and g11437 (n6747, n6728, n_6321);
  not g11438 (n_6333, n6746);
  not g11439 (n_6334, n6747);
  and g11440 (n6748, n_6333, n_6334);
  not g11441 (n_6336, \A[193] );
  and g11442 (n6749, n_6336, \A[194] );
  not g11443 (n_6338, \A[194] );
  and g11444 (n6750, \A[193] , n_6338);
  not g11445 (n_6340, n6750);
  and g11446 (n6751, \A[195] , n_6340);
  not g11447 (n_6341, n6749);
  and g11448 (n6752, n_6341, n6751);
  and g11449 (n6753, n_6341, n_6340);
  not g11450 (n_6342, \A[195] );
  not g11451 (n_6343, n6753);
  and g11452 (n6754, n_6342, n_6343);
  not g11453 (n_6344, n6752);
  not g11454 (n_6345, n6754);
  and g11455 (n6755, n_6344, n_6345);
  not g11456 (n_6347, \A[196] );
  and g11457 (n6756, n_6347, \A[197] );
  not g11458 (n_6349, \A[197] );
  and g11459 (n6757, \A[196] , n_6349);
  not g11460 (n_6351, n6757);
  and g11461 (n6758, \A[198] , n_6351);
  not g11462 (n_6352, n6756);
  and g11463 (n6759, n_6352, n6758);
  and g11464 (n6760, n_6352, n_6351);
  not g11465 (n_6353, \A[198] );
  not g11466 (n_6354, n6760);
  and g11467 (n6761, n_6353, n_6354);
  not g11468 (n_6355, n6759);
  not g11469 (n_6356, n6761);
  and g11470 (n6762, n_6355, n_6356);
  not g11471 (n_6357, n6755);
  and g11472 (n6763, n_6357, n6762);
  not g11473 (n_6358, n6762);
  and g11474 (n6764, n6755, n_6358);
  not g11475 (n_6359, n6763);
  not g11476 (n_6360, n6764);
  and g11477 (n6765, n_6359, n_6360);
  and g11478 (n6766, \A[196] , \A[197] );
  and g11479 (n6767, \A[198] , n_6354);
  not g11480 (n_6361, n6766);
  not g11481 (n_6362, n6767);
  and g11482 (n6768, n_6361, n_6362);
  and g11483 (n6769, \A[193] , \A[194] );
  and g11484 (n6770, \A[195] , n_6343);
  not g11485 (n_6363, n6769);
  not g11486 (n_6364, n6770);
  and g11487 (n6771, n_6363, n_6364);
  not g11488 (n_6365, n6768);
  and g11489 (n6772, n_6365, n6771);
  not g11490 (n_6366, n6771);
  and g11491 (n6773, n6768, n_6366);
  not g11492 (n_6367, n6772);
  not g11493 (n_6368, n6773);
  and g11494 (n6774, n_6367, n_6368);
  and g11495 (n6775, n_6357, n_6358);
  not g11496 (n_6369, n6774);
  and g11497 (n6776, n_6369, n6775);
  and g11498 (n6777, n_6365, n_6366);
  not g11499 (n_6370, n6776);
  not g11500 (n_6371, n6777);
  and g11501 (n6778, n_6370, n_6371);
  and g11502 (n6779, n_6367, n6775);
  and g11503 (n6780, n_6368, n6779);
  not g11504 (n_6372, n6775);
  and g11505 (n6781, n_6369, n_6372);
  not g11506 (n_6373, n6780);
  not g11507 (n_6374, n6781);
  and g11508 (n6782, n_6373, n_6374);
  not g11509 (n_6375, n6778);
  not g11510 (n_6376, n6782);
  and g11511 (n6783, n_6375, n_6376);
  not g11512 (n_6377, n6765);
  not g11513 (n_6378, n6783);
  and g11514 (n6784, n_6377, n_6378);
  not g11515 (n_6380, \A[187] );
  and g11516 (n6785, n_6380, \A[188] );
  not g11517 (n_6382, \A[188] );
  and g11518 (n6786, \A[187] , n_6382);
  not g11519 (n_6384, n6786);
  and g11520 (n6787, \A[189] , n_6384);
  not g11521 (n_6385, n6785);
  and g11522 (n6788, n_6385, n6787);
  and g11523 (n6789, n_6385, n_6384);
  not g11524 (n_6386, \A[189] );
  not g11525 (n_6387, n6789);
  and g11526 (n6790, n_6386, n_6387);
  not g11527 (n_6388, n6788);
  not g11528 (n_6389, n6790);
  and g11529 (n6791, n_6388, n_6389);
  not g11530 (n_6391, \A[190] );
  and g11531 (n6792, n_6391, \A[191] );
  not g11532 (n_6393, \A[191] );
  and g11533 (n6793, \A[190] , n_6393);
  not g11534 (n_6395, n6793);
  and g11535 (n6794, \A[192] , n_6395);
  not g11536 (n_6396, n6792);
  and g11537 (n6795, n_6396, n6794);
  and g11538 (n6796, n_6396, n_6395);
  not g11539 (n_6397, \A[192] );
  not g11540 (n_6398, n6796);
  and g11541 (n6797, n_6397, n_6398);
  not g11542 (n_6399, n6795);
  not g11543 (n_6400, n6797);
  and g11544 (n6798, n_6399, n_6400);
  not g11545 (n_6401, n6791);
  and g11546 (n6799, n_6401, n6798);
  not g11547 (n_6402, n6798);
  and g11548 (n6800, n6791, n_6402);
  not g11549 (n_6403, n6799);
  not g11550 (n_6404, n6800);
  and g11551 (n6801, n_6403, n_6404);
  and g11552 (n6802, \A[190] , \A[191] );
  and g11553 (n6803, \A[192] , n_6398);
  not g11554 (n_6405, n6802);
  not g11555 (n_6406, n6803);
  and g11556 (n6804, n_6405, n_6406);
  and g11557 (n6805, \A[187] , \A[188] );
  and g11558 (n6806, \A[189] , n_6387);
  not g11559 (n_6407, n6805);
  not g11560 (n_6408, n6806);
  and g11561 (n6807, n_6407, n_6408);
  not g11562 (n_6409, n6804);
  and g11563 (n6808, n_6409, n6807);
  not g11564 (n_6410, n6807);
  and g11565 (n6809, n6804, n_6410);
  not g11566 (n_6411, n6808);
  not g11567 (n_6412, n6809);
  and g11568 (n6810, n_6411, n_6412);
  and g11569 (n6811, n_6401, n_6402);
  not g11570 (n_6413, n6810);
  and g11571 (n6812, n_6413, n6811);
  and g11572 (n6813, n_6409, n_6410);
  not g11573 (n_6414, n6812);
  not g11574 (n_6415, n6813);
  and g11575 (n6814, n_6414, n_6415);
  and g11576 (n6815, n_6411, n6811);
  and g11577 (n6816, n_6412, n6815);
  not g11578 (n_6416, n6811);
  and g11579 (n6817, n_6413, n_6416);
  not g11580 (n_6417, n6816);
  not g11581 (n_6418, n6817);
  and g11582 (n6818, n_6417, n_6418);
  not g11583 (n_6419, n6814);
  not g11584 (n_6420, n6818);
  and g11585 (n6819, n_6419, n_6420);
  not g11586 (n_6421, n6801);
  not g11587 (n_6422, n6819);
  and g11588 (n6820, n_6421, n_6422);
  not g11589 (n_6423, n6784);
  and g11590 (n6821, n_6423, n6820);
  not g11591 (n_6424, n6820);
  and g11592 (n6822, n6784, n_6424);
  not g11593 (n_6425, n6821);
  not g11594 (n_6426, n6822);
  and g11595 (n6823, n_6425, n_6426);
  not g11596 (n_6428, \A[181] );
  and g11597 (n6824, n_6428, \A[182] );
  not g11598 (n_6430, \A[182] );
  and g11599 (n6825, \A[181] , n_6430);
  not g11600 (n_6432, n6825);
  and g11601 (n6826, \A[183] , n_6432);
  not g11602 (n_6433, n6824);
  and g11603 (n6827, n_6433, n6826);
  and g11604 (n6828, n_6433, n_6432);
  not g11605 (n_6434, \A[183] );
  not g11606 (n_6435, n6828);
  and g11607 (n6829, n_6434, n_6435);
  not g11608 (n_6436, n6827);
  not g11609 (n_6437, n6829);
  and g11610 (n6830, n_6436, n_6437);
  not g11611 (n_6439, \A[184] );
  and g11612 (n6831, n_6439, \A[185] );
  not g11613 (n_6441, \A[185] );
  and g11614 (n6832, \A[184] , n_6441);
  not g11615 (n_6443, n6832);
  and g11616 (n6833, \A[186] , n_6443);
  not g11617 (n_6444, n6831);
  and g11618 (n6834, n_6444, n6833);
  and g11619 (n6835, n_6444, n_6443);
  not g11620 (n_6445, \A[186] );
  not g11621 (n_6446, n6835);
  and g11622 (n6836, n_6445, n_6446);
  not g11623 (n_6447, n6834);
  not g11624 (n_6448, n6836);
  and g11625 (n6837, n_6447, n_6448);
  not g11626 (n_6449, n6830);
  and g11627 (n6838, n_6449, n6837);
  not g11628 (n_6450, n6837);
  and g11629 (n6839, n6830, n_6450);
  not g11630 (n_6451, n6838);
  not g11631 (n_6452, n6839);
  and g11632 (n6840, n_6451, n_6452);
  and g11633 (n6841, \A[184] , \A[185] );
  and g11634 (n6842, \A[186] , n_6446);
  not g11635 (n_6453, n6841);
  not g11636 (n_6454, n6842);
  and g11637 (n6843, n_6453, n_6454);
  and g11638 (n6844, \A[181] , \A[182] );
  and g11639 (n6845, \A[183] , n_6435);
  not g11640 (n_6455, n6844);
  not g11641 (n_6456, n6845);
  and g11642 (n6846, n_6455, n_6456);
  not g11643 (n_6457, n6843);
  and g11644 (n6847, n_6457, n6846);
  not g11645 (n_6458, n6846);
  and g11646 (n6848, n6843, n_6458);
  not g11647 (n_6459, n6847);
  not g11648 (n_6460, n6848);
  and g11649 (n6849, n_6459, n_6460);
  and g11650 (n6850, n_6449, n_6450);
  not g11651 (n_6461, n6849);
  and g11652 (n6851, n_6461, n6850);
  and g11653 (n6852, n_6457, n_6458);
  not g11654 (n_6462, n6851);
  not g11655 (n_6463, n6852);
  and g11656 (n6853, n_6462, n_6463);
  and g11657 (n6854, n_6459, n6850);
  and g11658 (n6855, n_6460, n6854);
  not g11659 (n_6464, n6850);
  and g11660 (n6856, n_6461, n_6464);
  not g11661 (n_6465, n6855);
  not g11662 (n_6466, n6856);
  and g11663 (n6857, n_6465, n_6466);
  not g11664 (n_6467, n6853);
  not g11665 (n_6468, n6857);
  and g11666 (n6858, n_6467, n_6468);
  not g11667 (n_6469, n6840);
  not g11668 (n_6470, n6858);
  and g11669 (n6859, n_6469, n_6470);
  not g11670 (n_6472, \A[175] );
  and g11671 (n6860, n_6472, \A[176] );
  not g11672 (n_6474, \A[176] );
  and g11673 (n6861, \A[175] , n_6474);
  not g11674 (n_6476, n6861);
  and g11675 (n6862, \A[177] , n_6476);
  not g11676 (n_6477, n6860);
  and g11677 (n6863, n_6477, n6862);
  and g11678 (n6864, n_6477, n_6476);
  not g11679 (n_6478, \A[177] );
  not g11680 (n_6479, n6864);
  and g11681 (n6865, n_6478, n_6479);
  not g11682 (n_6480, n6863);
  not g11683 (n_6481, n6865);
  and g11684 (n6866, n_6480, n_6481);
  not g11685 (n_6483, \A[178] );
  and g11686 (n6867, n_6483, \A[179] );
  not g11687 (n_6485, \A[179] );
  and g11688 (n6868, \A[178] , n_6485);
  not g11689 (n_6487, n6868);
  and g11690 (n6869, \A[180] , n_6487);
  not g11691 (n_6488, n6867);
  and g11692 (n6870, n_6488, n6869);
  and g11693 (n6871, n_6488, n_6487);
  not g11694 (n_6489, \A[180] );
  not g11695 (n_6490, n6871);
  and g11696 (n6872, n_6489, n_6490);
  not g11697 (n_6491, n6870);
  not g11698 (n_6492, n6872);
  and g11699 (n6873, n_6491, n_6492);
  not g11700 (n_6493, n6866);
  and g11701 (n6874, n_6493, n6873);
  not g11702 (n_6494, n6873);
  and g11703 (n6875, n6866, n_6494);
  not g11704 (n_6495, n6874);
  not g11705 (n_6496, n6875);
  and g11706 (n6876, n_6495, n_6496);
  and g11707 (n6877, \A[178] , \A[179] );
  and g11708 (n6878, \A[180] , n_6490);
  not g11709 (n_6497, n6877);
  not g11710 (n_6498, n6878);
  and g11711 (n6879, n_6497, n_6498);
  and g11712 (n6880, \A[175] , \A[176] );
  and g11713 (n6881, \A[177] , n_6479);
  not g11714 (n_6499, n6880);
  not g11715 (n_6500, n6881);
  and g11716 (n6882, n_6499, n_6500);
  not g11717 (n_6501, n6879);
  and g11718 (n6883, n_6501, n6882);
  not g11719 (n_6502, n6882);
  and g11720 (n6884, n6879, n_6502);
  not g11721 (n_6503, n6883);
  not g11722 (n_6504, n6884);
  and g11723 (n6885, n_6503, n_6504);
  and g11724 (n6886, n_6493, n_6494);
  not g11725 (n_6505, n6885);
  and g11726 (n6887, n_6505, n6886);
  and g11727 (n6888, n_6501, n_6502);
  not g11728 (n_6506, n6887);
  not g11729 (n_6507, n6888);
  and g11730 (n6889, n_6506, n_6507);
  and g11731 (n6890, n_6503, n6886);
  and g11732 (n6891, n_6504, n6890);
  not g11733 (n_6508, n6886);
  and g11734 (n6892, n_6505, n_6508);
  not g11735 (n_6509, n6891);
  not g11736 (n_6510, n6892);
  and g11737 (n6893, n_6509, n_6510);
  not g11738 (n_6511, n6889);
  not g11739 (n_6512, n6893);
  and g11740 (n6894, n_6511, n_6512);
  not g11741 (n_6513, n6876);
  not g11742 (n_6514, n6894);
  and g11743 (n6895, n_6513, n_6514);
  not g11744 (n_6515, n6859);
  and g11745 (n6896, n_6515, n6895);
  not g11746 (n_6516, n6895);
  and g11747 (n6897, n6859, n_6516);
  not g11748 (n_6517, n6896);
  not g11749 (n_6518, n6897);
  and g11750 (n6898, n_6517, n_6518);
  not g11751 (n_6519, n6823);
  and g11752 (n6899, n_6519, n6898);
  not g11753 (n_6520, n6898);
  and g11754 (n6900, n6823, n_6520);
  not g11755 (n_6521, n6899);
  not g11756 (n_6522, n6900);
  and g11757 (n6901, n_6521, n_6522);
  not g11758 (n_6523, n6748);
  not g11759 (n_6524, n6901);
  and g11760 (n6902, n_6523, n_6524);
  not g11761 (n_6525, n6745);
  and g11762 (n6903, n_6525, n6902);
  not g11763 (n_6526, n6740);
  and g11764 (n6904, n_6526, n6903);
  and g11765 (n6905, n_6526, n_6525);
  not g11766 (n_6527, n6902);
  not g11767 (n_6528, n6905);
  and g11768 (n6906, n_6527, n_6528);
  not g11769 (n_6529, n6904);
  not g11770 (n_6530, n6906);
  and g11771 (n6907, n_6529, n_6530);
  and g11772 (n6908, n_6421, n_6419);
  not g11773 (n_6531, n6908);
  and g11774 (n6909, n_6420, n_6531);
  and g11775 (n6910, n_6377, n_6421);
  and g11776 (n6911, n_6378, n6910);
  and g11777 (n6912, n_6422, n6911);
  and g11778 (n6913, n_6377, n_6375);
  not g11779 (n_6532, n6913);
  and g11780 (n6914, n_6376, n_6532);
  not g11781 (n_6533, n6912);
  not g11782 (n_6534, n6914);
  and g11783 (n6915, n_6533, n_6534);
  not g11788 (n_6535, n6915);
  not g11789 (n_6536, n6919);
  and g11790 (n6920, n_6535, n_6536);
  not g11791 (n_6537, n6920);
  and g11792 (n6921, n6909, n_6537);
  and g11793 (n6922, n_6533, n6914);
  and g11794 (n6923, n6912, n_6534);
  not g11795 (n_6538, n6922);
  not g11796 (n_6539, n6923);
  and g11797 (n6924, n_6538, n_6539);
  not g11798 (n_6540, n6909);
  not g11799 (n_6541, n6924);
  and g11800 (n6925, n_6540, n_6541);
  and g11801 (n6926, n_6519, n_6520);
  not g11802 (n_6542, n6925);
  and g11803 (n6927, n_6542, n6926);
  not g11804 (n_6543, n6921);
  and g11805 (n6928, n_6543, n6927);
  and g11806 (n6929, n_6543, n_6542);
  not g11807 (n_6544, n6926);
  not g11808 (n_6545, n6929);
  and g11809 (n6930, n_6544, n_6545);
  not g11810 (n_6546, n6928);
  not g11811 (n_6547, n6930);
  and g11812 (n6931, n_6546, n_6547);
  and g11813 (n6932, n_6513, n_6511);
  not g11814 (n_6548, n6932);
  and g11815 (n6933, n_6512, n_6548);
  and g11816 (n6934, n_6469, n_6513);
  and g11817 (n6935, n_6470, n6934);
  and g11818 (n6936, n_6514, n6935);
  and g11819 (n6937, n_6469, n_6467);
  not g11820 (n_6549, n6937);
  and g11821 (n6938, n_6468, n_6549);
  not g11822 (n_6550, n6936);
  and g11823 (n6939, n_6550, n6938);
  not g11824 (n_6551, n6938);
  and g11825 (n6940, n6936, n_6551);
  not g11826 (n_6552, n6939);
  not g11827 (n_6553, n6940);
  and g11828 (n6941, n_6552, n_6553);
  not g11829 (n_6554, n6933);
  not g11830 (n_6555, n6941);
  and g11831 (n6942, n_6554, n_6555);
  and g11832 (n6943, n_6550, n_6551);
  not g11837 (n_6556, n6943);
  not g11838 (n_6557, n6947);
  and g11839 (n6948, n_6556, n_6557);
  not g11840 (n_6558, n6948);
  and g11841 (n6949, n6933, n_6558);
  not g11842 (n_6559, n6942);
  not g11843 (n_6560, n6949);
  and g11844 (n6950, n_6559, n_6560);
  not g11845 (n_6561, n6931);
  and g11846 (n6951, n_6561, n6950);
  and g11847 (n6952, n_6542, n_6544);
  and g11848 (n6953, n_6543, n6952);
  and g11849 (n6954, n6926, n_6545);
  not g11850 (n_6562, n6953);
  not g11851 (n_6563, n6954);
  and g11852 (n6955, n_6562, n_6563);
  not g11853 (n_6564, n6950);
  not g11854 (n_6565, n6955);
  and g11855 (n6956, n_6564, n_6565);
  not g11856 (n_6566, n6951);
  not g11857 (n_6567, n6956);
  and g11858 (n6957, n_6566, n_6567);
  not g11859 (n_6568, n6907);
  and g11860 (n6958, n_6568, n6957);
  and g11861 (n6959, n_6525, n_6527);
  and g11862 (n6960, n_6526, n6959);
  and g11863 (n6961, n6902, n_6528);
  not g11864 (n_6569, n6960);
  not g11865 (n_6570, n6961);
  and g11866 (n6962, n_6569, n_6570);
  not g11867 (n_6571, n6957);
  not g11868 (n_6572, n6962);
  and g11869 (n6963, n_6571, n_6572);
  not g11870 (n_6573, n6958);
  not g11871 (n_6574, n6963);
  and g11872 (n6964, n_6573, n_6574);
  and g11873 (n6965, \A[238] , \A[239] );
  not g11874 (n_6577, \A[239] );
  and g11875 (n6966, \A[238] , n_6577);
  not g11876 (n_6578, \A[238] );
  and g11877 (n6967, n_6578, \A[239] );
  not g11878 (n_6579, n6966);
  not g11879 (n_6580, n6967);
  and g11880 (n6968, n_6579, n_6580);
  not g11881 (n_6582, n6968);
  and g11882 (n6969, \A[240] , n_6582);
  not g11883 (n_6583, n6965);
  not g11884 (n_6584, n6969);
  and g11885 (n6970, n_6583, n_6584);
  and g11886 (n6971, \A[235] , \A[236] );
  not g11887 (n_6587, \A[236] );
  and g11888 (n6972, \A[235] , n_6587);
  not g11889 (n_6588, \A[235] );
  and g11890 (n6973, n_6588, \A[236] );
  not g11891 (n_6589, n6972);
  not g11892 (n_6590, n6973);
  and g11893 (n6974, n_6589, n_6590);
  not g11894 (n_6592, n6974);
  and g11895 (n6975, \A[237] , n_6592);
  not g11896 (n_6593, n6971);
  not g11897 (n_6594, n6975);
  and g11898 (n6976, n_6593, n_6594);
  not g11899 (n_6595, n6976);
  and g11900 (n6977, n6970, n_6595);
  not g11901 (n_6596, n6970);
  and g11902 (n6978, n_6596, n6976);
  and g11903 (n6979, \A[237] , n_6589);
  and g11904 (n6980, n_6590, n6979);
  not g11905 (n_6597, \A[237] );
  and g11906 (n6981, n_6597, n_6592);
  not g11907 (n_6598, n6980);
  not g11908 (n_6599, n6981);
  and g11909 (n6982, n_6598, n_6599);
  and g11910 (n6983, \A[240] , n_6579);
  and g11911 (n6984, n_6580, n6983);
  not g11912 (n_6600, \A[240] );
  and g11913 (n6985, n_6600, n_6582);
  not g11914 (n_6601, n6984);
  not g11915 (n_6602, n6985);
  and g11916 (n6986, n_6601, n_6602);
  not g11917 (n_6603, n6982);
  not g11918 (n_6604, n6986);
  and g11919 (n6987, n_6603, n_6604);
  not g11920 (n_6605, n6978);
  and g11921 (n6988, n_6605, n6987);
  not g11922 (n_6606, n6977);
  and g11923 (n6989, n_6606, n6988);
  and g11924 (n6990, n_6606, n_6605);
  not g11925 (n_6607, n6987);
  not g11926 (n_6608, n6990);
  and g11927 (n6991, n_6607, n_6608);
  not g11928 (n_6609, n6989);
  not g11929 (n_6610, n6991);
  and g11930 (n6992, n_6609, n_6610);
  and g11931 (n6993, n_6603, n6986);
  and g11932 (n6994, n6982, n_6604);
  not g11933 (n_6611, n6993);
  not g11934 (n_6612, n6994);
  and g11935 (n6995, n_6611, n_6612);
  and g11936 (n6996, n6987, n_6608);
  and g11937 (n6997, n_6596, n_6595);
  not g11938 (n_6613, n6996);
  not g11939 (n_6614, n6997);
  and g11940 (n6998, n_6613, n_6614);
  not g11941 (n_6615, n6995);
  not g11942 (n_6616, n6998);
  and g11943 (n6999, n_6615, n_6616);
  not g11944 (n_6617, n6992);
  not g11945 (n_6618, n6999);
  and g11946 (n7000, n_6617, n_6618);
  and g11947 (n7001, n_6617, n_6616);
  and g11948 (n7002, \A[244] , \A[245] );
  not g11949 (n_6621, \A[245] );
  and g11950 (n7003, \A[244] , n_6621);
  not g11951 (n_6622, \A[244] );
  and g11952 (n7004, n_6622, \A[245] );
  not g11953 (n_6623, n7003);
  not g11954 (n_6624, n7004);
  and g11955 (n7005, n_6623, n_6624);
  not g11956 (n_6626, n7005);
  and g11957 (n7006, \A[246] , n_6626);
  not g11958 (n_6627, n7002);
  not g11959 (n_6628, n7006);
  and g11960 (n7007, n_6627, n_6628);
  and g11961 (n7008, \A[241] , \A[242] );
  not g11962 (n_6631, \A[242] );
  and g11963 (n7009, \A[241] , n_6631);
  not g11964 (n_6632, \A[241] );
  and g11965 (n7010, n_6632, \A[242] );
  not g11966 (n_6633, n7009);
  not g11967 (n_6634, n7010);
  and g11968 (n7011, n_6633, n_6634);
  not g11969 (n_6636, n7011);
  and g11970 (n7012, \A[243] , n_6636);
  not g11971 (n_6637, n7008);
  not g11972 (n_6638, n7012);
  and g11973 (n7013, n_6637, n_6638);
  not g11974 (n_6639, n7007);
  and g11975 (n7014, n_6639, n7013);
  not g11976 (n_6640, n7013);
  and g11977 (n7015, n7007, n_6640);
  not g11978 (n_6641, n7014);
  not g11979 (n_6642, n7015);
  and g11980 (n7016, n_6641, n_6642);
  and g11981 (n7017, \A[243] , n_6633);
  and g11982 (n7018, n_6634, n7017);
  not g11983 (n_6643, \A[243] );
  and g11984 (n7019, n_6643, n_6636);
  not g11985 (n_6644, n7018);
  not g11986 (n_6645, n7019);
  and g11987 (n7020, n_6644, n_6645);
  and g11988 (n7021, \A[246] , n_6623);
  and g11989 (n7022, n_6624, n7021);
  not g11990 (n_6646, \A[246] );
  and g11991 (n7023, n_6646, n_6626);
  not g11992 (n_6647, n7022);
  not g11993 (n_6648, n7023);
  and g11994 (n7024, n_6647, n_6648);
  not g11995 (n_6649, n7020);
  not g11996 (n_6650, n7024);
  and g11997 (n7025, n_6649, n_6650);
  not g11998 (n_6651, n7016);
  and g11999 (n7026, n_6651, n7025);
  and g12000 (n7027, n_6639, n_6640);
  not g12001 (n_6652, n7026);
  not g12002 (n_6653, n7027);
  and g12003 (n7028, n_6652, n_6653);
  and g12004 (n7029, n_6641, n7025);
  and g12005 (n7030, n_6642, n7029);
  not g12006 (n_6654, n7025);
  and g12007 (n7031, n_6651, n_6654);
  not g12008 (n_6655, n7030);
  not g12009 (n_6656, n7031);
  and g12010 (n7032, n_6655, n_6656);
  not g12011 (n_6657, n7028);
  not g12012 (n_6658, n7032);
  and g12013 (n7033, n_6657, n_6658);
  and g12014 (n7034, n_6649, n7024);
  and g12015 (n7035, n7020, n_6650);
  not g12016 (n_6659, n7034);
  not g12017 (n_6660, n7035);
  and g12018 (n7036, n_6659, n_6660);
  not g12019 (n_6661, n7036);
  and g12020 (n7037, n_6615, n_6661);
  not g12021 (n_6662, n7033);
  and g12022 (n7038, n_6662, n7037);
  not g12023 (n_6663, n7001);
  and g12024 (n7039, n_6663, n7038);
  and g12025 (n7040, n_6657, n_6661);
  not g12026 (n_6664, n7040);
  and g12027 (n7041, n_6658, n_6664);
  not g12028 (n_6665, n7039);
  not g12029 (n_6666, n7041);
  and g12030 (n7042, n_6665, n_6666);
  not g12035 (n_6667, n7042);
  not g12036 (n_6668, n7046);
  and g12037 (n7047, n_6667, n_6668);
  not g12038 (n_6669, n7047);
  and g12039 (n7048, n7000, n_6669);
  and g12040 (n7049, n_6665, n7041);
  and g12041 (n7050, n7039, n_6666);
  not g12042 (n_6670, n7049);
  not g12043 (n_6671, n7050);
  and g12044 (n7051, n_6670, n_6671);
  not g12045 (n_6672, n7000);
  not g12046 (n_6673, n7051);
  and g12047 (n7052, n_6672, n_6673);
  and g12048 (n7053, n_6662, n_6661);
  and g12049 (n7054, n_6615, n_6663);
  not g12050 (n_6674, n7053);
  and g12051 (n7055, n_6674, n7054);
  not g12052 (n_6675, n7054);
  and g12053 (n7056, n7053, n_6675);
  not g12054 (n_6676, n7055);
  not g12055 (n_6677, n7056);
  and g12056 (n7057, n_6676, n_6677);
  not g12057 (n_6679, \A[229] );
  and g12058 (n7058, n_6679, \A[230] );
  not g12059 (n_6681, \A[230] );
  and g12060 (n7059, \A[229] , n_6681);
  not g12061 (n_6683, n7059);
  and g12062 (n7060, \A[231] , n_6683);
  not g12063 (n_6684, n7058);
  and g12064 (n7061, n_6684, n7060);
  and g12065 (n7062, n_6684, n_6683);
  not g12066 (n_6685, \A[231] );
  not g12067 (n_6686, n7062);
  and g12068 (n7063, n_6685, n_6686);
  not g12069 (n_6687, n7061);
  not g12070 (n_6688, n7063);
  and g12071 (n7064, n_6687, n_6688);
  not g12072 (n_6690, \A[232] );
  and g12073 (n7065, n_6690, \A[233] );
  not g12074 (n_6692, \A[233] );
  and g12075 (n7066, \A[232] , n_6692);
  not g12076 (n_6694, n7066);
  and g12077 (n7067, \A[234] , n_6694);
  not g12078 (n_6695, n7065);
  and g12079 (n7068, n_6695, n7067);
  and g12080 (n7069, n_6695, n_6694);
  not g12081 (n_6696, \A[234] );
  not g12082 (n_6697, n7069);
  and g12083 (n7070, n_6696, n_6697);
  not g12084 (n_6698, n7068);
  not g12085 (n_6699, n7070);
  and g12086 (n7071, n_6698, n_6699);
  not g12087 (n_6700, n7064);
  and g12088 (n7072, n_6700, n7071);
  not g12089 (n_6701, n7071);
  and g12090 (n7073, n7064, n_6701);
  not g12091 (n_6702, n7072);
  not g12092 (n_6703, n7073);
  and g12093 (n7074, n_6702, n_6703);
  and g12094 (n7075, \A[232] , \A[233] );
  and g12095 (n7076, \A[234] , n_6697);
  not g12096 (n_6704, n7075);
  not g12097 (n_6705, n7076);
  and g12098 (n7077, n_6704, n_6705);
  and g12099 (n7078, \A[229] , \A[230] );
  and g12100 (n7079, \A[231] , n_6686);
  not g12101 (n_6706, n7078);
  not g12102 (n_6707, n7079);
  and g12103 (n7080, n_6706, n_6707);
  not g12104 (n_6708, n7077);
  and g12105 (n7081, n_6708, n7080);
  not g12106 (n_6709, n7080);
  and g12107 (n7082, n7077, n_6709);
  not g12108 (n_6710, n7081);
  not g12109 (n_6711, n7082);
  and g12110 (n7083, n_6710, n_6711);
  and g12111 (n7084, n_6700, n_6701);
  not g12112 (n_6712, n7083);
  and g12113 (n7085, n_6712, n7084);
  and g12114 (n7086, n_6708, n_6709);
  not g12115 (n_6713, n7085);
  not g12116 (n_6714, n7086);
  and g12117 (n7087, n_6713, n_6714);
  and g12118 (n7088, n_6710, n7084);
  and g12119 (n7089, n_6711, n7088);
  not g12120 (n_6715, n7084);
  and g12121 (n7090, n_6712, n_6715);
  not g12122 (n_6716, n7089);
  not g12123 (n_6717, n7090);
  and g12124 (n7091, n_6716, n_6717);
  not g12125 (n_6718, n7087);
  not g12126 (n_6719, n7091);
  and g12127 (n7092, n_6718, n_6719);
  not g12128 (n_6720, n7074);
  not g12129 (n_6721, n7092);
  and g12130 (n7093, n_6720, n_6721);
  not g12131 (n_6723, \A[223] );
  and g12132 (n7094, n_6723, \A[224] );
  not g12133 (n_6725, \A[224] );
  and g12134 (n7095, \A[223] , n_6725);
  not g12135 (n_6727, n7095);
  and g12136 (n7096, \A[225] , n_6727);
  not g12137 (n_6728, n7094);
  and g12138 (n7097, n_6728, n7096);
  and g12139 (n7098, n_6728, n_6727);
  not g12140 (n_6729, \A[225] );
  not g12141 (n_6730, n7098);
  and g12142 (n7099, n_6729, n_6730);
  not g12143 (n_6731, n7097);
  not g12144 (n_6732, n7099);
  and g12145 (n7100, n_6731, n_6732);
  not g12146 (n_6734, \A[226] );
  and g12147 (n7101, n_6734, \A[227] );
  not g12148 (n_6736, \A[227] );
  and g12149 (n7102, \A[226] , n_6736);
  not g12150 (n_6738, n7102);
  and g12151 (n7103, \A[228] , n_6738);
  not g12152 (n_6739, n7101);
  and g12153 (n7104, n_6739, n7103);
  and g12154 (n7105, n_6739, n_6738);
  not g12155 (n_6740, \A[228] );
  not g12156 (n_6741, n7105);
  and g12157 (n7106, n_6740, n_6741);
  not g12158 (n_6742, n7104);
  not g12159 (n_6743, n7106);
  and g12160 (n7107, n_6742, n_6743);
  not g12161 (n_6744, n7100);
  and g12162 (n7108, n_6744, n7107);
  not g12163 (n_6745, n7107);
  and g12164 (n7109, n7100, n_6745);
  not g12165 (n_6746, n7108);
  not g12166 (n_6747, n7109);
  and g12167 (n7110, n_6746, n_6747);
  and g12168 (n7111, \A[226] , \A[227] );
  and g12169 (n7112, \A[228] , n_6741);
  not g12170 (n_6748, n7111);
  not g12171 (n_6749, n7112);
  and g12172 (n7113, n_6748, n_6749);
  and g12173 (n7114, \A[223] , \A[224] );
  and g12174 (n7115, \A[225] , n_6730);
  not g12175 (n_6750, n7114);
  not g12176 (n_6751, n7115);
  and g12177 (n7116, n_6750, n_6751);
  not g12178 (n_6752, n7113);
  and g12179 (n7117, n_6752, n7116);
  not g12180 (n_6753, n7116);
  and g12181 (n7118, n7113, n_6753);
  not g12182 (n_6754, n7117);
  not g12183 (n_6755, n7118);
  and g12184 (n7119, n_6754, n_6755);
  and g12185 (n7120, n_6744, n_6745);
  not g12186 (n_6756, n7119);
  and g12187 (n7121, n_6756, n7120);
  and g12188 (n7122, n_6752, n_6753);
  not g12189 (n_6757, n7121);
  not g12190 (n_6758, n7122);
  and g12191 (n7123, n_6757, n_6758);
  and g12192 (n7124, n_6754, n7120);
  and g12193 (n7125, n_6755, n7124);
  not g12194 (n_6759, n7120);
  and g12195 (n7126, n_6756, n_6759);
  not g12196 (n_6760, n7125);
  not g12197 (n_6761, n7126);
  and g12198 (n7127, n_6760, n_6761);
  not g12199 (n_6762, n7123);
  not g12200 (n_6763, n7127);
  and g12201 (n7128, n_6762, n_6763);
  not g12202 (n_6764, n7110);
  not g12203 (n_6765, n7128);
  and g12204 (n7129, n_6764, n_6765);
  not g12205 (n_6766, n7093);
  and g12206 (n7130, n_6766, n7129);
  not g12207 (n_6767, n7129);
  and g12208 (n7131, n7093, n_6767);
  not g12209 (n_6768, n7130);
  not g12210 (n_6769, n7131);
  and g12211 (n7132, n_6768, n_6769);
  not g12212 (n_6770, n7057);
  not g12213 (n_6771, n7132);
  and g12214 (n7133, n_6770, n_6771);
  not g12215 (n_6772, n7052);
  and g12216 (n7134, n_6772, n7133);
  not g12217 (n_6773, n7048);
  and g12218 (n7135, n_6773, n7134);
  and g12219 (n7136, n_6773, n_6772);
  not g12220 (n_6774, n7133);
  not g12221 (n_6775, n7136);
  and g12222 (n7137, n_6774, n_6775);
  not g12223 (n_6776, n7135);
  not g12224 (n_6777, n7137);
  and g12225 (n7138, n_6776, n_6777);
  and g12226 (n7139, n_6764, n_6762);
  not g12227 (n_6778, n7139);
  and g12228 (n7140, n_6763, n_6778);
  and g12229 (n7141, n_6720, n_6764);
  and g12230 (n7142, n_6721, n7141);
  and g12231 (n7143, n_6765, n7142);
  and g12232 (n7144, n_6720, n_6718);
  not g12233 (n_6779, n7144);
  and g12234 (n7145, n_6719, n_6779);
  not g12235 (n_6780, n7143);
  and g12236 (n7146, n_6780, n7145);
  not g12237 (n_6781, n7145);
  and g12238 (n7147, n7143, n_6781);
  not g12239 (n_6782, n7146);
  not g12240 (n_6783, n7147);
  and g12241 (n7148, n_6782, n_6783);
  not g12242 (n_6784, n7140);
  not g12243 (n_6785, n7148);
  and g12244 (n7149, n_6784, n_6785);
  and g12245 (n7150, n_6780, n_6781);
  not g12250 (n_6786, n7150);
  not g12251 (n_6787, n7154);
  and g12252 (n7155, n_6786, n_6787);
  not g12253 (n_6788, n7155);
  and g12254 (n7156, n7140, n_6788);
  not g12255 (n_6789, n7149);
  not g12256 (n_6790, n7156);
  and g12257 (n7157, n_6789, n_6790);
  not g12258 (n_6791, n7138);
  and g12259 (n7158, n_6791, n7157);
  and g12260 (n7159, n_6772, n_6774);
  and g12261 (n7160, n_6773, n7159);
  and g12262 (n7161, n7133, n_6775);
  not g12263 (n_6792, n7160);
  not g12264 (n_6793, n7161);
  and g12265 (n7162, n_6792, n_6793);
  not g12266 (n_6794, n7157);
  not g12267 (n_6795, n7162);
  and g12268 (n7163, n_6794, n_6795);
  not g12269 (n_6796, n7158);
  not g12270 (n_6797, n7163);
  and g12271 (n7164, n_6796, n_6797);
  and g12272 (n7165, \A[250] , \A[251] );
  not g12273 (n_6800, \A[251] );
  and g12274 (n7166, \A[250] , n_6800);
  not g12275 (n_6801, \A[250] );
  and g12276 (n7167, n_6801, \A[251] );
  not g12277 (n_6802, n7166);
  not g12278 (n_6803, n7167);
  and g12279 (n7168, n_6802, n_6803);
  not g12280 (n_6805, n7168);
  and g12281 (n7169, \A[252] , n_6805);
  not g12282 (n_6806, n7165);
  not g12283 (n_6807, n7169);
  and g12284 (n7170, n_6806, n_6807);
  and g12285 (n7171, \A[247] , \A[248] );
  not g12286 (n_6810, \A[248] );
  and g12287 (n7172, \A[247] , n_6810);
  not g12288 (n_6811, \A[247] );
  and g12289 (n7173, n_6811, \A[248] );
  not g12290 (n_6812, n7172);
  not g12291 (n_6813, n7173);
  and g12292 (n7174, n_6812, n_6813);
  not g12293 (n_6815, n7174);
  and g12294 (n7175, \A[249] , n_6815);
  not g12295 (n_6816, n7171);
  not g12296 (n_6817, n7175);
  and g12297 (n7176, n_6816, n_6817);
  not g12298 (n_6818, n7176);
  and g12299 (n7177, n7170, n_6818);
  not g12300 (n_6819, n7170);
  and g12301 (n7178, n_6819, n7176);
  and g12302 (n7179, \A[249] , n_6812);
  and g12303 (n7180, n_6813, n7179);
  not g12304 (n_6820, \A[249] );
  and g12305 (n7181, n_6820, n_6815);
  not g12306 (n_6821, n7180);
  not g12307 (n_6822, n7181);
  and g12308 (n7182, n_6821, n_6822);
  and g12309 (n7183, \A[252] , n_6802);
  and g12310 (n7184, n_6803, n7183);
  not g12311 (n_6823, \A[252] );
  and g12312 (n7185, n_6823, n_6805);
  not g12313 (n_6824, n7184);
  not g12314 (n_6825, n7185);
  and g12315 (n7186, n_6824, n_6825);
  not g12316 (n_6826, n7182);
  not g12317 (n_6827, n7186);
  and g12318 (n7187, n_6826, n_6827);
  not g12319 (n_6828, n7178);
  and g12320 (n7188, n_6828, n7187);
  not g12321 (n_6829, n7177);
  and g12322 (n7189, n_6829, n7188);
  and g12323 (n7190, n_6829, n_6828);
  not g12324 (n_6830, n7187);
  not g12325 (n_6831, n7190);
  and g12326 (n7191, n_6830, n_6831);
  not g12327 (n_6832, n7189);
  not g12328 (n_6833, n7191);
  and g12329 (n7192, n_6832, n_6833);
  and g12330 (n7193, n_6826, n7186);
  and g12331 (n7194, n7182, n_6827);
  not g12332 (n_6834, n7193);
  not g12333 (n_6835, n7194);
  and g12334 (n7195, n_6834, n_6835);
  and g12335 (n7196, n7187, n_6831);
  and g12336 (n7197, n_6819, n_6818);
  not g12337 (n_6836, n7196);
  not g12338 (n_6837, n7197);
  and g12339 (n7198, n_6836, n_6837);
  not g12340 (n_6838, n7195);
  not g12341 (n_6839, n7198);
  and g12342 (n7199, n_6838, n_6839);
  not g12343 (n_6840, n7192);
  not g12344 (n_6841, n7199);
  and g12345 (n7200, n_6840, n_6841);
  and g12346 (n7201, n_6840, n_6839);
  and g12347 (n7202, \A[256] , \A[257] );
  not g12348 (n_6844, \A[257] );
  and g12349 (n7203, \A[256] , n_6844);
  not g12350 (n_6845, \A[256] );
  and g12351 (n7204, n_6845, \A[257] );
  not g12352 (n_6846, n7203);
  not g12353 (n_6847, n7204);
  and g12354 (n7205, n_6846, n_6847);
  not g12355 (n_6849, n7205);
  and g12356 (n7206, \A[258] , n_6849);
  not g12357 (n_6850, n7202);
  not g12358 (n_6851, n7206);
  and g12359 (n7207, n_6850, n_6851);
  and g12360 (n7208, \A[253] , \A[254] );
  not g12361 (n_6854, \A[254] );
  and g12362 (n7209, \A[253] , n_6854);
  not g12363 (n_6855, \A[253] );
  and g12364 (n7210, n_6855, \A[254] );
  not g12365 (n_6856, n7209);
  not g12366 (n_6857, n7210);
  and g12367 (n7211, n_6856, n_6857);
  not g12368 (n_6859, n7211);
  and g12369 (n7212, \A[255] , n_6859);
  not g12370 (n_6860, n7208);
  not g12371 (n_6861, n7212);
  and g12372 (n7213, n_6860, n_6861);
  not g12373 (n_6862, n7207);
  and g12374 (n7214, n_6862, n7213);
  not g12375 (n_6863, n7213);
  and g12376 (n7215, n7207, n_6863);
  not g12377 (n_6864, n7214);
  not g12378 (n_6865, n7215);
  and g12379 (n7216, n_6864, n_6865);
  and g12380 (n7217, \A[255] , n_6856);
  and g12381 (n7218, n_6857, n7217);
  not g12382 (n_6866, \A[255] );
  and g12383 (n7219, n_6866, n_6859);
  not g12384 (n_6867, n7218);
  not g12385 (n_6868, n7219);
  and g12386 (n7220, n_6867, n_6868);
  and g12387 (n7221, \A[258] , n_6846);
  and g12388 (n7222, n_6847, n7221);
  not g12389 (n_6869, \A[258] );
  and g12390 (n7223, n_6869, n_6849);
  not g12391 (n_6870, n7222);
  not g12392 (n_6871, n7223);
  and g12393 (n7224, n_6870, n_6871);
  not g12394 (n_6872, n7220);
  not g12395 (n_6873, n7224);
  and g12396 (n7225, n_6872, n_6873);
  not g12397 (n_6874, n7216);
  and g12398 (n7226, n_6874, n7225);
  and g12399 (n7227, n_6862, n_6863);
  not g12400 (n_6875, n7226);
  not g12401 (n_6876, n7227);
  and g12402 (n7228, n_6875, n_6876);
  and g12403 (n7229, n_6864, n7225);
  and g12404 (n7230, n_6865, n7229);
  not g12405 (n_6877, n7225);
  and g12406 (n7231, n_6874, n_6877);
  not g12407 (n_6878, n7230);
  not g12408 (n_6879, n7231);
  and g12409 (n7232, n_6878, n_6879);
  not g12410 (n_6880, n7228);
  not g12411 (n_6881, n7232);
  and g12412 (n7233, n_6880, n_6881);
  and g12413 (n7234, n_6872, n7224);
  and g12414 (n7235, n7220, n_6873);
  not g12415 (n_6882, n7234);
  not g12416 (n_6883, n7235);
  and g12417 (n7236, n_6882, n_6883);
  not g12418 (n_6884, n7236);
  and g12419 (n7237, n_6838, n_6884);
  not g12420 (n_6885, n7233);
  and g12421 (n7238, n_6885, n7237);
  not g12422 (n_6886, n7201);
  and g12423 (n7239, n_6886, n7238);
  and g12424 (n7240, n_6880, n_6884);
  not g12425 (n_6887, n7240);
  and g12426 (n7241, n_6881, n_6887);
  not g12427 (n_6888, n7239);
  and g12428 (n7242, n_6888, n7241);
  not g12429 (n_6889, n7241);
  and g12430 (n7243, n7239, n_6889);
  not g12431 (n_6890, n7242);
  not g12432 (n_6891, n7243);
  and g12433 (n7244, n_6890, n_6891);
  not g12434 (n_6892, n7200);
  not g12435 (n_6893, n7244);
  and g12436 (n7245, n_6892, n_6893);
  and g12437 (n7246, n_6888, n_6889);
  not g12442 (n_6894, n7246);
  not g12443 (n_6895, n7250);
  and g12444 (n7251, n_6894, n_6895);
  not g12445 (n_6896, n7251);
  and g12446 (n7252, n7200, n_6896);
  not g12447 (n_6897, n7245);
  not g12448 (n_6898, n7252);
  and g12449 (n7253, n_6897, n_6898);
  and g12450 (n7254, \A[262] , \A[263] );
  not g12451 (n_6901, \A[263] );
  and g12452 (n7255, \A[262] , n_6901);
  not g12453 (n_6902, \A[262] );
  and g12454 (n7256, n_6902, \A[263] );
  not g12455 (n_6903, n7255);
  not g12456 (n_6904, n7256);
  and g12457 (n7257, n_6903, n_6904);
  not g12458 (n_6906, n7257);
  and g12459 (n7258, \A[264] , n_6906);
  not g12460 (n_6907, n7254);
  not g12461 (n_6908, n7258);
  and g12462 (n7259, n_6907, n_6908);
  and g12463 (n7260, \A[259] , \A[260] );
  not g12464 (n_6911, \A[260] );
  and g12465 (n7261, \A[259] , n_6911);
  not g12466 (n_6912, \A[259] );
  and g12467 (n7262, n_6912, \A[260] );
  not g12468 (n_6913, n7261);
  not g12469 (n_6914, n7262);
  and g12470 (n7263, n_6913, n_6914);
  not g12471 (n_6916, n7263);
  and g12472 (n7264, \A[261] , n_6916);
  not g12473 (n_6917, n7260);
  not g12474 (n_6918, n7264);
  and g12475 (n7265, n_6917, n_6918);
  not g12476 (n_6919, n7265);
  and g12477 (n7266, n7259, n_6919);
  not g12478 (n_6920, n7259);
  and g12479 (n7267, n_6920, n7265);
  and g12480 (n7268, \A[261] , n_6913);
  and g12481 (n7269, n_6914, n7268);
  not g12482 (n_6921, \A[261] );
  and g12483 (n7270, n_6921, n_6916);
  not g12484 (n_6922, n7269);
  not g12485 (n_6923, n7270);
  and g12486 (n7271, n_6922, n_6923);
  and g12487 (n7272, \A[264] , n_6903);
  and g12488 (n7273, n_6904, n7272);
  not g12489 (n_6924, \A[264] );
  and g12490 (n7274, n_6924, n_6906);
  not g12491 (n_6925, n7273);
  not g12492 (n_6926, n7274);
  and g12493 (n7275, n_6925, n_6926);
  not g12494 (n_6927, n7271);
  not g12495 (n_6928, n7275);
  and g12496 (n7276, n_6927, n_6928);
  not g12497 (n_6929, n7267);
  and g12498 (n7277, n_6929, n7276);
  not g12499 (n_6930, n7266);
  and g12500 (n7278, n_6930, n7277);
  and g12501 (n7279, n_6930, n_6929);
  not g12502 (n_6931, n7276);
  not g12503 (n_6932, n7279);
  and g12504 (n7280, n_6931, n_6932);
  not g12505 (n_6933, n7278);
  not g12506 (n_6934, n7280);
  and g12507 (n7281, n_6933, n_6934);
  and g12508 (n7282, n_6927, n7275);
  and g12509 (n7283, n7271, n_6928);
  not g12510 (n_6935, n7282);
  not g12511 (n_6936, n7283);
  and g12512 (n7284, n_6935, n_6936);
  and g12513 (n7285, n7276, n_6932);
  and g12514 (n7286, n_6920, n_6919);
  not g12515 (n_6937, n7285);
  not g12516 (n_6938, n7286);
  and g12517 (n7287, n_6937, n_6938);
  not g12518 (n_6939, n7284);
  not g12519 (n_6940, n7287);
  and g12520 (n7288, n_6939, n_6940);
  not g12521 (n_6941, n7281);
  not g12522 (n_6942, n7288);
  and g12523 (n7289, n_6941, n_6942);
  and g12524 (n7290, n_6941, n_6940);
  and g12525 (n7291, \A[268] , \A[269] );
  not g12526 (n_6945, \A[269] );
  and g12527 (n7292, \A[268] , n_6945);
  not g12528 (n_6946, \A[268] );
  and g12529 (n7293, n_6946, \A[269] );
  not g12530 (n_6947, n7292);
  not g12531 (n_6948, n7293);
  and g12532 (n7294, n_6947, n_6948);
  not g12533 (n_6950, n7294);
  and g12534 (n7295, \A[270] , n_6950);
  not g12535 (n_6951, n7291);
  not g12536 (n_6952, n7295);
  and g12537 (n7296, n_6951, n_6952);
  and g12538 (n7297, \A[265] , \A[266] );
  not g12539 (n_6955, \A[266] );
  and g12540 (n7298, \A[265] , n_6955);
  not g12541 (n_6956, \A[265] );
  and g12542 (n7299, n_6956, \A[266] );
  not g12543 (n_6957, n7298);
  not g12544 (n_6958, n7299);
  and g12545 (n7300, n_6957, n_6958);
  not g12546 (n_6960, n7300);
  and g12547 (n7301, \A[267] , n_6960);
  not g12548 (n_6961, n7297);
  not g12549 (n_6962, n7301);
  and g12550 (n7302, n_6961, n_6962);
  not g12551 (n_6963, n7296);
  and g12552 (n7303, n_6963, n7302);
  not g12553 (n_6964, n7302);
  and g12554 (n7304, n7296, n_6964);
  not g12555 (n_6965, n7303);
  not g12556 (n_6966, n7304);
  and g12557 (n7305, n_6965, n_6966);
  and g12558 (n7306, \A[267] , n_6957);
  and g12559 (n7307, n_6958, n7306);
  not g12560 (n_6967, \A[267] );
  and g12561 (n7308, n_6967, n_6960);
  not g12562 (n_6968, n7307);
  not g12563 (n_6969, n7308);
  and g12564 (n7309, n_6968, n_6969);
  and g12565 (n7310, \A[270] , n_6947);
  and g12566 (n7311, n_6948, n7310);
  not g12567 (n_6970, \A[270] );
  and g12568 (n7312, n_6970, n_6950);
  not g12569 (n_6971, n7311);
  not g12570 (n_6972, n7312);
  and g12571 (n7313, n_6971, n_6972);
  not g12572 (n_6973, n7309);
  not g12573 (n_6974, n7313);
  and g12574 (n7314, n_6973, n_6974);
  not g12575 (n_6975, n7305);
  and g12576 (n7315, n_6975, n7314);
  and g12577 (n7316, n_6963, n_6964);
  not g12578 (n_6976, n7315);
  not g12579 (n_6977, n7316);
  and g12580 (n7317, n_6976, n_6977);
  and g12581 (n7318, n_6965, n7314);
  and g12582 (n7319, n_6966, n7318);
  not g12583 (n_6978, n7314);
  and g12584 (n7320, n_6975, n_6978);
  not g12585 (n_6979, n7319);
  not g12586 (n_6980, n7320);
  and g12587 (n7321, n_6979, n_6980);
  not g12588 (n_6981, n7317);
  not g12589 (n_6982, n7321);
  and g12590 (n7322, n_6981, n_6982);
  and g12591 (n7323, n_6973, n7313);
  and g12592 (n7324, n7309, n_6974);
  not g12593 (n_6983, n7323);
  not g12594 (n_6984, n7324);
  and g12595 (n7325, n_6983, n_6984);
  not g12596 (n_6985, n7325);
  and g12597 (n7326, n_6939, n_6985);
  not g12598 (n_6986, n7322);
  and g12599 (n7327, n_6986, n7326);
  not g12600 (n_6987, n7290);
  and g12601 (n7328, n_6987, n7327);
  and g12602 (n7329, n_6981, n_6985);
  not g12603 (n_6988, n7329);
  and g12604 (n7330, n_6982, n_6988);
  not g12605 (n_6989, n7328);
  not g12606 (n_6990, n7330);
  and g12607 (n7331, n_6989, n_6990);
  not g12612 (n_6991, n7331);
  not g12613 (n_6992, n7335);
  and g12614 (n7336, n_6991, n_6992);
  not g12615 (n_6993, n7336);
  and g12616 (n7337, n7289, n_6993);
  and g12617 (n7338, n_6989, n7330);
  and g12618 (n7339, n7328, n_6990);
  not g12619 (n_6994, n7338);
  not g12620 (n_6995, n7339);
  and g12621 (n7340, n_6994, n_6995);
  not g12622 (n_6996, n7289);
  not g12623 (n_6997, n7340);
  and g12624 (n7341, n_6996, n_6997);
  and g12625 (n7342, n_6986, n_6985);
  and g12626 (n7343, n_6939, n_6987);
  not g12627 (n_6998, n7342);
  and g12628 (n7344, n_6998, n7343);
  not g12629 (n_6999, n7343);
  and g12630 (n7345, n7342, n_6999);
  not g12631 (n_7000, n7344);
  not g12632 (n_7001, n7345);
  and g12633 (n7346, n_7000, n_7001);
  and g12634 (n7347, n_6885, n_6884);
  and g12635 (n7348, n_6838, n_6886);
  not g12636 (n_7002, n7347);
  and g12637 (n7349, n_7002, n7348);
  not g12638 (n_7003, n7348);
  and g12639 (n7350, n7347, n_7003);
  not g12640 (n_7004, n7349);
  not g12641 (n_7005, n7350);
  and g12642 (n7351, n_7004, n_7005);
  not g12643 (n_7006, n7346);
  not g12644 (n_7007, n7351);
  and g12645 (n7352, n_7006, n_7007);
  not g12646 (n_7008, n7341);
  not g12647 (n_7009, n7352);
  and g12648 (n7353, n_7008, n_7009);
  not g12649 (n_7010, n7337);
  and g12650 (n7354, n_7010, n7353);
  and g12651 (n7355, n_7010, n_7008);
  not g12652 (n_7011, n7355);
  and g12653 (n7356, n7352, n_7011);
  not g12654 (n_7012, n7354);
  not g12655 (n_7013, n7356);
  and g12656 (n7357, n_7012, n_7013);
  not g12657 (n_7014, n7253);
  not g12658 (n_7015, n7357);
  and g12659 (n7358, n_7014, n_7015);
  and g12660 (n7359, n_7008, n7352);
  and g12661 (n7360, n_7010, n7359);
  and g12662 (n7361, n_7009, n_7011);
  not g12663 (n_7016, n7360);
  not g12664 (n_7017, n7361);
  and g12665 (n7362, n_7016, n_7017);
  not g12666 (n_7018, n7362);
  and g12667 (n7363, n7253, n_7018);
  and g12668 (n7364, n_7006, n7351);
  and g12669 (n7365, n7346, n_7007);
  not g12670 (n_7019, n7364);
  not g12671 (n_7020, n7365);
  and g12672 (n7366, n_7019, n_7020);
  and g12673 (n7367, n_6770, n7132);
  and g12674 (n7368, n7057, n_6771);
  not g12675 (n_7021, n7367);
  not g12676 (n_7022, n7368);
  and g12677 (n7369, n_7021, n_7022);
  not g12678 (n_7023, n7366);
  not g12679 (n_7024, n7369);
  and g12680 (n7370, n_7023, n_7024);
  not g12681 (n_7025, n7363);
  not g12682 (n_7026, n7370);
  and g12683 (n7371, n_7025, n_7026);
  not g12684 (n_7027, n7358);
  and g12685 (n7372, n_7027, n7371);
  and g12686 (n7373, n_7027, n_7025);
  not g12687 (n_7028, n7373);
  and g12688 (n7374, n7370, n_7028);
  not g12689 (n_7029, n7372);
  not g12690 (n_7030, n7374);
  and g12691 (n7375, n_7029, n_7030);
  not g12692 (n_7031, n7164);
  not g12693 (n_7032, n7375);
  and g12694 (n7376, n_7031, n_7032);
  and g12695 (n7377, n_7025, n7370);
  and g12696 (n7378, n_7027, n7377);
  and g12697 (n7379, n_7026, n_7028);
  not g12698 (n_7033, n7378);
  not g12699 (n_7034, n7379);
  and g12700 (n7380, n_7033, n_7034);
  not g12701 (n_7035, n7380);
  and g12702 (n7381, n7164, n_7035);
  and g12703 (n7382, n_7023, n7369);
  and g12704 (n7383, n7366, n_7024);
  not g12705 (n_7036, n7382);
  not g12706 (n_7037, n7383);
  and g12707 (n7384, n_7036, n_7037);
  and g12708 (n7385, n_6523, n6901);
  and g12709 (n7386, n6748, n_6524);
  not g12710 (n_7038, n7385);
  not g12711 (n_7039, n7386);
  and g12712 (n7387, n_7038, n_7039);
  not g12713 (n_7040, n7384);
  not g12714 (n_7041, n7387);
  and g12715 (n7388, n_7040, n_7041);
  not g12716 (n_7042, n7381);
  not g12717 (n_7043, n7388);
  and g12718 (n7389, n_7042, n_7043);
  not g12719 (n_7044, n7376);
  and g12720 (n7390, n_7044, n7389);
  and g12721 (n7391, n_7044, n_7042);
  not g12722 (n_7045, n7391);
  and g12723 (n7392, n7388, n_7045);
  not g12724 (n_7046, n7390);
  not g12725 (n_7047, n7392);
  and g12726 (n7393, n_7046, n_7047);
  not g12727 (n_7048, n6964);
  not g12728 (n_7049, n7393);
  and g12729 (n7394, n_7048, n_7049);
  and g12730 (n7395, n_7042, n7388);
  and g12731 (n7396, n_7044, n7395);
  and g12732 (n7397, n_7043, n_7045);
  not g12733 (n_7050, n7396);
  not g12734 (n_7051, n7397);
  and g12735 (n7398, n_7050, n_7051);
  not g12736 (n_7052, n7398);
  and g12737 (n7399, n6964, n_7052);
  and g12738 (n7400, n_7040, n7387);
  and g12739 (n7401, n7384, n_7041);
  not g12740 (n_7053, n7400);
  not g12741 (n_7054, n7401);
  and g12742 (n7402, n_7053, n_7054);
  not g12743 (n_7056, \A[169] );
  and g12744 (n7403, n_7056, \A[170] );
  not g12745 (n_7058, \A[170] );
  and g12746 (n7404, \A[169] , n_7058);
  not g12747 (n_7060, n7404);
  and g12748 (n7405, \A[171] , n_7060);
  not g12749 (n_7061, n7403);
  and g12750 (n7406, n_7061, n7405);
  and g12751 (n7407, n_7061, n_7060);
  not g12752 (n_7062, \A[171] );
  not g12753 (n_7063, n7407);
  and g12754 (n7408, n_7062, n_7063);
  not g12755 (n_7064, n7406);
  not g12756 (n_7065, n7408);
  and g12757 (n7409, n_7064, n_7065);
  not g12758 (n_7067, \A[172] );
  and g12759 (n7410, n_7067, \A[173] );
  not g12760 (n_7069, \A[173] );
  and g12761 (n7411, \A[172] , n_7069);
  not g12762 (n_7071, n7411);
  and g12763 (n7412, \A[174] , n_7071);
  not g12764 (n_7072, n7410);
  and g12765 (n7413, n_7072, n7412);
  and g12766 (n7414, n_7072, n_7071);
  not g12767 (n_7073, \A[174] );
  not g12768 (n_7074, n7414);
  and g12769 (n7415, n_7073, n_7074);
  not g12770 (n_7075, n7413);
  not g12771 (n_7076, n7415);
  and g12772 (n7416, n_7075, n_7076);
  not g12773 (n_7077, n7409);
  and g12774 (n7417, n_7077, n7416);
  not g12775 (n_7078, n7416);
  and g12776 (n7418, n7409, n_7078);
  not g12777 (n_7079, n7417);
  not g12778 (n_7080, n7418);
  and g12779 (n7419, n_7079, n_7080);
  and g12780 (n7420, \A[172] , \A[173] );
  and g12781 (n7421, \A[174] , n_7074);
  not g12782 (n_7081, n7420);
  not g12783 (n_7082, n7421);
  and g12784 (n7422, n_7081, n_7082);
  and g12785 (n7423, \A[169] , \A[170] );
  and g12786 (n7424, \A[171] , n_7063);
  not g12787 (n_7083, n7423);
  not g12788 (n_7084, n7424);
  and g12789 (n7425, n_7083, n_7084);
  not g12790 (n_7085, n7422);
  and g12791 (n7426, n_7085, n7425);
  not g12792 (n_7086, n7425);
  and g12793 (n7427, n7422, n_7086);
  not g12794 (n_7087, n7426);
  not g12795 (n_7088, n7427);
  and g12796 (n7428, n_7087, n_7088);
  and g12797 (n7429, n_7077, n_7078);
  not g12798 (n_7089, n7428);
  and g12799 (n7430, n_7089, n7429);
  and g12800 (n7431, n_7085, n_7086);
  not g12801 (n_7090, n7430);
  not g12802 (n_7091, n7431);
  and g12803 (n7432, n_7090, n_7091);
  and g12804 (n7433, n_7087, n7429);
  and g12805 (n7434, n_7088, n7433);
  not g12806 (n_7092, n7429);
  and g12807 (n7435, n_7089, n_7092);
  not g12808 (n_7093, n7434);
  not g12809 (n_7094, n7435);
  and g12810 (n7436, n_7093, n_7094);
  not g12811 (n_7095, n7432);
  not g12812 (n_7096, n7436);
  and g12813 (n7437, n_7095, n_7096);
  not g12814 (n_7097, n7419);
  not g12815 (n_7098, n7437);
  and g12816 (n7438, n_7097, n_7098);
  not g12817 (n_7100, \A[163] );
  and g12818 (n7439, n_7100, \A[164] );
  not g12819 (n_7102, \A[164] );
  and g12820 (n7440, \A[163] , n_7102);
  not g12821 (n_7104, n7440);
  and g12822 (n7441, \A[165] , n_7104);
  not g12823 (n_7105, n7439);
  and g12824 (n7442, n_7105, n7441);
  and g12825 (n7443, n_7105, n_7104);
  not g12826 (n_7106, \A[165] );
  not g12827 (n_7107, n7443);
  and g12828 (n7444, n_7106, n_7107);
  not g12829 (n_7108, n7442);
  not g12830 (n_7109, n7444);
  and g12831 (n7445, n_7108, n_7109);
  not g12832 (n_7111, \A[166] );
  and g12833 (n7446, n_7111, \A[167] );
  not g12834 (n_7113, \A[167] );
  and g12835 (n7447, \A[166] , n_7113);
  not g12836 (n_7115, n7447);
  and g12837 (n7448, \A[168] , n_7115);
  not g12838 (n_7116, n7446);
  and g12839 (n7449, n_7116, n7448);
  and g12840 (n7450, n_7116, n_7115);
  not g12841 (n_7117, \A[168] );
  not g12842 (n_7118, n7450);
  and g12843 (n7451, n_7117, n_7118);
  not g12844 (n_7119, n7449);
  not g12845 (n_7120, n7451);
  and g12846 (n7452, n_7119, n_7120);
  not g12847 (n_7121, n7445);
  and g12848 (n7453, n_7121, n7452);
  not g12849 (n_7122, n7452);
  and g12850 (n7454, n7445, n_7122);
  not g12851 (n_7123, n7453);
  not g12852 (n_7124, n7454);
  and g12853 (n7455, n_7123, n_7124);
  and g12854 (n7456, \A[166] , \A[167] );
  and g12855 (n7457, \A[168] , n_7118);
  not g12856 (n_7125, n7456);
  not g12857 (n_7126, n7457);
  and g12858 (n7458, n_7125, n_7126);
  and g12859 (n7459, \A[163] , \A[164] );
  and g12860 (n7460, \A[165] , n_7107);
  not g12861 (n_7127, n7459);
  not g12862 (n_7128, n7460);
  and g12863 (n7461, n_7127, n_7128);
  not g12864 (n_7129, n7458);
  and g12865 (n7462, n_7129, n7461);
  not g12866 (n_7130, n7461);
  and g12867 (n7463, n7458, n_7130);
  not g12868 (n_7131, n7462);
  not g12869 (n_7132, n7463);
  and g12870 (n7464, n_7131, n_7132);
  and g12871 (n7465, n_7121, n_7122);
  not g12872 (n_7133, n7464);
  and g12873 (n7466, n_7133, n7465);
  and g12874 (n7467, n_7129, n_7130);
  not g12875 (n_7134, n7466);
  not g12876 (n_7135, n7467);
  and g12877 (n7468, n_7134, n_7135);
  and g12878 (n7469, n_7131, n7465);
  and g12879 (n7470, n_7132, n7469);
  not g12880 (n_7136, n7465);
  and g12881 (n7471, n_7133, n_7136);
  not g12882 (n_7137, n7470);
  not g12883 (n_7138, n7471);
  and g12884 (n7472, n_7137, n_7138);
  not g12885 (n_7139, n7468);
  not g12886 (n_7140, n7472);
  and g12887 (n7473, n_7139, n_7140);
  not g12888 (n_7141, n7455);
  not g12889 (n_7142, n7473);
  and g12890 (n7474, n_7141, n_7142);
  not g12891 (n_7143, n7438);
  and g12892 (n7475, n_7143, n7474);
  not g12893 (n_7144, n7474);
  and g12894 (n7476, n7438, n_7144);
  not g12895 (n_7145, n7475);
  not g12896 (n_7146, n7476);
  and g12897 (n7477, n_7145, n_7146);
  not g12898 (n_7148, \A[157] );
  and g12899 (n7478, n_7148, \A[158] );
  not g12900 (n_7150, \A[158] );
  and g12901 (n7479, \A[157] , n_7150);
  not g12902 (n_7152, n7479);
  and g12903 (n7480, \A[159] , n_7152);
  not g12904 (n_7153, n7478);
  and g12905 (n7481, n_7153, n7480);
  and g12906 (n7482, n_7153, n_7152);
  not g12907 (n_7154, \A[159] );
  not g12908 (n_7155, n7482);
  and g12909 (n7483, n_7154, n_7155);
  not g12910 (n_7156, n7481);
  not g12911 (n_7157, n7483);
  and g12912 (n7484, n_7156, n_7157);
  not g12913 (n_7159, \A[160] );
  and g12914 (n7485, n_7159, \A[161] );
  not g12915 (n_7161, \A[161] );
  and g12916 (n7486, \A[160] , n_7161);
  not g12917 (n_7163, n7486);
  and g12918 (n7487, \A[162] , n_7163);
  not g12919 (n_7164, n7485);
  and g12920 (n7488, n_7164, n7487);
  and g12921 (n7489, n_7164, n_7163);
  not g12922 (n_7165, \A[162] );
  not g12923 (n_7166, n7489);
  and g12924 (n7490, n_7165, n_7166);
  not g12925 (n_7167, n7488);
  not g12926 (n_7168, n7490);
  and g12927 (n7491, n_7167, n_7168);
  not g12928 (n_7169, n7484);
  and g12929 (n7492, n_7169, n7491);
  not g12930 (n_7170, n7491);
  and g12931 (n7493, n7484, n_7170);
  not g12932 (n_7171, n7492);
  not g12933 (n_7172, n7493);
  and g12934 (n7494, n_7171, n_7172);
  and g12935 (n7495, \A[160] , \A[161] );
  and g12936 (n7496, \A[162] , n_7166);
  not g12937 (n_7173, n7495);
  not g12938 (n_7174, n7496);
  and g12939 (n7497, n_7173, n_7174);
  and g12940 (n7498, \A[157] , \A[158] );
  and g12941 (n7499, \A[159] , n_7155);
  not g12942 (n_7175, n7498);
  not g12943 (n_7176, n7499);
  and g12944 (n7500, n_7175, n_7176);
  not g12945 (n_7177, n7497);
  and g12946 (n7501, n_7177, n7500);
  not g12947 (n_7178, n7500);
  and g12948 (n7502, n7497, n_7178);
  not g12949 (n_7179, n7501);
  not g12950 (n_7180, n7502);
  and g12951 (n7503, n_7179, n_7180);
  and g12952 (n7504, n_7169, n_7170);
  not g12953 (n_7181, n7503);
  and g12954 (n7505, n_7181, n7504);
  and g12955 (n7506, n_7177, n_7178);
  not g12956 (n_7182, n7505);
  not g12957 (n_7183, n7506);
  and g12958 (n7507, n_7182, n_7183);
  and g12959 (n7508, n_7179, n7504);
  and g12960 (n7509, n_7180, n7508);
  not g12961 (n_7184, n7504);
  and g12962 (n7510, n_7181, n_7184);
  not g12963 (n_7185, n7509);
  not g12964 (n_7186, n7510);
  and g12965 (n7511, n_7185, n_7186);
  not g12966 (n_7187, n7507);
  not g12967 (n_7188, n7511);
  and g12968 (n7512, n_7187, n_7188);
  not g12969 (n_7189, n7494);
  not g12970 (n_7190, n7512);
  and g12971 (n7513, n_7189, n_7190);
  not g12972 (n_7192, \A[151] );
  and g12973 (n7514, n_7192, \A[152] );
  not g12974 (n_7194, \A[152] );
  and g12975 (n7515, \A[151] , n_7194);
  not g12976 (n_7196, n7515);
  and g12977 (n7516, \A[153] , n_7196);
  not g12978 (n_7197, n7514);
  and g12979 (n7517, n_7197, n7516);
  and g12980 (n7518, n_7197, n_7196);
  not g12981 (n_7198, \A[153] );
  not g12982 (n_7199, n7518);
  and g12983 (n7519, n_7198, n_7199);
  not g12984 (n_7200, n7517);
  not g12985 (n_7201, n7519);
  and g12986 (n7520, n_7200, n_7201);
  not g12987 (n_7203, \A[154] );
  and g12988 (n7521, n_7203, \A[155] );
  not g12989 (n_7205, \A[155] );
  and g12990 (n7522, \A[154] , n_7205);
  not g12991 (n_7207, n7522);
  and g12992 (n7523, \A[156] , n_7207);
  not g12993 (n_7208, n7521);
  and g12994 (n7524, n_7208, n7523);
  and g12995 (n7525, n_7208, n_7207);
  not g12996 (n_7209, \A[156] );
  not g12997 (n_7210, n7525);
  and g12998 (n7526, n_7209, n_7210);
  not g12999 (n_7211, n7524);
  not g13000 (n_7212, n7526);
  and g13001 (n7527, n_7211, n_7212);
  not g13002 (n_7213, n7520);
  and g13003 (n7528, n_7213, n7527);
  not g13004 (n_7214, n7527);
  and g13005 (n7529, n7520, n_7214);
  not g13006 (n_7215, n7528);
  not g13007 (n_7216, n7529);
  and g13008 (n7530, n_7215, n_7216);
  and g13009 (n7531, \A[154] , \A[155] );
  and g13010 (n7532, \A[156] , n_7210);
  not g13011 (n_7217, n7531);
  not g13012 (n_7218, n7532);
  and g13013 (n7533, n_7217, n_7218);
  and g13014 (n7534, \A[151] , \A[152] );
  and g13015 (n7535, \A[153] , n_7199);
  not g13016 (n_7219, n7534);
  not g13017 (n_7220, n7535);
  and g13018 (n7536, n_7219, n_7220);
  not g13019 (n_7221, n7533);
  and g13020 (n7537, n_7221, n7536);
  not g13021 (n_7222, n7536);
  and g13022 (n7538, n7533, n_7222);
  not g13023 (n_7223, n7537);
  not g13024 (n_7224, n7538);
  and g13025 (n7539, n_7223, n_7224);
  and g13026 (n7540, n_7213, n_7214);
  not g13027 (n_7225, n7539);
  and g13028 (n7541, n_7225, n7540);
  and g13029 (n7542, n_7221, n_7222);
  not g13030 (n_7226, n7541);
  not g13031 (n_7227, n7542);
  and g13032 (n7543, n_7226, n_7227);
  and g13033 (n7544, n_7223, n7540);
  and g13034 (n7545, n_7224, n7544);
  not g13035 (n_7228, n7540);
  and g13036 (n7546, n_7225, n_7228);
  not g13037 (n_7229, n7545);
  not g13038 (n_7230, n7546);
  and g13039 (n7547, n_7229, n_7230);
  not g13040 (n_7231, n7543);
  not g13041 (n_7232, n7547);
  and g13042 (n7548, n_7231, n_7232);
  not g13043 (n_7233, n7530);
  not g13044 (n_7234, n7548);
  and g13045 (n7549, n_7233, n_7234);
  not g13046 (n_7235, n7513);
  and g13047 (n7550, n_7235, n7549);
  not g13048 (n_7236, n7549);
  and g13049 (n7551, n7513, n_7236);
  not g13050 (n_7237, n7550);
  not g13051 (n_7238, n7551);
  and g13052 (n7552, n_7237, n_7238);
  not g13053 (n_7239, n7477);
  and g13054 (n7553, n_7239, n7552);
  not g13055 (n_7240, n7552);
  and g13056 (n7554, n7477, n_7240);
  not g13057 (n_7241, n7553);
  not g13058 (n_7242, n7554);
  and g13059 (n7555, n_7241, n_7242);
  not g13060 (n_7244, \A[145] );
  and g13061 (n7556, n_7244, \A[146] );
  not g13062 (n_7246, \A[146] );
  and g13063 (n7557, \A[145] , n_7246);
  not g13064 (n_7248, n7557);
  and g13065 (n7558, \A[147] , n_7248);
  not g13066 (n_7249, n7556);
  and g13067 (n7559, n_7249, n7558);
  and g13068 (n7560, n_7249, n_7248);
  not g13069 (n_7250, \A[147] );
  not g13070 (n_7251, n7560);
  and g13071 (n7561, n_7250, n_7251);
  not g13072 (n_7252, n7559);
  not g13073 (n_7253, n7561);
  and g13074 (n7562, n_7252, n_7253);
  not g13075 (n_7255, \A[148] );
  and g13076 (n7563, n_7255, \A[149] );
  not g13077 (n_7257, \A[149] );
  and g13078 (n7564, \A[148] , n_7257);
  not g13079 (n_7259, n7564);
  and g13080 (n7565, \A[150] , n_7259);
  not g13081 (n_7260, n7563);
  and g13082 (n7566, n_7260, n7565);
  and g13083 (n7567, n_7260, n_7259);
  not g13084 (n_7261, \A[150] );
  not g13085 (n_7262, n7567);
  and g13086 (n7568, n_7261, n_7262);
  not g13087 (n_7263, n7566);
  not g13088 (n_7264, n7568);
  and g13089 (n7569, n_7263, n_7264);
  not g13090 (n_7265, n7562);
  and g13091 (n7570, n_7265, n7569);
  not g13092 (n_7266, n7569);
  and g13093 (n7571, n7562, n_7266);
  not g13094 (n_7267, n7570);
  not g13095 (n_7268, n7571);
  and g13096 (n7572, n_7267, n_7268);
  and g13097 (n7573, \A[148] , \A[149] );
  and g13098 (n7574, \A[150] , n_7262);
  not g13099 (n_7269, n7573);
  not g13100 (n_7270, n7574);
  and g13101 (n7575, n_7269, n_7270);
  and g13102 (n7576, \A[145] , \A[146] );
  and g13103 (n7577, \A[147] , n_7251);
  not g13104 (n_7271, n7576);
  not g13105 (n_7272, n7577);
  and g13106 (n7578, n_7271, n_7272);
  not g13107 (n_7273, n7575);
  and g13108 (n7579, n_7273, n7578);
  not g13109 (n_7274, n7578);
  and g13110 (n7580, n7575, n_7274);
  not g13111 (n_7275, n7579);
  not g13112 (n_7276, n7580);
  and g13113 (n7581, n_7275, n_7276);
  and g13114 (n7582, n_7265, n_7266);
  not g13115 (n_7277, n7581);
  and g13116 (n7583, n_7277, n7582);
  and g13117 (n7584, n_7273, n_7274);
  not g13118 (n_7278, n7583);
  not g13119 (n_7279, n7584);
  and g13120 (n7585, n_7278, n_7279);
  and g13121 (n7586, n_7275, n7582);
  and g13122 (n7587, n_7276, n7586);
  not g13123 (n_7280, n7582);
  and g13124 (n7588, n_7277, n_7280);
  not g13125 (n_7281, n7587);
  not g13126 (n_7282, n7588);
  and g13127 (n7589, n_7281, n_7282);
  not g13128 (n_7283, n7585);
  not g13129 (n_7284, n7589);
  and g13130 (n7590, n_7283, n_7284);
  not g13131 (n_7285, n7572);
  not g13132 (n_7286, n7590);
  and g13133 (n7591, n_7285, n_7286);
  not g13134 (n_7288, \A[139] );
  and g13135 (n7592, n_7288, \A[140] );
  not g13136 (n_7290, \A[140] );
  and g13137 (n7593, \A[139] , n_7290);
  not g13138 (n_7292, n7593);
  and g13139 (n7594, \A[141] , n_7292);
  not g13140 (n_7293, n7592);
  and g13141 (n7595, n_7293, n7594);
  and g13142 (n7596, n_7293, n_7292);
  not g13143 (n_7294, \A[141] );
  not g13144 (n_7295, n7596);
  and g13145 (n7597, n_7294, n_7295);
  not g13146 (n_7296, n7595);
  not g13147 (n_7297, n7597);
  and g13148 (n7598, n_7296, n_7297);
  not g13149 (n_7299, \A[142] );
  and g13150 (n7599, n_7299, \A[143] );
  not g13151 (n_7301, \A[143] );
  and g13152 (n7600, \A[142] , n_7301);
  not g13153 (n_7303, n7600);
  and g13154 (n7601, \A[144] , n_7303);
  not g13155 (n_7304, n7599);
  and g13156 (n7602, n_7304, n7601);
  and g13157 (n7603, n_7304, n_7303);
  not g13158 (n_7305, \A[144] );
  not g13159 (n_7306, n7603);
  and g13160 (n7604, n_7305, n_7306);
  not g13161 (n_7307, n7602);
  not g13162 (n_7308, n7604);
  and g13163 (n7605, n_7307, n_7308);
  not g13164 (n_7309, n7598);
  and g13165 (n7606, n_7309, n7605);
  not g13166 (n_7310, n7605);
  and g13167 (n7607, n7598, n_7310);
  not g13168 (n_7311, n7606);
  not g13169 (n_7312, n7607);
  and g13170 (n7608, n_7311, n_7312);
  and g13171 (n7609, \A[142] , \A[143] );
  and g13172 (n7610, \A[144] , n_7306);
  not g13173 (n_7313, n7609);
  not g13174 (n_7314, n7610);
  and g13175 (n7611, n_7313, n_7314);
  and g13176 (n7612, \A[139] , \A[140] );
  and g13177 (n7613, \A[141] , n_7295);
  not g13178 (n_7315, n7612);
  not g13179 (n_7316, n7613);
  and g13180 (n7614, n_7315, n_7316);
  not g13181 (n_7317, n7611);
  and g13182 (n7615, n_7317, n7614);
  not g13183 (n_7318, n7614);
  and g13184 (n7616, n7611, n_7318);
  not g13185 (n_7319, n7615);
  not g13186 (n_7320, n7616);
  and g13187 (n7617, n_7319, n_7320);
  and g13188 (n7618, n_7309, n_7310);
  not g13189 (n_7321, n7617);
  and g13190 (n7619, n_7321, n7618);
  and g13191 (n7620, n_7317, n_7318);
  not g13192 (n_7322, n7619);
  not g13193 (n_7323, n7620);
  and g13194 (n7621, n_7322, n_7323);
  and g13195 (n7622, n_7319, n7618);
  and g13196 (n7623, n_7320, n7622);
  not g13197 (n_7324, n7618);
  and g13198 (n7624, n_7321, n_7324);
  not g13199 (n_7325, n7623);
  not g13200 (n_7326, n7624);
  and g13201 (n7625, n_7325, n_7326);
  not g13202 (n_7327, n7621);
  not g13203 (n_7328, n7625);
  and g13204 (n7626, n_7327, n_7328);
  not g13205 (n_7329, n7608);
  not g13206 (n_7330, n7626);
  and g13207 (n7627, n_7329, n_7330);
  not g13208 (n_7331, n7591);
  and g13209 (n7628, n_7331, n7627);
  not g13210 (n_7332, n7627);
  and g13211 (n7629, n7591, n_7332);
  not g13212 (n_7333, n7628);
  not g13213 (n_7334, n7629);
  and g13214 (n7630, n_7333, n_7334);
  not g13215 (n_7336, \A[133] );
  and g13216 (n7631, n_7336, \A[134] );
  not g13217 (n_7338, \A[134] );
  and g13218 (n7632, \A[133] , n_7338);
  not g13219 (n_7340, n7632);
  and g13220 (n7633, \A[135] , n_7340);
  not g13221 (n_7341, n7631);
  and g13222 (n7634, n_7341, n7633);
  and g13223 (n7635, n_7341, n_7340);
  not g13224 (n_7342, \A[135] );
  not g13225 (n_7343, n7635);
  and g13226 (n7636, n_7342, n_7343);
  not g13227 (n_7344, n7634);
  not g13228 (n_7345, n7636);
  and g13229 (n7637, n_7344, n_7345);
  not g13230 (n_7347, \A[136] );
  and g13231 (n7638, n_7347, \A[137] );
  not g13232 (n_7349, \A[137] );
  and g13233 (n7639, \A[136] , n_7349);
  not g13234 (n_7351, n7639);
  and g13235 (n7640, \A[138] , n_7351);
  not g13236 (n_7352, n7638);
  and g13237 (n7641, n_7352, n7640);
  and g13238 (n7642, n_7352, n_7351);
  not g13239 (n_7353, \A[138] );
  not g13240 (n_7354, n7642);
  and g13241 (n7643, n_7353, n_7354);
  not g13242 (n_7355, n7641);
  not g13243 (n_7356, n7643);
  and g13244 (n7644, n_7355, n_7356);
  not g13245 (n_7357, n7637);
  and g13246 (n7645, n_7357, n7644);
  not g13247 (n_7358, n7644);
  and g13248 (n7646, n7637, n_7358);
  not g13249 (n_7359, n7645);
  not g13250 (n_7360, n7646);
  and g13251 (n7647, n_7359, n_7360);
  and g13252 (n7648, \A[136] , \A[137] );
  and g13253 (n7649, \A[138] , n_7354);
  not g13254 (n_7361, n7648);
  not g13255 (n_7362, n7649);
  and g13256 (n7650, n_7361, n_7362);
  and g13257 (n7651, \A[133] , \A[134] );
  and g13258 (n7652, \A[135] , n_7343);
  not g13259 (n_7363, n7651);
  not g13260 (n_7364, n7652);
  and g13261 (n7653, n_7363, n_7364);
  not g13262 (n_7365, n7650);
  and g13263 (n7654, n_7365, n7653);
  not g13264 (n_7366, n7653);
  and g13265 (n7655, n7650, n_7366);
  not g13266 (n_7367, n7654);
  not g13267 (n_7368, n7655);
  and g13268 (n7656, n_7367, n_7368);
  and g13269 (n7657, n_7357, n_7358);
  not g13270 (n_7369, n7656);
  and g13271 (n7658, n_7369, n7657);
  and g13272 (n7659, n_7365, n_7366);
  not g13273 (n_7370, n7658);
  not g13274 (n_7371, n7659);
  and g13275 (n7660, n_7370, n_7371);
  and g13276 (n7661, n_7367, n7657);
  and g13277 (n7662, n_7368, n7661);
  not g13278 (n_7372, n7657);
  and g13279 (n7663, n_7369, n_7372);
  not g13280 (n_7373, n7662);
  not g13281 (n_7374, n7663);
  and g13282 (n7664, n_7373, n_7374);
  not g13283 (n_7375, n7660);
  not g13284 (n_7376, n7664);
  and g13285 (n7665, n_7375, n_7376);
  not g13286 (n_7377, n7647);
  not g13287 (n_7378, n7665);
  and g13288 (n7666, n_7377, n_7378);
  not g13289 (n_7380, \A[127] );
  and g13290 (n7667, n_7380, \A[128] );
  not g13291 (n_7382, \A[128] );
  and g13292 (n7668, \A[127] , n_7382);
  not g13293 (n_7384, n7668);
  and g13294 (n7669, \A[129] , n_7384);
  not g13295 (n_7385, n7667);
  and g13296 (n7670, n_7385, n7669);
  and g13297 (n7671, n_7385, n_7384);
  not g13298 (n_7386, \A[129] );
  not g13299 (n_7387, n7671);
  and g13300 (n7672, n_7386, n_7387);
  not g13301 (n_7388, n7670);
  not g13302 (n_7389, n7672);
  and g13303 (n7673, n_7388, n_7389);
  not g13304 (n_7391, \A[130] );
  and g13305 (n7674, n_7391, \A[131] );
  not g13306 (n_7393, \A[131] );
  and g13307 (n7675, \A[130] , n_7393);
  not g13308 (n_7395, n7675);
  and g13309 (n7676, \A[132] , n_7395);
  not g13310 (n_7396, n7674);
  and g13311 (n7677, n_7396, n7676);
  and g13312 (n7678, n_7396, n_7395);
  not g13313 (n_7397, \A[132] );
  not g13314 (n_7398, n7678);
  and g13315 (n7679, n_7397, n_7398);
  not g13316 (n_7399, n7677);
  not g13317 (n_7400, n7679);
  and g13318 (n7680, n_7399, n_7400);
  not g13319 (n_7401, n7673);
  and g13320 (n7681, n_7401, n7680);
  not g13321 (n_7402, n7680);
  and g13322 (n7682, n7673, n_7402);
  not g13323 (n_7403, n7681);
  not g13324 (n_7404, n7682);
  and g13325 (n7683, n_7403, n_7404);
  and g13326 (n7684, \A[130] , \A[131] );
  and g13327 (n7685, \A[132] , n_7398);
  not g13328 (n_7405, n7684);
  not g13329 (n_7406, n7685);
  and g13330 (n7686, n_7405, n_7406);
  and g13331 (n7687, \A[127] , \A[128] );
  and g13332 (n7688, \A[129] , n_7387);
  not g13333 (n_7407, n7687);
  not g13334 (n_7408, n7688);
  and g13335 (n7689, n_7407, n_7408);
  not g13336 (n_7409, n7686);
  and g13337 (n7690, n_7409, n7689);
  not g13338 (n_7410, n7689);
  and g13339 (n7691, n7686, n_7410);
  not g13340 (n_7411, n7690);
  not g13341 (n_7412, n7691);
  and g13342 (n7692, n_7411, n_7412);
  and g13343 (n7693, n_7401, n_7402);
  not g13344 (n_7413, n7692);
  and g13345 (n7694, n_7413, n7693);
  and g13346 (n7695, n_7409, n_7410);
  not g13347 (n_7414, n7694);
  not g13348 (n_7415, n7695);
  and g13349 (n7696, n_7414, n_7415);
  and g13350 (n7697, n_7411, n7693);
  and g13351 (n7698, n_7412, n7697);
  not g13352 (n_7416, n7693);
  and g13353 (n7699, n_7413, n_7416);
  not g13354 (n_7417, n7698);
  not g13355 (n_7418, n7699);
  and g13356 (n7700, n_7417, n_7418);
  not g13357 (n_7419, n7696);
  not g13358 (n_7420, n7700);
  and g13359 (n7701, n_7419, n_7420);
  not g13360 (n_7421, n7683);
  not g13361 (n_7422, n7701);
  and g13362 (n7702, n_7421, n_7422);
  not g13363 (n_7423, n7666);
  and g13364 (n7703, n_7423, n7702);
  not g13365 (n_7424, n7702);
  and g13366 (n7704, n7666, n_7424);
  not g13367 (n_7425, n7703);
  not g13368 (n_7426, n7704);
  and g13369 (n7705, n_7425, n_7426);
  not g13370 (n_7427, n7630);
  and g13371 (n7706, n_7427, n7705);
  not g13372 (n_7428, n7705);
  and g13373 (n7707, n7630, n_7428);
  not g13374 (n_7429, n7706);
  not g13375 (n_7430, n7707);
  and g13376 (n7708, n_7429, n_7430);
  not g13377 (n_7431, n7555);
  and g13378 (n7709, n_7431, n7708);
  not g13379 (n_7432, n7708);
  and g13380 (n7710, n7555, n_7432);
  not g13381 (n_7433, n7709);
  not g13382 (n_7434, n7710);
  and g13383 (n7711, n_7433, n_7434);
  not g13384 (n_7436, \A[121] );
  and g13385 (n7712, n_7436, \A[122] );
  not g13386 (n_7438, \A[122] );
  and g13387 (n7713, \A[121] , n_7438);
  not g13388 (n_7440, n7713);
  and g13389 (n7714, \A[123] , n_7440);
  not g13390 (n_7441, n7712);
  and g13391 (n7715, n_7441, n7714);
  and g13392 (n7716, n_7441, n_7440);
  not g13393 (n_7442, \A[123] );
  not g13394 (n_7443, n7716);
  and g13395 (n7717, n_7442, n_7443);
  not g13396 (n_7444, n7715);
  not g13397 (n_7445, n7717);
  and g13398 (n7718, n_7444, n_7445);
  not g13399 (n_7447, \A[124] );
  and g13400 (n7719, n_7447, \A[125] );
  not g13401 (n_7449, \A[125] );
  and g13402 (n7720, \A[124] , n_7449);
  not g13403 (n_7451, n7720);
  and g13404 (n7721, \A[126] , n_7451);
  not g13405 (n_7452, n7719);
  and g13406 (n7722, n_7452, n7721);
  and g13407 (n7723, n_7452, n_7451);
  not g13408 (n_7453, \A[126] );
  not g13409 (n_7454, n7723);
  and g13410 (n7724, n_7453, n_7454);
  not g13411 (n_7455, n7722);
  not g13412 (n_7456, n7724);
  and g13413 (n7725, n_7455, n_7456);
  not g13414 (n_7457, n7718);
  and g13415 (n7726, n_7457, n7725);
  not g13416 (n_7458, n7725);
  and g13417 (n7727, n7718, n_7458);
  not g13418 (n_7459, n7726);
  not g13419 (n_7460, n7727);
  and g13420 (n7728, n_7459, n_7460);
  and g13421 (n7729, \A[124] , \A[125] );
  and g13422 (n7730, \A[126] , n_7454);
  not g13423 (n_7461, n7729);
  not g13424 (n_7462, n7730);
  and g13425 (n7731, n_7461, n_7462);
  and g13426 (n7732, \A[121] , \A[122] );
  and g13427 (n7733, \A[123] , n_7443);
  not g13428 (n_7463, n7732);
  not g13429 (n_7464, n7733);
  and g13430 (n7734, n_7463, n_7464);
  not g13431 (n_7465, n7731);
  and g13432 (n7735, n_7465, n7734);
  not g13433 (n_7466, n7734);
  and g13434 (n7736, n7731, n_7466);
  not g13435 (n_7467, n7735);
  not g13436 (n_7468, n7736);
  and g13437 (n7737, n_7467, n_7468);
  and g13438 (n7738, n_7457, n_7458);
  not g13439 (n_7469, n7737);
  and g13440 (n7739, n_7469, n7738);
  and g13441 (n7740, n_7465, n_7466);
  not g13442 (n_7470, n7739);
  not g13443 (n_7471, n7740);
  and g13444 (n7741, n_7470, n_7471);
  and g13445 (n7742, n_7467, n7738);
  and g13446 (n7743, n_7468, n7742);
  not g13447 (n_7472, n7738);
  and g13448 (n7744, n_7469, n_7472);
  not g13449 (n_7473, n7743);
  not g13450 (n_7474, n7744);
  and g13451 (n7745, n_7473, n_7474);
  not g13452 (n_7475, n7741);
  not g13453 (n_7476, n7745);
  and g13454 (n7746, n_7475, n_7476);
  not g13455 (n_7477, n7728);
  not g13456 (n_7478, n7746);
  and g13457 (n7747, n_7477, n_7478);
  not g13458 (n_7480, \A[115] );
  and g13459 (n7748, n_7480, \A[116] );
  not g13460 (n_7482, \A[116] );
  and g13461 (n7749, \A[115] , n_7482);
  not g13462 (n_7484, n7749);
  and g13463 (n7750, \A[117] , n_7484);
  not g13464 (n_7485, n7748);
  and g13465 (n7751, n_7485, n7750);
  and g13466 (n7752, n_7485, n_7484);
  not g13467 (n_7486, \A[117] );
  not g13468 (n_7487, n7752);
  and g13469 (n7753, n_7486, n_7487);
  not g13470 (n_7488, n7751);
  not g13471 (n_7489, n7753);
  and g13472 (n7754, n_7488, n_7489);
  not g13473 (n_7491, \A[118] );
  and g13474 (n7755, n_7491, \A[119] );
  not g13475 (n_7493, \A[119] );
  and g13476 (n7756, \A[118] , n_7493);
  not g13477 (n_7495, n7756);
  and g13478 (n7757, \A[120] , n_7495);
  not g13479 (n_7496, n7755);
  and g13480 (n7758, n_7496, n7757);
  and g13481 (n7759, n_7496, n_7495);
  not g13482 (n_7497, \A[120] );
  not g13483 (n_7498, n7759);
  and g13484 (n7760, n_7497, n_7498);
  not g13485 (n_7499, n7758);
  not g13486 (n_7500, n7760);
  and g13487 (n7761, n_7499, n_7500);
  not g13488 (n_7501, n7754);
  and g13489 (n7762, n_7501, n7761);
  not g13490 (n_7502, n7761);
  and g13491 (n7763, n7754, n_7502);
  not g13492 (n_7503, n7762);
  not g13493 (n_7504, n7763);
  and g13494 (n7764, n_7503, n_7504);
  and g13495 (n7765, \A[118] , \A[119] );
  and g13496 (n7766, \A[120] , n_7498);
  not g13497 (n_7505, n7765);
  not g13498 (n_7506, n7766);
  and g13499 (n7767, n_7505, n_7506);
  and g13500 (n7768, \A[115] , \A[116] );
  and g13501 (n7769, \A[117] , n_7487);
  not g13502 (n_7507, n7768);
  not g13503 (n_7508, n7769);
  and g13504 (n7770, n_7507, n_7508);
  not g13505 (n_7509, n7767);
  and g13506 (n7771, n_7509, n7770);
  not g13507 (n_7510, n7770);
  and g13508 (n7772, n7767, n_7510);
  not g13509 (n_7511, n7771);
  not g13510 (n_7512, n7772);
  and g13511 (n7773, n_7511, n_7512);
  and g13512 (n7774, n_7501, n_7502);
  not g13513 (n_7513, n7773);
  and g13514 (n7775, n_7513, n7774);
  and g13515 (n7776, n_7509, n_7510);
  not g13516 (n_7514, n7775);
  not g13517 (n_7515, n7776);
  and g13518 (n7777, n_7514, n_7515);
  and g13519 (n7778, n_7511, n7774);
  and g13520 (n7779, n_7512, n7778);
  not g13521 (n_7516, n7774);
  and g13522 (n7780, n_7513, n_7516);
  not g13523 (n_7517, n7779);
  not g13524 (n_7518, n7780);
  and g13525 (n7781, n_7517, n_7518);
  not g13526 (n_7519, n7777);
  not g13527 (n_7520, n7781);
  and g13528 (n7782, n_7519, n_7520);
  not g13529 (n_7521, n7764);
  not g13530 (n_7522, n7782);
  and g13531 (n7783, n_7521, n_7522);
  not g13532 (n_7523, n7747);
  and g13533 (n7784, n_7523, n7783);
  not g13534 (n_7524, n7783);
  and g13535 (n7785, n7747, n_7524);
  not g13536 (n_7525, n7784);
  not g13537 (n_7526, n7785);
  and g13538 (n7786, n_7525, n_7526);
  not g13539 (n_7528, \A[109] );
  and g13540 (n7787, n_7528, \A[110] );
  not g13541 (n_7530, \A[110] );
  and g13542 (n7788, \A[109] , n_7530);
  not g13543 (n_7532, n7788);
  and g13544 (n7789, \A[111] , n_7532);
  not g13545 (n_7533, n7787);
  and g13546 (n7790, n_7533, n7789);
  and g13547 (n7791, n_7533, n_7532);
  not g13548 (n_7534, \A[111] );
  not g13549 (n_7535, n7791);
  and g13550 (n7792, n_7534, n_7535);
  not g13551 (n_7536, n7790);
  not g13552 (n_7537, n7792);
  and g13553 (n7793, n_7536, n_7537);
  not g13554 (n_7539, \A[112] );
  and g13555 (n7794, n_7539, \A[113] );
  not g13556 (n_7541, \A[113] );
  and g13557 (n7795, \A[112] , n_7541);
  not g13558 (n_7543, n7795);
  and g13559 (n7796, \A[114] , n_7543);
  not g13560 (n_7544, n7794);
  and g13561 (n7797, n_7544, n7796);
  and g13562 (n7798, n_7544, n_7543);
  not g13563 (n_7545, \A[114] );
  not g13564 (n_7546, n7798);
  and g13565 (n7799, n_7545, n_7546);
  not g13566 (n_7547, n7797);
  not g13567 (n_7548, n7799);
  and g13568 (n7800, n_7547, n_7548);
  not g13569 (n_7549, n7793);
  and g13570 (n7801, n_7549, n7800);
  not g13571 (n_7550, n7800);
  and g13572 (n7802, n7793, n_7550);
  not g13573 (n_7551, n7801);
  not g13574 (n_7552, n7802);
  and g13575 (n7803, n_7551, n_7552);
  and g13576 (n7804, \A[112] , \A[113] );
  and g13577 (n7805, \A[114] , n_7546);
  not g13578 (n_7553, n7804);
  not g13579 (n_7554, n7805);
  and g13580 (n7806, n_7553, n_7554);
  and g13581 (n7807, \A[109] , \A[110] );
  and g13582 (n7808, \A[111] , n_7535);
  not g13583 (n_7555, n7807);
  not g13584 (n_7556, n7808);
  and g13585 (n7809, n_7555, n_7556);
  not g13586 (n_7557, n7806);
  and g13587 (n7810, n_7557, n7809);
  not g13588 (n_7558, n7809);
  and g13589 (n7811, n7806, n_7558);
  not g13590 (n_7559, n7810);
  not g13591 (n_7560, n7811);
  and g13592 (n7812, n_7559, n_7560);
  and g13593 (n7813, n_7549, n_7550);
  not g13594 (n_7561, n7812);
  and g13595 (n7814, n_7561, n7813);
  and g13596 (n7815, n_7557, n_7558);
  not g13597 (n_7562, n7814);
  not g13598 (n_7563, n7815);
  and g13599 (n7816, n_7562, n_7563);
  and g13600 (n7817, n_7559, n7813);
  and g13601 (n7818, n_7560, n7817);
  not g13602 (n_7564, n7813);
  and g13603 (n7819, n_7561, n_7564);
  not g13604 (n_7565, n7818);
  not g13605 (n_7566, n7819);
  and g13606 (n7820, n_7565, n_7566);
  not g13607 (n_7567, n7816);
  not g13608 (n_7568, n7820);
  and g13609 (n7821, n_7567, n_7568);
  not g13610 (n_7569, n7803);
  not g13611 (n_7570, n7821);
  and g13612 (n7822, n_7569, n_7570);
  not g13613 (n_7572, \A[103] );
  and g13614 (n7823, n_7572, \A[104] );
  not g13615 (n_7574, \A[104] );
  and g13616 (n7824, \A[103] , n_7574);
  not g13617 (n_7576, n7824);
  and g13618 (n7825, \A[105] , n_7576);
  not g13619 (n_7577, n7823);
  and g13620 (n7826, n_7577, n7825);
  and g13621 (n7827, n_7577, n_7576);
  not g13622 (n_7578, \A[105] );
  not g13623 (n_7579, n7827);
  and g13624 (n7828, n_7578, n_7579);
  not g13625 (n_7580, n7826);
  not g13626 (n_7581, n7828);
  and g13627 (n7829, n_7580, n_7581);
  not g13628 (n_7583, \A[106] );
  and g13629 (n7830, n_7583, \A[107] );
  not g13630 (n_7585, \A[107] );
  and g13631 (n7831, \A[106] , n_7585);
  not g13632 (n_7587, n7831);
  and g13633 (n7832, \A[108] , n_7587);
  not g13634 (n_7588, n7830);
  and g13635 (n7833, n_7588, n7832);
  and g13636 (n7834, n_7588, n_7587);
  not g13637 (n_7589, \A[108] );
  not g13638 (n_7590, n7834);
  and g13639 (n7835, n_7589, n_7590);
  not g13640 (n_7591, n7833);
  not g13641 (n_7592, n7835);
  and g13642 (n7836, n_7591, n_7592);
  not g13643 (n_7593, n7829);
  and g13644 (n7837, n_7593, n7836);
  not g13645 (n_7594, n7836);
  and g13646 (n7838, n7829, n_7594);
  not g13647 (n_7595, n7837);
  not g13648 (n_7596, n7838);
  and g13649 (n7839, n_7595, n_7596);
  and g13650 (n7840, \A[106] , \A[107] );
  and g13651 (n7841, \A[108] , n_7590);
  not g13652 (n_7597, n7840);
  not g13653 (n_7598, n7841);
  and g13654 (n7842, n_7597, n_7598);
  and g13655 (n7843, \A[103] , \A[104] );
  and g13656 (n7844, \A[105] , n_7579);
  not g13657 (n_7599, n7843);
  not g13658 (n_7600, n7844);
  and g13659 (n7845, n_7599, n_7600);
  not g13660 (n_7601, n7842);
  and g13661 (n7846, n_7601, n7845);
  not g13662 (n_7602, n7845);
  and g13663 (n7847, n7842, n_7602);
  not g13664 (n_7603, n7846);
  not g13665 (n_7604, n7847);
  and g13666 (n7848, n_7603, n_7604);
  and g13667 (n7849, n_7593, n_7594);
  not g13668 (n_7605, n7848);
  and g13669 (n7850, n_7605, n7849);
  and g13670 (n7851, n_7601, n_7602);
  not g13671 (n_7606, n7850);
  not g13672 (n_7607, n7851);
  and g13673 (n7852, n_7606, n_7607);
  and g13674 (n7853, n_7603, n7849);
  and g13675 (n7854, n_7604, n7853);
  not g13676 (n_7608, n7849);
  and g13677 (n7855, n_7605, n_7608);
  not g13678 (n_7609, n7854);
  not g13679 (n_7610, n7855);
  and g13680 (n7856, n_7609, n_7610);
  not g13681 (n_7611, n7852);
  not g13682 (n_7612, n7856);
  and g13683 (n7857, n_7611, n_7612);
  not g13684 (n_7613, n7839);
  not g13685 (n_7614, n7857);
  and g13686 (n7858, n_7613, n_7614);
  not g13687 (n_7615, n7822);
  and g13688 (n7859, n_7615, n7858);
  not g13689 (n_7616, n7858);
  and g13690 (n7860, n7822, n_7616);
  not g13691 (n_7617, n7859);
  not g13692 (n_7618, n7860);
  and g13693 (n7861, n_7617, n_7618);
  not g13694 (n_7619, n7786);
  and g13695 (n7862, n_7619, n7861);
  not g13696 (n_7620, n7861);
  and g13697 (n7863, n7786, n_7620);
  not g13698 (n_7621, n7862);
  not g13699 (n_7622, n7863);
  and g13700 (n7864, n_7621, n_7622);
  not g13701 (n_7624, \A[97] );
  and g13702 (n7865, n_7624, \A[98] );
  not g13703 (n_7626, \A[98] );
  and g13704 (n7866, \A[97] , n_7626);
  not g13705 (n_7628, n7866);
  and g13706 (n7867, \A[99] , n_7628);
  not g13707 (n_7629, n7865);
  and g13708 (n7868, n_7629, n7867);
  and g13709 (n7869, n_7629, n_7628);
  not g13710 (n_7630, \A[99] );
  not g13711 (n_7631, n7869);
  and g13712 (n7870, n_7630, n_7631);
  not g13713 (n_7632, n7868);
  not g13714 (n_7633, n7870);
  and g13715 (n7871, n_7632, n_7633);
  not g13716 (n_7635, \A[100] );
  and g13717 (n7872, n_7635, \A[101] );
  not g13718 (n_7637, \A[101] );
  and g13719 (n7873, \A[100] , n_7637);
  not g13720 (n_7639, n7873);
  and g13721 (n7874, \A[102] , n_7639);
  not g13722 (n_7640, n7872);
  and g13723 (n7875, n_7640, n7874);
  and g13724 (n7876, n_7640, n_7639);
  not g13725 (n_7641, \A[102] );
  not g13726 (n_7642, n7876);
  and g13727 (n7877, n_7641, n_7642);
  not g13728 (n_7643, n7875);
  not g13729 (n_7644, n7877);
  and g13730 (n7878, n_7643, n_7644);
  not g13731 (n_7645, n7871);
  and g13732 (n7879, n_7645, n7878);
  not g13733 (n_7646, n7878);
  and g13734 (n7880, n7871, n_7646);
  not g13735 (n_7647, n7879);
  not g13736 (n_7648, n7880);
  and g13737 (n7881, n_7647, n_7648);
  and g13738 (n7882, \A[100] , \A[101] );
  and g13739 (n7883, \A[102] , n_7642);
  not g13740 (n_7649, n7882);
  not g13741 (n_7650, n7883);
  and g13742 (n7884, n_7649, n_7650);
  and g13743 (n7885, \A[97] , \A[98] );
  and g13744 (n7886, \A[99] , n_7631);
  not g13745 (n_7651, n7885);
  not g13746 (n_7652, n7886);
  and g13747 (n7887, n_7651, n_7652);
  not g13748 (n_7653, n7884);
  and g13749 (n7888, n_7653, n7887);
  not g13750 (n_7654, n7887);
  and g13751 (n7889, n7884, n_7654);
  not g13752 (n_7655, n7888);
  not g13753 (n_7656, n7889);
  and g13754 (n7890, n_7655, n_7656);
  and g13755 (n7891, n_7645, n_7646);
  not g13756 (n_7657, n7890);
  and g13757 (n7892, n_7657, n7891);
  and g13758 (n7893, n_7653, n_7654);
  not g13759 (n_7658, n7892);
  not g13760 (n_7659, n7893);
  and g13761 (n7894, n_7658, n_7659);
  and g13762 (n7895, n_7655, n7891);
  and g13763 (n7896, n_7656, n7895);
  not g13764 (n_7660, n7891);
  and g13765 (n7897, n_7657, n_7660);
  not g13766 (n_7661, n7896);
  not g13767 (n_7662, n7897);
  and g13768 (n7898, n_7661, n_7662);
  not g13769 (n_7663, n7894);
  not g13770 (n_7664, n7898);
  and g13771 (n7899, n_7663, n_7664);
  not g13772 (n_7665, n7881);
  not g13773 (n_7666, n7899);
  and g13774 (n7900, n_7665, n_7666);
  not g13775 (n_7668, \A[91] );
  and g13776 (n7901, n_7668, \A[92] );
  not g13777 (n_7670, \A[92] );
  and g13778 (n7902, \A[91] , n_7670);
  not g13779 (n_7672, n7902);
  and g13780 (n7903, \A[93] , n_7672);
  not g13781 (n_7673, n7901);
  and g13782 (n7904, n_7673, n7903);
  and g13783 (n7905, n_7673, n_7672);
  not g13784 (n_7674, \A[93] );
  not g13785 (n_7675, n7905);
  and g13786 (n7906, n_7674, n_7675);
  not g13787 (n_7676, n7904);
  not g13788 (n_7677, n7906);
  and g13789 (n7907, n_7676, n_7677);
  not g13790 (n_7679, \A[94] );
  and g13791 (n7908, n_7679, \A[95] );
  not g13792 (n_7681, \A[95] );
  and g13793 (n7909, \A[94] , n_7681);
  not g13794 (n_7683, n7909);
  and g13795 (n7910, \A[96] , n_7683);
  not g13796 (n_7684, n7908);
  and g13797 (n7911, n_7684, n7910);
  and g13798 (n7912, n_7684, n_7683);
  not g13799 (n_7685, \A[96] );
  not g13800 (n_7686, n7912);
  and g13801 (n7913, n_7685, n_7686);
  not g13802 (n_7687, n7911);
  not g13803 (n_7688, n7913);
  and g13804 (n7914, n_7687, n_7688);
  not g13805 (n_7689, n7907);
  and g13806 (n7915, n_7689, n7914);
  not g13807 (n_7690, n7914);
  and g13808 (n7916, n7907, n_7690);
  not g13809 (n_7691, n7915);
  not g13810 (n_7692, n7916);
  and g13811 (n7917, n_7691, n_7692);
  and g13812 (n7918, \A[94] , \A[95] );
  and g13813 (n7919, \A[96] , n_7686);
  not g13814 (n_7693, n7918);
  not g13815 (n_7694, n7919);
  and g13816 (n7920, n_7693, n_7694);
  and g13817 (n7921, \A[91] , \A[92] );
  and g13818 (n7922, \A[93] , n_7675);
  not g13819 (n_7695, n7921);
  not g13820 (n_7696, n7922);
  and g13821 (n7923, n_7695, n_7696);
  not g13822 (n_7697, n7920);
  and g13823 (n7924, n_7697, n7923);
  not g13824 (n_7698, n7923);
  and g13825 (n7925, n7920, n_7698);
  not g13826 (n_7699, n7924);
  not g13827 (n_7700, n7925);
  and g13828 (n7926, n_7699, n_7700);
  and g13829 (n7927, n_7689, n_7690);
  not g13830 (n_7701, n7926);
  and g13831 (n7928, n_7701, n7927);
  and g13832 (n7929, n_7697, n_7698);
  not g13833 (n_7702, n7928);
  not g13834 (n_7703, n7929);
  and g13835 (n7930, n_7702, n_7703);
  and g13836 (n7931, n_7699, n7927);
  and g13837 (n7932, n_7700, n7931);
  not g13838 (n_7704, n7927);
  and g13839 (n7933, n_7701, n_7704);
  not g13840 (n_7705, n7932);
  not g13841 (n_7706, n7933);
  and g13842 (n7934, n_7705, n_7706);
  not g13843 (n_7707, n7930);
  not g13844 (n_7708, n7934);
  and g13845 (n7935, n_7707, n_7708);
  not g13846 (n_7709, n7917);
  not g13847 (n_7710, n7935);
  and g13848 (n7936, n_7709, n_7710);
  not g13849 (n_7711, n7900);
  and g13850 (n7937, n_7711, n7936);
  not g13851 (n_7712, n7936);
  and g13852 (n7938, n7900, n_7712);
  not g13853 (n_7713, n7937);
  not g13854 (n_7714, n7938);
  and g13855 (n7939, n_7713, n_7714);
  not g13856 (n_7716, \A[85] );
  and g13857 (n7940, n_7716, \A[86] );
  not g13858 (n_7718, \A[86] );
  and g13859 (n7941, \A[85] , n_7718);
  not g13860 (n_7720, n7941);
  and g13861 (n7942, \A[87] , n_7720);
  not g13862 (n_7721, n7940);
  and g13863 (n7943, n_7721, n7942);
  and g13864 (n7944, n_7721, n_7720);
  not g13865 (n_7722, \A[87] );
  not g13866 (n_7723, n7944);
  and g13867 (n7945, n_7722, n_7723);
  not g13868 (n_7724, n7943);
  not g13869 (n_7725, n7945);
  and g13870 (n7946, n_7724, n_7725);
  not g13871 (n_7727, \A[88] );
  and g13872 (n7947, n_7727, \A[89] );
  not g13873 (n_7729, \A[89] );
  and g13874 (n7948, \A[88] , n_7729);
  not g13875 (n_7731, n7948);
  and g13876 (n7949, \A[90] , n_7731);
  not g13877 (n_7732, n7947);
  and g13878 (n7950, n_7732, n7949);
  and g13879 (n7951, n_7732, n_7731);
  not g13880 (n_7733, \A[90] );
  not g13881 (n_7734, n7951);
  and g13882 (n7952, n_7733, n_7734);
  not g13883 (n_7735, n7950);
  not g13884 (n_7736, n7952);
  and g13885 (n7953, n_7735, n_7736);
  not g13886 (n_7737, n7946);
  and g13887 (n7954, n_7737, n7953);
  not g13888 (n_7738, n7953);
  and g13889 (n7955, n7946, n_7738);
  not g13890 (n_7739, n7954);
  not g13891 (n_7740, n7955);
  and g13892 (n7956, n_7739, n_7740);
  and g13893 (n7957, \A[88] , \A[89] );
  and g13894 (n7958, \A[90] , n_7734);
  not g13895 (n_7741, n7957);
  not g13896 (n_7742, n7958);
  and g13897 (n7959, n_7741, n_7742);
  and g13898 (n7960, \A[85] , \A[86] );
  and g13899 (n7961, \A[87] , n_7723);
  not g13900 (n_7743, n7960);
  not g13901 (n_7744, n7961);
  and g13902 (n7962, n_7743, n_7744);
  not g13903 (n_7745, n7959);
  and g13904 (n7963, n_7745, n7962);
  not g13905 (n_7746, n7962);
  and g13906 (n7964, n7959, n_7746);
  not g13907 (n_7747, n7963);
  not g13908 (n_7748, n7964);
  and g13909 (n7965, n_7747, n_7748);
  and g13910 (n7966, n_7737, n_7738);
  not g13911 (n_7749, n7965);
  and g13912 (n7967, n_7749, n7966);
  and g13913 (n7968, n_7745, n_7746);
  not g13914 (n_7750, n7967);
  not g13915 (n_7751, n7968);
  and g13916 (n7969, n_7750, n_7751);
  and g13917 (n7970, n_7747, n7966);
  and g13918 (n7971, n_7748, n7970);
  not g13919 (n_7752, n7966);
  and g13920 (n7972, n_7749, n_7752);
  not g13921 (n_7753, n7971);
  not g13922 (n_7754, n7972);
  and g13923 (n7973, n_7753, n_7754);
  not g13924 (n_7755, n7969);
  not g13925 (n_7756, n7973);
  and g13926 (n7974, n_7755, n_7756);
  not g13927 (n_7757, n7956);
  not g13928 (n_7758, n7974);
  and g13929 (n7975, n_7757, n_7758);
  not g13930 (n_7760, \A[79] );
  and g13931 (n7976, n_7760, \A[80] );
  not g13932 (n_7762, \A[80] );
  and g13933 (n7977, \A[79] , n_7762);
  not g13934 (n_7764, n7977);
  and g13935 (n7978, \A[81] , n_7764);
  not g13936 (n_7765, n7976);
  and g13937 (n7979, n_7765, n7978);
  and g13938 (n7980, n_7765, n_7764);
  not g13939 (n_7766, \A[81] );
  not g13940 (n_7767, n7980);
  and g13941 (n7981, n_7766, n_7767);
  not g13942 (n_7768, n7979);
  not g13943 (n_7769, n7981);
  and g13944 (n7982, n_7768, n_7769);
  not g13945 (n_7771, \A[82] );
  and g13946 (n7983, n_7771, \A[83] );
  not g13947 (n_7773, \A[83] );
  and g13948 (n7984, \A[82] , n_7773);
  not g13949 (n_7775, n7984);
  and g13950 (n7985, \A[84] , n_7775);
  not g13951 (n_7776, n7983);
  and g13952 (n7986, n_7776, n7985);
  and g13953 (n7987, n_7776, n_7775);
  not g13954 (n_7777, \A[84] );
  not g13955 (n_7778, n7987);
  and g13956 (n7988, n_7777, n_7778);
  not g13957 (n_7779, n7986);
  not g13958 (n_7780, n7988);
  and g13959 (n7989, n_7779, n_7780);
  not g13960 (n_7781, n7982);
  and g13961 (n7990, n_7781, n7989);
  not g13962 (n_7782, n7989);
  and g13963 (n7991, n7982, n_7782);
  not g13964 (n_7783, n7990);
  not g13965 (n_7784, n7991);
  and g13966 (n7992, n_7783, n_7784);
  and g13967 (n7993, \A[82] , \A[83] );
  and g13968 (n7994, \A[84] , n_7778);
  not g13969 (n_7785, n7993);
  not g13970 (n_7786, n7994);
  and g13971 (n7995, n_7785, n_7786);
  and g13972 (n7996, \A[79] , \A[80] );
  and g13973 (n7997, \A[81] , n_7767);
  not g13974 (n_7787, n7996);
  not g13975 (n_7788, n7997);
  and g13976 (n7998, n_7787, n_7788);
  not g13977 (n_7789, n7995);
  and g13978 (n7999, n_7789, n7998);
  not g13979 (n_7790, n7998);
  and g13980 (n8000, n7995, n_7790);
  not g13981 (n_7791, n7999);
  not g13982 (n_7792, n8000);
  and g13983 (n8001, n_7791, n_7792);
  and g13984 (n8002, n_7781, n_7782);
  not g13985 (n_7793, n8001);
  and g13986 (n8003, n_7793, n8002);
  and g13987 (n8004, n_7789, n_7790);
  not g13988 (n_7794, n8003);
  not g13989 (n_7795, n8004);
  and g13990 (n8005, n_7794, n_7795);
  and g13991 (n8006, n_7791, n8002);
  and g13992 (n8007, n_7792, n8006);
  not g13993 (n_7796, n8002);
  and g13994 (n8008, n_7793, n_7796);
  not g13995 (n_7797, n8007);
  not g13996 (n_7798, n8008);
  and g13997 (n8009, n_7797, n_7798);
  not g13998 (n_7799, n8005);
  not g13999 (n_7800, n8009);
  and g14000 (n8010, n_7799, n_7800);
  not g14001 (n_7801, n7992);
  not g14002 (n_7802, n8010);
  and g14003 (n8011, n_7801, n_7802);
  not g14004 (n_7803, n7975);
  and g14005 (n8012, n_7803, n8011);
  not g14006 (n_7804, n8011);
  and g14007 (n8013, n7975, n_7804);
  not g14008 (n_7805, n8012);
  not g14009 (n_7806, n8013);
  and g14010 (n8014, n_7805, n_7806);
  not g14011 (n_7807, n7939);
  and g14012 (n8015, n_7807, n8014);
  not g14013 (n_7808, n8014);
  and g14014 (n8016, n7939, n_7808);
  not g14015 (n_7809, n8015);
  not g14016 (n_7810, n8016);
  and g14017 (n8017, n_7809, n_7810);
  not g14018 (n_7811, n7864);
  and g14019 (n8018, n_7811, n8017);
  not g14020 (n_7812, n8017);
  and g14021 (n8019, n7864, n_7812);
  not g14022 (n_7813, n8018);
  not g14023 (n_7814, n8019);
  and g14024 (n8020, n_7813, n_7814);
  not g14025 (n_7815, n7711);
  and g14026 (n8021, n_7815, n8020);
  not g14027 (n_7816, n8020);
  and g14028 (n8022, n7711, n_7816);
  not g14029 (n_7817, n8021);
  not g14030 (n_7818, n8022);
  and g14031 (n8023, n_7817, n_7818);
  not g14032 (n_7819, n7402);
  not g14033 (n_7820, n8023);
  and g14034 (n8024, n_7819, n_7820);
  not g14035 (n_7821, n7399);
  and g14036 (n8025, n_7821, n8024);
  not g14037 (n_7822, n7394);
  and g14038 (n8026, n_7822, n8025);
  and g14039 (n8027, n_7822, n_7821);
  not g14040 (n_7823, n8024);
  not g14041 (n_7824, n8027);
  and g14042 (n8028, n_7823, n_7824);
  not g14043 (n_7825, n8026);
  not g14044 (n_7826, n8028);
  and g14045 (n8029, n_7825, n_7826);
  and g14046 (n8030, n_7329, n_7327);
  not g14047 (n_7827, n8030);
  and g14048 (n8031, n_7328, n_7827);
  and g14049 (n8032, n_7285, n_7329);
  and g14050 (n8033, n_7286, n8032);
  and g14051 (n8034, n_7330, n8033);
  and g14052 (n8035, n_7285, n_7283);
  not g14053 (n_7828, n8035);
  and g14054 (n8036, n_7284, n_7828);
  not g14055 (n_7829, n8034);
  not g14056 (n_7830, n8036);
  and g14057 (n8037, n_7829, n_7830);
  not g14062 (n_7831, n8037);
  not g14063 (n_7832, n8041);
  and g14064 (n8042, n_7831, n_7832);
  not g14065 (n_7833, n8042);
  and g14066 (n8043, n8031, n_7833);
  and g14067 (n8044, n_7829, n8036);
  and g14068 (n8045, n8034, n_7830);
  not g14069 (n_7834, n8044);
  not g14070 (n_7835, n8045);
  and g14071 (n8046, n_7834, n_7835);
  not g14072 (n_7836, n8031);
  not g14073 (n_7837, n8046);
  and g14074 (n8047, n_7836, n_7837);
  and g14075 (n8048, n_7427, n_7428);
  not g14076 (n_7838, n8047);
  and g14077 (n8049, n_7838, n8048);
  not g14078 (n_7839, n8043);
  and g14079 (n8050, n_7839, n8049);
  and g14080 (n8051, n_7839, n_7838);
  not g14081 (n_7840, n8048);
  not g14082 (n_7841, n8051);
  and g14083 (n8052, n_7840, n_7841);
  not g14084 (n_7842, n8050);
  not g14085 (n_7843, n8052);
  and g14086 (n8053, n_7842, n_7843);
  and g14087 (n8054, n_7421, n_7419);
  not g14088 (n_7844, n8054);
  and g14089 (n8055, n_7420, n_7844);
  and g14090 (n8056, n_7377, n_7421);
  and g14091 (n8057, n_7378, n8056);
  and g14092 (n8058, n_7422, n8057);
  and g14093 (n8059, n_7377, n_7375);
  not g14094 (n_7845, n8059);
  and g14095 (n8060, n_7376, n_7845);
  not g14096 (n_7846, n8058);
  and g14097 (n8061, n_7846, n8060);
  not g14098 (n_7847, n8060);
  and g14099 (n8062, n8058, n_7847);
  not g14100 (n_7848, n8061);
  not g14101 (n_7849, n8062);
  and g14102 (n8063, n_7848, n_7849);
  not g14103 (n_7850, n8055);
  not g14104 (n_7851, n8063);
  and g14105 (n8064, n_7850, n_7851);
  and g14106 (n8065, n_7846, n_7847);
  not g14111 (n_7852, n8065);
  not g14112 (n_7853, n8069);
  and g14113 (n8070, n_7852, n_7853);
  not g14114 (n_7854, n8070);
  and g14115 (n8071, n8055, n_7854);
  not g14116 (n_7855, n8064);
  not g14117 (n_7856, n8071);
  and g14118 (n8072, n_7855, n_7856);
  not g14119 (n_7857, n8053);
  and g14120 (n8073, n_7857, n8072);
  and g14121 (n8074, n_7838, n_7840);
  and g14122 (n8075, n_7839, n8074);
  and g14123 (n8076, n8048, n_7841);
  not g14124 (n_7858, n8075);
  not g14125 (n_7859, n8076);
  and g14126 (n8077, n_7858, n_7859);
  not g14127 (n_7860, n8072);
  not g14128 (n_7861, n8077);
  and g14129 (n8078, n_7860, n_7861);
  not g14130 (n_7862, n8073);
  not g14131 (n_7863, n8078);
  and g14132 (n8079, n_7862, n_7863);
  and g14133 (n8080, n_7233, n_7231);
  not g14134 (n_7864, n8080);
  and g14135 (n8081, n_7232, n_7864);
  and g14136 (n8082, n_7189, n_7233);
  and g14137 (n8083, n_7190, n8082);
  and g14138 (n8084, n_7234, n8083);
  and g14139 (n8085, n_7189, n_7187);
  not g14140 (n_7865, n8085);
  and g14141 (n8086, n_7188, n_7865);
  not g14142 (n_7866, n8084);
  and g14143 (n8087, n_7866, n8086);
  not g14144 (n_7867, n8086);
  and g14145 (n8088, n8084, n_7867);
  not g14146 (n_7868, n8087);
  not g14147 (n_7869, n8088);
  and g14148 (n8089, n_7868, n_7869);
  not g14149 (n_7870, n8081);
  not g14150 (n_7871, n8089);
  and g14151 (n8090, n_7870, n_7871);
  and g14152 (n8091, n_7866, n_7867);
  not g14157 (n_7872, n8091);
  not g14158 (n_7873, n8095);
  and g14159 (n8096, n_7872, n_7873);
  not g14160 (n_7874, n8096);
  and g14161 (n8097, n8081, n_7874);
  not g14162 (n_7875, n8090);
  not g14163 (n_7876, n8097);
  and g14164 (n8098, n_7875, n_7876);
  and g14165 (n8099, n_7141, n_7139);
  not g14166 (n_7877, n8099);
  and g14167 (n8100, n_7140, n_7877);
  and g14168 (n8101, n_7097, n_7141);
  and g14169 (n8102, n_7098, n8101);
  and g14170 (n8103, n_7142, n8102);
  and g14171 (n8104, n_7097, n_7095);
  not g14172 (n_7878, n8104);
  and g14173 (n8105, n_7096, n_7878);
  not g14174 (n_7879, n8103);
  not g14175 (n_7880, n8105);
  and g14176 (n8106, n_7879, n_7880);
  not g14181 (n_7881, n8106);
  not g14182 (n_7882, n8110);
  and g14183 (n8111, n_7881, n_7882);
  not g14184 (n_7883, n8111);
  and g14185 (n8112, n8100, n_7883);
  and g14186 (n8113, n_7879, n8105);
  and g14187 (n8114, n8103, n_7880);
  not g14188 (n_7884, n8113);
  not g14189 (n_7885, n8114);
  and g14190 (n8115, n_7884, n_7885);
  not g14191 (n_7886, n8100);
  not g14192 (n_7887, n8115);
  and g14193 (n8116, n_7886, n_7887);
  and g14194 (n8117, n_7239, n_7240);
  not g14195 (n_7888, n8116);
  not g14196 (n_7889, n8117);
  and g14197 (n8118, n_7888, n_7889);
  not g14198 (n_7890, n8112);
  and g14199 (n8119, n_7890, n8118);
  and g14200 (n8120, n_7890, n_7888);
  not g14201 (n_7891, n8120);
  and g14202 (n8121, n8117, n_7891);
  not g14203 (n_7892, n8119);
  not g14204 (n_7893, n8121);
  and g14205 (n8122, n_7892, n_7893);
  not g14206 (n_7894, n8098);
  not g14207 (n_7895, n8122);
  and g14208 (n8123, n_7894, n_7895);
  and g14209 (n8124, n_7888, n8117);
  and g14210 (n8125, n_7890, n8124);
  and g14211 (n8126, n_7889, n_7891);
  not g14212 (n_7896, n8125);
  not g14213 (n_7897, n8126);
  and g14214 (n8127, n_7896, n_7897);
  not g14215 (n_7898, n8127);
  and g14216 (n8128, n8098, n_7898);
  and g14217 (n8129, n_7431, n_7432);
  not g14218 (n_7899, n8128);
  not g14219 (n_7900, n8129);
  and g14220 (n8130, n_7899, n_7900);
  not g14221 (n_7901, n8123);
  and g14222 (n8131, n_7901, n8130);
  and g14223 (n8132, n_7901, n_7899);
  not g14224 (n_7902, n8132);
  and g14225 (n8133, n8129, n_7902);
  not g14226 (n_7903, n8131);
  not g14227 (n_7904, n8133);
  and g14228 (n8134, n_7903, n_7904);
  not g14229 (n_7905, n8079);
  not g14230 (n_7906, n8134);
  and g14231 (n8135, n_7905, n_7906);
  and g14232 (n8136, n_7899, n8129);
  and g14233 (n8137, n_7901, n8136);
  and g14234 (n8138, n_7900, n_7902);
  not g14235 (n_7907, n8137);
  not g14236 (n_7908, n8138);
  and g14237 (n8139, n_7907, n_7908);
  not g14238 (n_7909, n8139);
  and g14239 (n8140, n8079, n_7909);
  and g14240 (n8141, n_7815, n_7816);
  not g14241 (n_7910, n8140);
  and g14242 (n8142, n_7910, n8141);
  not g14243 (n_7911, n8135);
  and g14244 (n8143, n_7911, n8142);
  and g14245 (n8144, n_7911, n_7910);
  not g14246 (n_7912, n8141);
  not g14247 (n_7913, n8144);
  and g14248 (n8145, n_7912, n_7913);
  not g14249 (n_7914, n8143);
  not g14250 (n_7915, n8145);
  and g14251 (n8146, n_7914, n_7915);
  and g14252 (n8147, n_7613, n_7611);
  not g14253 (n_7916, n8147);
  and g14254 (n8148, n_7612, n_7916);
  and g14255 (n8149, n_7569, n_7613);
  and g14256 (n8150, n_7570, n8149);
  and g14257 (n8151, n_7614, n8150);
  and g14258 (n8152, n_7569, n_7567);
  not g14259 (n_7917, n8152);
  and g14260 (n8153, n_7568, n_7917);
  not g14261 (n_7918, n8151);
  and g14262 (n8154, n_7918, n8153);
  not g14263 (n_7919, n8153);
  and g14264 (n8155, n8151, n_7919);
  not g14265 (n_7920, n8154);
  not g14266 (n_7921, n8155);
  and g14267 (n8156, n_7920, n_7921);
  not g14268 (n_7922, n8148);
  not g14269 (n_7923, n8156);
  and g14270 (n8157, n_7922, n_7923);
  and g14271 (n8158, n_7918, n_7919);
  not g14276 (n_7924, n8158);
  not g14277 (n_7925, n8162);
  and g14278 (n8163, n_7924, n_7925);
  not g14279 (n_7926, n8163);
  and g14280 (n8164, n8148, n_7926);
  not g14281 (n_7927, n8157);
  not g14282 (n_7928, n8164);
  and g14283 (n8165, n_7927, n_7928);
  and g14284 (n8166, n_7521, n_7519);
  not g14285 (n_7929, n8166);
  and g14286 (n8167, n_7520, n_7929);
  and g14287 (n8168, n_7477, n_7521);
  and g14288 (n8169, n_7478, n8168);
  and g14289 (n8170, n_7522, n8169);
  and g14290 (n8171, n_7477, n_7475);
  not g14291 (n_7930, n8171);
  and g14292 (n8172, n_7476, n_7930);
  not g14293 (n_7931, n8170);
  not g14294 (n_7932, n8172);
  and g14295 (n8173, n_7931, n_7932);
  not g14300 (n_7933, n8173);
  not g14301 (n_7934, n8177);
  and g14302 (n8178, n_7933, n_7934);
  not g14303 (n_7935, n8178);
  and g14304 (n8179, n8167, n_7935);
  and g14305 (n8180, n_7931, n8172);
  and g14306 (n8181, n8170, n_7932);
  not g14307 (n_7936, n8180);
  not g14308 (n_7937, n8181);
  and g14309 (n8182, n_7936, n_7937);
  not g14310 (n_7938, n8167);
  not g14311 (n_7939, n8182);
  and g14312 (n8183, n_7938, n_7939);
  and g14313 (n8184, n_7619, n_7620);
  not g14314 (n_7940, n8183);
  not g14315 (n_7941, n8184);
  and g14316 (n8185, n_7940, n_7941);
  not g14317 (n_7942, n8179);
  and g14318 (n8186, n_7942, n8185);
  and g14319 (n8187, n_7942, n_7940);
  not g14320 (n_7943, n8187);
  and g14321 (n8188, n8184, n_7943);
  not g14322 (n_7944, n8186);
  not g14323 (n_7945, n8188);
  and g14324 (n8189, n_7944, n_7945);
  not g14325 (n_7946, n8165);
  not g14326 (n_7947, n8189);
  and g14327 (n8190, n_7946, n_7947);
  and g14328 (n8191, n_7940, n8184);
  and g14329 (n8192, n_7942, n8191);
  and g14330 (n8193, n_7941, n_7943);
  not g14331 (n_7948, n8192);
  not g14332 (n_7949, n8193);
  and g14333 (n8194, n_7948, n_7949);
  not g14334 (n_7950, n8194);
  and g14335 (n8195, n8165, n_7950);
  and g14336 (n8196, n_7811, n_7812);
  not g14337 (n_7951, n8195);
  and g14338 (n8197, n_7951, n8196);
  not g14339 (n_7952, n8190);
  and g14340 (n8198, n_7952, n8197);
  and g14341 (n8199, n_7952, n_7951);
  not g14342 (n_7953, n8196);
  not g14343 (n_7954, n8199);
  and g14344 (n8200, n_7953, n_7954);
  not g14345 (n_7955, n8198);
  not g14346 (n_7956, n8200);
  and g14347 (n8201, n_7955, n_7956);
  and g14348 (n8202, n_7709, n_7707);
  not g14349 (n_7957, n8202);
  and g14350 (n8203, n_7708, n_7957);
  and g14351 (n8204, n_7665, n_7709);
  and g14352 (n8205, n_7666, n8204);
  and g14353 (n8206, n_7710, n8205);
  and g14354 (n8207, n_7665, n_7663);
  not g14355 (n_7958, n8207);
  and g14356 (n8208, n_7664, n_7958);
  not g14357 (n_7959, n8206);
  not g14358 (n_7960, n8208);
  and g14359 (n8209, n_7959, n_7960);
  not g14364 (n_7961, n8209);
  not g14365 (n_7962, n8213);
  and g14366 (n8214, n_7961, n_7962);
  not g14367 (n_7963, n8214);
  and g14368 (n8215, n8203, n_7963);
  and g14369 (n8216, n_7959, n8208);
  and g14370 (n8217, n8206, n_7960);
  not g14371 (n_7964, n8216);
  not g14372 (n_7965, n8217);
  and g14373 (n8218, n_7964, n_7965);
  not g14374 (n_7966, n8203);
  not g14375 (n_7967, n8218);
  and g14376 (n8219, n_7966, n_7967);
  and g14377 (n8220, n_7807, n_7808);
  not g14378 (n_7968, n8219);
  and g14379 (n8221, n_7968, n8220);
  not g14380 (n_7969, n8215);
  and g14381 (n8222, n_7969, n8221);
  and g14382 (n8223, n_7969, n_7968);
  not g14383 (n_7970, n8220);
  not g14384 (n_7971, n8223);
  and g14385 (n8224, n_7970, n_7971);
  not g14386 (n_7972, n8222);
  not g14387 (n_7973, n8224);
  and g14388 (n8225, n_7972, n_7973);
  and g14389 (n8226, n_7801, n_7799);
  not g14390 (n_7974, n8226);
  and g14391 (n8227, n_7800, n_7974);
  and g14392 (n8228, n_7757, n_7801);
  and g14393 (n8229, n_7758, n8228);
  and g14394 (n8230, n_7802, n8229);
  and g14395 (n8231, n_7757, n_7755);
  not g14396 (n_7975, n8231);
  and g14397 (n8232, n_7756, n_7975);
  not g14398 (n_7976, n8230);
  and g14399 (n8233, n_7976, n8232);
  not g14400 (n_7977, n8232);
  and g14401 (n8234, n8230, n_7977);
  not g14402 (n_7978, n8233);
  not g14403 (n_7979, n8234);
  and g14404 (n8235, n_7978, n_7979);
  not g14405 (n_7980, n8227);
  not g14406 (n_7981, n8235);
  and g14407 (n8236, n_7980, n_7981);
  and g14408 (n8237, n_7976, n_7977);
  not g14413 (n_7982, n8237);
  not g14414 (n_7983, n8241);
  and g14415 (n8242, n_7982, n_7983);
  not g14416 (n_7984, n8242);
  and g14417 (n8243, n8227, n_7984);
  not g14418 (n_7985, n8236);
  not g14419 (n_7986, n8243);
  and g14420 (n8244, n_7985, n_7986);
  not g14421 (n_7987, n8225);
  and g14422 (n8245, n_7987, n8244);
  and g14423 (n8246, n_7968, n_7970);
  and g14424 (n8247, n_7969, n8246);
  and g14425 (n8248, n8220, n_7971);
  not g14426 (n_7988, n8247);
  not g14427 (n_7989, n8248);
  and g14428 (n8249, n_7988, n_7989);
  not g14429 (n_7990, n8244);
  not g14430 (n_7991, n8249);
  and g14431 (n8250, n_7990, n_7991);
  not g14432 (n_7992, n8245);
  not g14433 (n_7993, n8250);
  and g14434 (n8251, n_7992, n_7993);
  not g14435 (n_7994, n8201);
  and g14436 (n8252, n_7994, n8251);
  and g14437 (n8253, n_7951, n_7953);
  and g14438 (n8254, n_7952, n8253);
  and g14439 (n8255, n8196, n_7954);
  not g14440 (n_7995, n8254);
  not g14441 (n_7996, n8255);
  and g14442 (n8256, n_7995, n_7996);
  not g14443 (n_7997, n8251);
  not g14444 (n_7998, n8256);
  and g14445 (n8257, n_7997, n_7998);
  not g14446 (n_7999, n8252);
  not g14447 (n_8000, n8257);
  and g14448 (n8258, n_7999, n_8000);
  not g14449 (n_8001, n8146);
  and g14450 (n8259, n_8001, n8258);
  and g14451 (n8260, n_7910, n_7912);
  and g14452 (n8261, n_7911, n8260);
  and g14453 (n8262, n8141, n_7913);
  not g14454 (n_8002, n8261);
  not g14455 (n_8003, n8262);
  and g14456 (n8263, n_8002, n_8003);
  not g14457 (n_8004, n8258);
  not g14458 (n_8005, n8263);
  and g14459 (n8264, n_8004, n_8005);
  not g14460 (n_8006, n8259);
  not g14461 (n_8007, n8264);
  and g14462 (n8265, n_8006, n_8007);
  not g14463 (n_8008, n8029);
  and g14464 (n8266, n_8008, n8265);
  and g14465 (n8267, n_7821, n_7823);
  and g14466 (n8268, n_7822, n8267);
  and g14467 (n8269, n8024, n_7824);
  not g14468 (n_8009, n8268);
  not g14469 (n_8010, n8269);
  and g14470 (n8270, n_8009, n_8010);
  not g14471 (n_8011, n8265);
  not g14472 (n_8012, n8270);
  and g14473 (n8271, n_8011, n_8012);
  not g14474 (n_8013, n8266);
  not g14475 (n_8014, n8271);
  and g14476 (n8272, n_8013, n_8014);
  and g14477 (n8273, \A[334] , \A[335] );
  not g14478 (n_8017, \A[335] );
  and g14479 (n8274, \A[334] , n_8017);
  not g14480 (n_8018, \A[334] );
  and g14481 (n8275, n_8018, \A[335] );
  not g14482 (n_8019, n8274);
  not g14483 (n_8020, n8275);
  and g14484 (n8276, n_8019, n_8020);
  not g14485 (n_8022, n8276);
  and g14486 (n8277, \A[336] , n_8022);
  not g14487 (n_8023, n8273);
  not g14488 (n_8024, n8277);
  and g14489 (n8278, n_8023, n_8024);
  and g14490 (n8279, \A[331] , \A[332] );
  not g14491 (n_8027, \A[332] );
  and g14492 (n8280, \A[331] , n_8027);
  not g14493 (n_8028, \A[331] );
  and g14494 (n8281, n_8028, \A[332] );
  not g14495 (n_8029, n8280);
  not g14496 (n_8030, n8281);
  and g14497 (n8282, n_8029, n_8030);
  not g14498 (n_8032, n8282);
  and g14499 (n8283, \A[333] , n_8032);
  not g14500 (n_8033, n8279);
  not g14501 (n_8034, n8283);
  and g14502 (n8284, n_8033, n_8034);
  not g14503 (n_8035, n8284);
  and g14504 (n8285, n8278, n_8035);
  not g14505 (n_8036, n8278);
  and g14506 (n8286, n_8036, n8284);
  and g14507 (n8287, \A[333] , n_8029);
  and g14508 (n8288, n_8030, n8287);
  not g14509 (n_8037, \A[333] );
  and g14510 (n8289, n_8037, n_8032);
  not g14511 (n_8038, n8288);
  not g14512 (n_8039, n8289);
  and g14513 (n8290, n_8038, n_8039);
  and g14514 (n8291, \A[336] , n_8019);
  and g14515 (n8292, n_8020, n8291);
  not g14516 (n_8040, \A[336] );
  and g14517 (n8293, n_8040, n_8022);
  not g14518 (n_8041, n8292);
  not g14519 (n_8042, n8293);
  and g14520 (n8294, n_8041, n_8042);
  not g14521 (n_8043, n8290);
  not g14522 (n_8044, n8294);
  and g14523 (n8295, n_8043, n_8044);
  not g14524 (n_8045, n8286);
  and g14525 (n8296, n_8045, n8295);
  not g14526 (n_8046, n8285);
  and g14527 (n8297, n_8046, n8296);
  and g14528 (n8298, n_8046, n_8045);
  not g14529 (n_8047, n8295);
  not g14530 (n_8048, n8298);
  and g14531 (n8299, n_8047, n_8048);
  not g14532 (n_8049, n8297);
  not g14533 (n_8050, n8299);
  and g14534 (n8300, n_8049, n_8050);
  and g14535 (n8301, n_8043, n8294);
  and g14536 (n8302, n8290, n_8044);
  not g14537 (n_8051, n8301);
  not g14538 (n_8052, n8302);
  and g14539 (n8303, n_8051, n_8052);
  and g14540 (n8304, n8295, n_8048);
  and g14541 (n8305, n_8036, n_8035);
  not g14542 (n_8053, n8304);
  not g14543 (n_8054, n8305);
  and g14544 (n8306, n_8053, n_8054);
  not g14545 (n_8055, n8303);
  not g14546 (n_8056, n8306);
  and g14547 (n8307, n_8055, n_8056);
  not g14548 (n_8057, n8300);
  not g14549 (n_8058, n8307);
  and g14550 (n8308, n_8057, n_8058);
  and g14551 (n8309, n_8057, n_8056);
  and g14552 (n8310, \A[340] , \A[341] );
  not g14553 (n_8061, \A[341] );
  and g14554 (n8311, \A[340] , n_8061);
  not g14555 (n_8062, \A[340] );
  and g14556 (n8312, n_8062, \A[341] );
  not g14557 (n_8063, n8311);
  not g14558 (n_8064, n8312);
  and g14559 (n8313, n_8063, n_8064);
  not g14560 (n_8066, n8313);
  and g14561 (n8314, \A[342] , n_8066);
  not g14562 (n_8067, n8310);
  not g14563 (n_8068, n8314);
  and g14564 (n8315, n_8067, n_8068);
  and g14565 (n8316, \A[337] , \A[338] );
  not g14566 (n_8071, \A[338] );
  and g14567 (n8317, \A[337] , n_8071);
  not g14568 (n_8072, \A[337] );
  and g14569 (n8318, n_8072, \A[338] );
  not g14570 (n_8073, n8317);
  not g14571 (n_8074, n8318);
  and g14572 (n8319, n_8073, n_8074);
  not g14573 (n_8076, n8319);
  and g14574 (n8320, \A[339] , n_8076);
  not g14575 (n_8077, n8316);
  not g14576 (n_8078, n8320);
  and g14577 (n8321, n_8077, n_8078);
  not g14578 (n_8079, n8315);
  and g14579 (n8322, n_8079, n8321);
  not g14580 (n_8080, n8321);
  and g14581 (n8323, n8315, n_8080);
  not g14582 (n_8081, n8322);
  not g14583 (n_8082, n8323);
  and g14584 (n8324, n_8081, n_8082);
  and g14585 (n8325, \A[339] , n_8073);
  and g14586 (n8326, n_8074, n8325);
  not g14587 (n_8083, \A[339] );
  and g14588 (n8327, n_8083, n_8076);
  not g14589 (n_8084, n8326);
  not g14590 (n_8085, n8327);
  and g14591 (n8328, n_8084, n_8085);
  and g14592 (n8329, \A[342] , n_8063);
  and g14593 (n8330, n_8064, n8329);
  not g14594 (n_8086, \A[342] );
  and g14595 (n8331, n_8086, n_8066);
  not g14596 (n_8087, n8330);
  not g14597 (n_8088, n8331);
  and g14598 (n8332, n_8087, n_8088);
  not g14599 (n_8089, n8328);
  not g14600 (n_8090, n8332);
  and g14601 (n8333, n_8089, n_8090);
  not g14602 (n_8091, n8324);
  and g14603 (n8334, n_8091, n8333);
  and g14604 (n8335, n_8079, n_8080);
  not g14605 (n_8092, n8334);
  not g14606 (n_8093, n8335);
  and g14607 (n8336, n_8092, n_8093);
  and g14608 (n8337, n_8081, n8333);
  and g14609 (n8338, n_8082, n8337);
  not g14610 (n_8094, n8333);
  and g14611 (n8339, n_8091, n_8094);
  not g14612 (n_8095, n8338);
  not g14613 (n_8096, n8339);
  and g14614 (n8340, n_8095, n_8096);
  not g14615 (n_8097, n8336);
  not g14616 (n_8098, n8340);
  and g14617 (n8341, n_8097, n_8098);
  and g14618 (n8342, n_8089, n8332);
  and g14619 (n8343, n8328, n_8090);
  not g14620 (n_8099, n8342);
  not g14621 (n_8100, n8343);
  and g14622 (n8344, n_8099, n_8100);
  not g14623 (n_8101, n8344);
  and g14624 (n8345, n_8055, n_8101);
  not g14625 (n_8102, n8341);
  and g14626 (n8346, n_8102, n8345);
  not g14627 (n_8103, n8309);
  and g14628 (n8347, n_8103, n8346);
  and g14629 (n8348, n_8097, n_8101);
  not g14630 (n_8104, n8348);
  and g14631 (n8349, n_8098, n_8104);
  not g14632 (n_8105, n8347);
  not g14633 (n_8106, n8349);
  and g14634 (n8350, n_8105, n_8106);
  not g14639 (n_8107, n8350);
  not g14640 (n_8108, n8354);
  and g14641 (n8355, n_8107, n_8108);
  not g14642 (n_8109, n8355);
  and g14643 (n8356, n8308, n_8109);
  and g14644 (n8357, n_8105, n8349);
  and g14645 (n8358, n8347, n_8106);
  not g14646 (n_8110, n8357);
  not g14647 (n_8111, n8358);
  and g14648 (n8359, n_8110, n_8111);
  not g14649 (n_8112, n8308);
  not g14650 (n_8113, n8359);
  and g14651 (n8360, n_8112, n_8113);
  and g14652 (n8361, n_8102, n_8101);
  and g14653 (n8362, n_8055, n_8103);
  not g14654 (n_8114, n8361);
  and g14655 (n8363, n_8114, n8362);
  not g14656 (n_8115, n8362);
  and g14657 (n8364, n8361, n_8115);
  not g14658 (n_8116, n8363);
  not g14659 (n_8117, n8364);
  and g14660 (n8365, n_8116, n_8117);
  not g14661 (n_8119, \A[325] );
  and g14662 (n8366, n_8119, \A[326] );
  not g14663 (n_8121, \A[326] );
  and g14664 (n8367, \A[325] , n_8121);
  not g14665 (n_8123, n8367);
  and g14666 (n8368, \A[327] , n_8123);
  not g14667 (n_8124, n8366);
  and g14668 (n8369, n_8124, n8368);
  and g14669 (n8370, n_8124, n_8123);
  not g14670 (n_8125, \A[327] );
  not g14671 (n_8126, n8370);
  and g14672 (n8371, n_8125, n_8126);
  not g14673 (n_8127, n8369);
  not g14674 (n_8128, n8371);
  and g14675 (n8372, n_8127, n_8128);
  not g14676 (n_8130, \A[328] );
  and g14677 (n8373, n_8130, \A[329] );
  not g14678 (n_8132, \A[329] );
  and g14679 (n8374, \A[328] , n_8132);
  not g14680 (n_8134, n8374);
  and g14681 (n8375, \A[330] , n_8134);
  not g14682 (n_8135, n8373);
  and g14683 (n8376, n_8135, n8375);
  and g14684 (n8377, n_8135, n_8134);
  not g14685 (n_8136, \A[330] );
  not g14686 (n_8137, n8377);
  and g14687 (n8378, n_8136, n_8137);
  not g14688 (n_8138, n8376);
  not g14689 (n_8139, n8378);
  and g14690 (n8379, n_8138, n_8139);
  not g14691 (n_8140, n8372);
  and g14692 (n8380, n_8140, n8379);
  not g14693 (n_8141, n8379);
  and g14694 (n8381, n8372, n_8141);
  not g14695 (n_8142, n8380);
  not g14696 (n_8143, n8381);
  and g14697 (n8382, n_8142, n_8143);
  and g14698 (n8383, \A[328] , \A[329] );
  and g14699 (n8384, \A[330] , n_8137);
  not g14700 (n_8144, n8383);
  not g14701 (n_8145, n8384);
  and g14702 (n8385, n_8144, n_8145);
  and g14703 (n8386, \A[325] , \A[326] );
  and g14704 (n8387, \A[327] , n_8126);
  not g14705 (n_8146, n8386);
  not g14706 (n_8147, n8387);
  and g14707 (n8388, n_8146, n_8147);
  not g14708 (n_8148, n8385);
  and g14709 (n8389, n_8148, n8388);
  not g14710 (n_8149, n8388);
  and g14711 (n8390, n8385, n_8149);
  not g14712 (n_8150, n8389);
  not g14713 (n_8151, n8390);
  and g14714 (n8391, n_8150, n_8151);
  and g14715 (n8392, n_8140, n_8141);
  not g14716 (n_8152, n8391);
  and g14717 (n8393, n_8152, n8392);
  and g14718 (n8394, n_8148, n_8149);
  not g14719 (n_8153, n8393);
  not g14720 (n_8154, n8394);
  and g14721 (n8395, n_8153, n_8154);
  and g14722 (n8396, n_8150, n8392);
  and g14723 (n8397, n_8151, n8396);
  not g14724 (n_8155, n8392);
  and g14725 (n8398, n_8152, n_8155);
  not g14726 (n_8156, n8397);
  not g14727 (n_8157, n8398);
  and g14728 (n8399, n_8156, n_8157);
  not g14729 (n_8158, n8395);
  not g14730 (n_8159, n8399);
  and g14731 (n8400, n_8158, n_8159);
  not g14732 (n_8160, n8382);
  not g14733 (n_8161, n8400);
  and g14734 (n8401, n_8160, n_8161);
  not g14735 (n_8163, \A[319] );
  and g14736 (n8402, n_8163, \A[320] );
  not g14737 (n_8165, \A[320] );
  and g14738 (n8403, \A[319] , n_8165);
  not g14739 (n_8167, n8403);
  and g14740 (n8404, \A[321] , n_8167);
  not g14741 (n_8168, n8402);
  and g14742 (n8405, n_8168, n8404);
  and g14743 (n8406, n_8168, n_8167);
  not g14744 (n_8169, \A[321] );
  not g14745 (n_8170, n8406);
  and g14746 (n8407, n_8169, n_8170);
  not g14747 (n_8171, n8405);
  not g14748 (n_8172, n8407);
  and g14749 (n8408, n_8171, n_8172);
  not g14750 (n_8174, \A[322] );
  and g14751 (n8409, n_8174, \A[323] );
  not g14752 (n_8176, \A[323] );
  and g14753 (n8410, \A[322] , n_8176);
  not g14754 (n_8178, n8410);
  and g14755 (n8411, \A[324] , n_8178);
  not g14756 (n_8179, n8409);
  and g14757 (n8412, n_8179, n8411);
  and g14758 (n8413, n_8179, n_8178);
  not g14759 (n_8180, \A[324] );
  not g14760 (n_8181, n8413);
  and g14761 (n8414, n_8180, n_8181);
  not g14762 (n_8182, n8412);
  not g14763 (n_8183, n8414);
  and g14764 (n8415, n_8182, n_8183);
  not g14765 (n_8184, n8408);
  and g14766 (n8416, n_8184, n8415);
  not g14767 (n_8185, n8415);
  and g14768 (n8417, n8408, n_8185);
  not g14769 (n_8186, n8416);
  not g14770 (n_8187, n8417);
  and g14771 (n8418, n_8186, n_8187);
  and g14772 (n8419, \A[322] , \A[323] );
  and g14773 (n8420, \A[324] , n_8181);
  not g14774 (n_8188, n8419);
  not g14775 (n_8189, n8420);
  and g14776 (n8421, n_8188, n_8189);
  and g14777 (n8422, \A[319] , \A[320] );
  and g14778 (n8423, \A[321] , n_8170);
  not g14779 (n_8190, n8422);
  not g14780 (n_8191, n8423);
  and g14781 (n8424, n_8190, n_8191);
  not g14782 (n_8192, n8421);
  and g14783 (n8425, n_8192, n8424);
  not g14784 (n_8193, n8424);
  and g14785 (n8426, n8421, n_8193);
  not g14786 (n_8194, n8425);
  not g14787 (n_8195, n8426);
  and g14788 (n8427, n_8194, n_8195);
  and g14789 (n8428, n_8184, n_8185);
  not g14790 (n_8196, n8427);
  and g14791 (n8429, n_8196, n8428);
  and g14792 (n8430, n_8192, n_8193);
  not g14793 (n_8197, n8429);
  not g14794 (n_8198, n8430);
  and g14795 (n8431, n_8197, n_8198);
  and g14796 (n8432, n_8194, n8428);
  and g14797 (n8433, n_8195, n8432);
  not g14798 (n_8199, n8428);
  and g14799 (n8434, n_8196, n_8199);
  not g14800 (n_8200, n8433);
  not g14801 (n_8201, n8434);
  and g14802 (n8435, n_8200, n_8201);
  not g14803 (n_8202, n8431);
  not g14804 (n_8203, n8435);
  and g14805 (n8436, n_8202, n_8203);
  not g14806 (n_8204, n8418);
  not g14807 (n_8205, n8436);
  and g14808 (n8437, n_8204, n_8205);
  not g14809 (n_8206, n8401);
  and g14810 (n8438, n_8206, n8437);
  not g14811 (n_8207, n8437);
  and g14812 (n8439, n8401, n_8207);
  not g14813 (n_8208, n8438);
  not g14814 (n_8209, n8439);
  and g14815 (n8440, n_8208, n_8209);
  not g14816 (n_8210, n8365);
  not g14817 (n_8211, n8440);
  and g14818 (n8441, n_8210, n_8211);
  not g14819 (n_8212, n8360);
  and g14820 (n8442, n_8212, n8441);
  not g14821 (n_8213, n8356);
  and g14822 (n8443, n_8213, n8442);
  and g14823 (n8444, n_8213, n_8212);
  not g14824 (n_8214, n8441);
  not g14825 (n_8215, n8444);
  and g14826 (n8445, n_8214, n_8215);
  not g14827 (n_8216, n8443);
  not g14828 (n_8217, n8445);
  and g14829 (n8446, n_8216, n_8217);
  and g14830 (n8447, n_8204, n_8202);
  not g14831 (n_8218, n8447);
  and g14832 (n8448, n_8203, n_8218);
  and g14833 (n8449, n_8160, n_8204);
  and g14834 (n8450, n_8161, n8449);
  and g14835 (n8451, n_8205, n8450);
  and g14836 (n8452, n_8160, n_8158);
  not g14837 (n_8219, n8452);
  and g14838 (n8453, n_8159, n_8219);
  not g14839 (n_8220, n8451);
  and g14840 (n8454, n_8220, n8453);
  not g14841 (n_8221, n8453);
  and g14842 (n8455, n8451, n_8221);
  not g14843 (n_8222, n8454);
  not g14844 (n_8223, n8455);
  and g14845 (n8456, n_8222, n_8223);
  not g14846 (n_8224, n8448);
  not g14847 (n_8225, n8456);
  and g14848 (n8457, n_8224, n_8225);
  and g14849 (n8458, n_8220, n_8221);
  not g14854 (n_8226, n8458);
  not g14855 (n_8227, n8462);
  and g14856 (n8463, n_8226, n_8227);
  not g14857 (n_8228, n8463);
  and g14858 (n8464, n8448, n_8228);
  not g14859 (n_8229, n8457);
  not g14860 (n_8230, n8464);
  and g14861 (n8465, n_8229, n_8230);
  not g14862 (n_8231, n8446);
  and g14863 (n8466, n_8231, n8465);
  and g14864 (n8467, n_8212, n_8214);
  and g14865 (n8468, n_8213, n8467);
  and g14866 (n8469, n8441, n_8215);
  not g14867 (n_8232, n8468);
  not g14868 (n_8233, n8469);
  and g14869 (n8470, n_8232, n_8233);
  not g14870 (n_8234, n8465);
  not g14871 (n_8235, n8470);
  and g14872 (n8471, n_8234, n_8235);
  not g14873 (n_8236, n8466);
  not g14874 (n_8237, n8471);
  and g14875 (n8472, n_8236, n_8237);
  and g14876 (n8473, \A[346] , \A[347] );
  not g14877 (n_8240, \A[347] );
  and g14878 (n8474, \A[346] , n_8240);
  not g14879 (n_8241, \A[346] );
  and g14880 (n8475, n_8241, \A[347] );
  not g14881 (n_8242, n8474);
  not g14882 (n_8243, n8475);
  and g14883 (n8476, n_8242, n_8243);
  not g14884 (n_8245, n8476);
  and g14885 (n8477, \A[348] , n_8245);
  not g14886 (n_8246, n8473);
  not g14887 (n_8247, n8477);
  and g14888 (n8478, n_8246, n_8247);
  and g14889 (n8479, \A[343] , \A[344] );
  not g14890 (n_8250, \A[344] );
  and g14891 (n8480, \A[343] , n_8250);
  not g14892 (n_8251, \A[343] );
  and g14893 (n8481, n_8251, \A[344] );
  not g14894 (n_8252, n8480);
  not g14895 (n_8253, n8481);
  and g14896 (n8482, n_8252, n_8253);
  not g14897 (n_8255, n8482);
  and g14898 (n8483, \A[345] , n_8255);
  not g14899 (n_8256, n8479);
  not g14900 (n_8257, n8483);
  and g14901 (n8484, n_8256, n_8257);
  not g14902 (n_8258, n8484);
  and g14903 (n8485, n8478, n_8258);
  not g14904 (n_8259, n8478);
  and g14905 (n8486, n_8259, n8484);
  and g14906 (n8487, \A[345] , n_8252);
  and g14907 (n8488, n_8253, n8487);
  not g14908 (n_8260, \A[345] );
  and g14909 (n8489, n_8260, n_8255);
  not g14910 (n_8261, n8488);
  not g14911 (n_8262, n8489);
  and g14912 (n8490, n_8261, n_8262);
  and g14913 (n8491, \A[348] , n_8242);
  and g14914 (n8492, n_8243, n8491);
  not g14915 (n_8263, \A[348] );
  and g14916 (n8493, n_8263, n_8245);
  not g14917 (n_8264, n8492);
  not g14918 (n_8265, n8493);
  and g14919 (n8494, n_8264, n_8265);
  not g14920 (n_8266, n8490);
  not g14921 (n_8267, n8494);
  and g14922 (n8495, n_8266, n_8267);
  not g14923 (n_8268, n8486);
  and g14924 (n8496, n_8268, n8495);
  not g14925 (n_8269, n8485);
  and g14926 (n8497, n_8269, n8496);
  and g14927 (n8498, n_8269, n_8268);
  not g14928 (n_8270, n8495);
  not g14929 (n_8271, n8498);
  and g14930 (n8499, n_8270, n_8271);
  not g14931 (n_8272, n8497);
  not g14932 (n_8273, n8499);
  and g14933 (n8500, n_8272, n_8273);
  and g14934 (n8501, n_8266, n8494);
  and g14935 (n8502, n8490, n_8267);
  not g14936 (n_8274, n8501);
  not g14937 (n_8275, n8502);
  and g14938 (n8503, n_8274, n_8275);
  and g14939 (n8504, n8495, n_8271);
  and g14940 (n8505, n_8259, n_8258);
  not g14941 (n_8276, n8504);
  not g14942 (n_8277, n8505);
  and g14943 (n8506, n_8276, n_8277);
  not g14944 (n_8278, n8503);
  not g14945 (n_8279, n8506);
  and g14946 (n8507, n_8278, n_8279);
  not g14947 (n_8280, n8500);
  not g14948 (n_8281, n8507);
  and g14949 (n8508, n_8280, n_8281);
  and g14950 (n8509, n_8280, n_8279);
  and g14951 (n8510, \A[352] , \A[353] );
  not g14952 (n_8284, \A[353] );
  and g14953 (n8511, \A[352] , n_8284);
  not g14954 (n_8285, \A[352] );
  and g14955 (n8512, n_8285, \A[353] );
  not g14956 (n_8286, n8511);
  not g14957 (n_8287, n8512);
  and g14958 (n8513, n_8286, n_8287);
  not g14959 (n_8289, n8513);
  and g14960 (n8514, \A[354] , n_8289);
  not g14961 (n_8290, n8510);
  not g14962 (n_8291, n8514);
  and g14963 (n8515, n_8290, n_8291);
  and g14964 (n8516, \A[349] , \A[350] );
  not g14965 (n_8294, \A[350] );
  and g14966 (n8517, \A[349] , n_8294);
  not g14967 (n_8295, \A[349] );
  and g14968 (n8518, n_8295, \A[350] );
  not g14969 (n_8296, n8517);
  not g14970 (n_8297, n8518);
  and g14971 (n8519, n_8296, n_8297);
  not g14972 (n_8299, n8519);
  and g14973 (n8520, \A[351] , n_8299);
  not g14974 (n_8300, n8516);
  not g14975 (n_8301, n8520);
  and g14976 (n8521, n_8300, n_8301);
  not g14977 (n_8302, n8515);
  and g14978 (n8522, n_8302, n8521);
  not g14979 (n_8303, n8521);
  and g14980 (n8523, n8515, n_8303);
  not g14981 (n_8304, n8522);
  not g14982 (n_8305, n8523);
  and g14983 (n8524, n_8304, n_8305);
  and g14984 (n8525, \A[351] , n_8296);
  and g14985 (n8526, n_8297, n8525);
  not g14986 (n_8306, \A[351] );
  and g14987 (n8527, n_8306, n_8299);
  not g14988 (n_8307, n8526);
  not g14989 (n_8308, n8527);
  and g14990 (n8528, n_8307, n_8308);
  and g14991 (n8529, \A[354] , n_8286);
  and g14992 (n8530, n_8287, n8529);
  not g14993 (n_8309, \A[354] );
  and g14994 (n8531, n_8309, n_8289);
  not g14995 (n_8310, n8530);
  not g14996 (n_8311, n8531);
  and g14997 (n8532, n_8310, n_8311);
  not g14998 (n_8312, n8528);
  not g14999 (n_8313, n8532);
  and g15000 (n8533, n_8312, n_8313);
  not g15001 (n_8314, n8524);
  and g15002 (n8534, n_8314, n8533);
  and g15003 (n8535, n_8302, n_8303);
  not g15004 (n_8315, n8534);
  not g15005 (n_8316, n8535);
  and g15006 (n8536, n_8315, n_8316);
  and g15007 (n8537, n_8304, n8533);
  and g15008 (n8538, n_8305, n8537);
  not g15009 (n_8317, n8533);
  and g15010 (n8539, n_8314, n_8317);
  not g15011 (n_8318, n8538);
  not g15012 (n_8319, n8539);
  and g15013 (n8540, n_8318, n_8319);
  not g15014 (n_8320, n8536);
  not g15015 (n_8321, n8540);
  and g15016 (n8541, n_8320, n_8321);
  and g15017 (n8542, n_8312, n8532);
  and g15018 (n8543, n8528, n_8313);
  not g15019 (n_8322, n8542);
  not g15020 (n_8323, n8543);
  and g15021 (n8544, n_8322, n_8323);
  not g15022 (n_8324, n8544);
  and g15023 (n8545, n_8278, n_8324);
  not g15024 (n_8325, n8541);
  and g15025 (n8546, n_8325, n8545);
  not g15026 (n_8326, n8509);
  and g15027 (n8547, n_8326, n8546);
  and g15028 (n8548, n_8320, n_8324);
  not g15029 (n_8327, n8548);
  and g15030 (n8549, n_8321, n_8327);
  not g15031 (n_8328, n8547);
  and g15032 (n8550, n_8328, n8549);
  not g15033 (n_8329, n8549);
  and g15034 (n8551, n8547, n_8329);
  not g15035 (n_8330, n8550);
  not g15036 (n_8331, n8551);
  and g15037 (n8552, n_8330, n_8331);
  not g15038 (n_8332, n8508);
  not g15039 (n_8333, n8552);
  and g15040 (n8553, n_8332, n_8333);
  and g15041 (n8554, n_8328, n_8329);
  not g15046 (n_8334, n8554);
  not g15047 (n_8335, n8558);
  and g15048 (n8559, n_8334, n_8335);
  not g15049 (n_8336, n8559);
  and g15050 (n8560, n8508, n_8336);
  not g15051 (n_8337, n8553);
  not g15052 (n_8338, n8560);
  and g15053 (n8561, n_8337, n_8338);
  and g15054 (n8562, \A[358] , \A[359] );
  not g15055 (n_8341, \A[359] );
  and g15056 (n8563, \A[358] , n_8341);
  not g15057 (n_8342, \A[358] );
  and g15058 (n8564, n_8342, \A[359] );
  not g15059 (n_8343, n8563);
  not g15060 (n_8344, n8564);
  and g15061 (n8565, n_8343, n_8344);
  not g15062 (n_8346, n8565);
  and g15063 (n8566, \A[360] , n_8346);
  not g15064 (n_8347, n8562);
  not g15065 (n_8348, n8566);
  and g15066 (n8567, n_8347, n_8348);
  and g15067 (n8568, \A[355] , \A[356] );
  not g15068 (n_8351, \A[356] );
  and g15069 (n8569, \A[355] , n_8351);
  not g15070 (n_8352, \A[355] );
  and g15071 (n8570, n_8352, \A[356] );
  not g15072 (n_8353, n8569);
  not g15073 (n_8354, n8570);
  and g15074 (n8571, n_8353, n_8354);
  not g15075 (n_8356, n8571);
  and g15076 (n8572, \A[357] , n_8356);
  not g15077 (n_8357, n8568);
  not g15078 (n_8358, n8572);
  and g15079 (n8573, n_8357, n_8358);
  not g15080 (n_8359, n8573);
  and g15081 (n8574, n8567, n_8359);
  not g15082 (n_8360, n8567);
  and g15083 (n8575, n_8360, n8573);
  and g15084 (n8576, \A[357] , n_8353);
  and g15085 (n8577, n_8354, n8576);
  not g15086 (n_8361, \A[357] );
  and g15087 (n8578, n_8361, n_8356);
  not g15088 (n_8362, n8577);
  not g15089 (n_8363, n8578);
  and g15090 (n8579, n_8362, n_8363);
  and g15091 (n8580, \A[360] , n_8343);
  and g15092 (n8581, n_8344, n8580);
  not g15093 (n_8364, \A[360] );
  and g15094 (n8582, n_8364, n_8346);
  not g15095 (n_8365, n8581);
  not g15096 (n_8366, n8582);
  and g15097 (n8583, n_8365, n_8366);
  not g15098 (n_8367, n8579);
  not g15099 (n_8368, n8583);
  and g15100 (n8584, n_8367, n_8368);
  not g15101 (n_8369, n8575);
  and g15102 (n8585, n_8369, n8584);
  not g15103 (n_8370, n8574);
  and g15104 (n8586, n_8370, n8585);
  and g15105 (n8587, n_8370, n_8369);
  not g15106 (n_8371, n8584);
  not g15107 (n_8372, n8587);
  and g15108 (n8588, n_8371, n_8372);
  not g15109 (n_8373, n8586);
  not g15110 (n_8374, n8588);
  and g15111 (n8589, n_8373, n_8374);
  and g15112 (n8590, n_8367, n8583);
  and g15113 (n8591, n8579, n_8368);
  not g15114 (n_8375, n8590);
  not g15115 (n_8376, n8591);
  and g15116 (n8592, n_8375, n_8376);
  and g15117 (n8593, n8584, n_8372);
  and g15118 (n8594, n_8360, n_8359);
  not g15119 (n_8377, n8593);
  not g15120 (n_8378, n8594);
  and g15121 (n8595, n_8377, n_8378);
  not g15122 (n_8379, n8592);
  not g15123 (n_8380, n8595);
  and g15124 (n8596, n_8379, n_8380);
  not g15125 (n_8381, n8589);
  not g15126 (n_8382, n8596);
  and g15127 (n8597, n_8381, n_8382);
  and g15128 (n8598, n_8381, n_8380);
  and g15129 (n8599, \A[364] , \A[365] );
  not g15130 (n_8385, \A[365] );
  and g15131 (n8600, \A[364] , n_8385);
  not g15132 (n_8386, \A[364] );
  and g15133 (n8601, n_8386, \A[365] );
  not g15134 (n_8387, n8600);
  not g15135 (n_8388, n8601);
  and g15136 (n8602, n_8387, n_8388);
  not g15137 (n_8390, n8602);
  and g15138 (n8603, \A[366] , n_8390);
  not g15139 (n_8391, n8599);
  not g15140 (n_8392, n8603);
  and g15141 (n8604, n_8391, n_8392);
  and g15142 (n8605, \A[361] , \A[362] );
  not g15143 (n_8395, \A[362] );
  and g15144 (n8606, \A[361] , n_8395);
  not g15145 (n_8396, \A[361] );
  and g15146 (n8607, n_8396, \A[362] );
  not g15147 (n_8397, n8606);
  not g15148 (n_8398, n8607);
  and g15149 (n8608, n_8397, n_8398);
  not g15150 (n_8400, n8608);
  and g15151 (n8609, \A[363] , n_8400);
  not g15152 (n_8401, n8605);
  not g15153 (n_8402, n8609);
  and g15154 (n8610, n_8401, n_8402);
  not g15155 (n_8403, n8604);
  and g15156 (n8611, n_8403, n8610);
  not g15157 (n_8404, n8610);
  and g15158 (n8612, n8604, n_8404);
  not g15159 (n_8405, n8611);
  not g15160 (n_8406, n8612);
  and g15161 (n8613, n_8405, n_8406);
  and g15162 (n8614, \A[363] , n_8397);
  and g15163 (n8615, n_8398, n8614);
  not g15164 (n_8407, \A[363] );
  and g15165 (n8616, n_8407, n_8400);
  not g15166 (n_8408, n8615);
  not g15167 (n_8409, n8616);
  and g15168 (n8617, n_8408, n_8409);
  and g15169 (n8618, \A[366] , n_8387);
  and g15170 (n8619, n_8388, n8618);
  not g15171 (n_8410, \A[366] );
  and g15172 (n8620, n_8410, n_8390);
  not g15173 (n_8411, n8619);
  not g15174 (n_8412, n8620);
  and g15175 (n8621, n_8411, n_8412);
  not g15176 (n_8413, n8617);
  not g15177 (n_8414, n8621);
  and g15178 (n8622, n_8413, n_8414);
  not g15179 (n_8415, n8613);
  and g15180 (n8623, n_8415, n8622);
  and g15181 (n8624, n_8403, n_8404);
  not g15182 (n_8416, n8623);
  not g15183 (n_8417, n8624);
  and g15184 (n8625, n_8416, n_8417);
  and g15185 (n8626, n_8405, n8622);
  and g15186 (n8627, n_8406, n8626);
  not g15187 (n_8418, n8622);
  and g15188 (n8628, n_8415, n_8418);
  not g15189 (n_8419, n8627);
  not g15190 (n_8420, n8628);
  and g15191 (n8629, n_8419, n_8420);
  not g15192 (n_8421, n8625);
  not g15193 (n_8422, n8629);
  and g15194 (n8630, n_8421, n_8422);
  and g15195 (n8631, n_8413, n8621);
  and g15196 (n8632, n8617, n_8414);
  not g15197 (n_8423, n8631);
  not g15198 (n_8424, n8632);
  and g15199 (n8633, n_8423, n_8424);
  not g15200 (n_8425, n8633);
  and g15201 (n8634, n_8379, n_8425);
  not g15202 (n_8426, n8630);
  and g15203 (n8635, n_8426, n8634);
  not g15204 (n_8427, n8598);
  and g15205 (n8636, n_8427, n8635);
  and g15206 (n8637, n_8421, n_8425);
  not g15207 (n_8428, n8637);
  and g15208 (n8638, n_8422, n_8428);
  not g15209 (n_8429, n8636);
  not g15210 (n_8430, n8638);
  and g15211 (n8639, n_8429, n_8430);
  not g15216 (n_8431, n8639);
  not g15217 (n_8432, n8643);
  and g15218 (n8644, n_8431, n_8432);
  not g15219 (n_8433, n8644);
  and g15220 (n8645, n8597, n_8433);
  and g15221 (n8646, n_8429, n8638);
  and g15222 (n8647, n8636, n_8430);
  not g15223 (n_8434, n8646);
  not g15224 (n_8435, n8647);
  and g15225 (n8648, n_8434, n_8435);
  not g15226 (n_8436, n8597);
  not g15227 (n_8437, n8648);
  and g15228 (n8649, n_8436, n_8437);
  and g15229 (n8650, n_8426, n_8425);
  and g15230 (n8651, n_8379, n_8427);
  not g15231 (n_8438, n8650);
  and g15232 (n8652, n_8438, n8651);
  not g15233 (n_8439, n8651);
  and g15234 (n8653, n8650, n_8439);
  not g15235 (n_8440, n8652);
  not g15236 (n_8441, n8653);
  and g15237 (n8654, n_8440, n_8441);
  and g15238 (n8655, n_8325, n_8324);
  and g15239 (n8656, n_8278, n_8326);
  not g15240 (n_8442, n8655);
  and g15241 (n8657, n_8442, n8656);
  not g15242 (n_8443, n8656);
  and g15243 (n8658, n8655, n_8443);
  not g15244 (n_8444, n8657);
  not g15245 (n_8445, n8658);
  and g15246 (n8659, n_8444, n_8445);
  not g15247 (n_8446, n8654);
  not g15248 (n_8447, n8659);
  and g15249 (n8660, n_8446, n_8447);
  not g15250 (n_8448, n8649);
  not g15251 (n_8449, n8660);
  and g15252 (n8661, n_8448, n_8449);
  not g15253 (n_8450, n8645);
  and g15254 (n8662, n_8450, n8661);
  and g15255 (n8663, n_8450, n_8448);
  not g15256 (n_8451, n8663);
  and g15257 (n8664, n8660, n_8451);
  not g15258 (n_8452, n8662);
  not g15259 (n_8453, n8664);
  and g15260 (n8665, n_8452, n_8453);
  not g15261 (n_8454, n8561);
  not g15262 (n_8455, n8665);
  and g15263 (n8666, n_8454, n_8455);
  and g15264 (n8667, n_8448, n8660);
  and g15265 (n8668, n_8450, n8667);
  and g15266 (n8669, n_8449, n_8451);
  not g15267 (n_8456, n8668);
  not g15268 (n_8457, n8669);
  and g15269 (n8670, n_8456, n_8457);
  not g15270 (n_8458, n8670);
  and g15271 (n8671, n8561, n_8458);
  and g15272 (n8672, n_8446, n8659);
  and g15273 (n8673, n8654, n_8447);
  not g15274 (n_8459, n8672);
  not g15275 (n_8460, n8673);
  and g15276 (n8674, n_8459, n_8460);
  and g15277 (n8675, n_8210, n8440);
  and g15278 (n8676, n8365, n_8211);
  not g15279 (n_8461, n8675);
  not g15280 (n_8462, n8676);
  and g15281 (n8677, n_8461, n_8462);
  not g15282 (n_8463, n8674);
  not g15283 (n_8464, n8677);
  and g15284 (n8678, n_8463, n_8464);
  not g15285 (n_8465, n8671);
  not g15286 (n_8466, n8678);
  and g15287 (n8679, n_8465, n_8466);
  not g15288 (n_8467, n8666);
  and g15289 (n8680, n_8467, n8679);
  and g15290 (n8681, n_8467, n_8465);
  not g15291 (n_8468, n8681);
  and g15292 (n8682, n8678, n_8468);
  not g15293 (n_8469, n8680);
  not g15294 (n_8470, n8682);
  and g15295 (n8683, n_8469, n_8470);
  not g15296 (n_8471, n8472);
  not g15297 (n_8472, n8683);
  and g15298 (n8684, n_8471, n_8472);
  and g15299 (n8685, n_8465, n8678);
  and g15300 (n8686, n_8467, n8685);
  and g15301 (n8687, n_8466, n_8468);
  not g15302 (n_8473, n8686);
  not g15303 (n_8474, n8687);
  and g15304 (n8688, n_8473, n_8474);
  not g15305 (n_8475, n8688);
  and g15306 (n8689, n8472, n_8475);
  and g15307 (n8690, n_8463, n8677);
  and g15308 (n8691, n8674, n_8464);
  not g15309 (n_8476, n8690);
  not g15310 (n_8477, n8691);
  and g15311 (n8692, n_8476, n_8477);
  not g15312 (n_8479, \A[313] );
  and g15313 (n8693, n_8479, \A[314] );
  not g15314 (n_8481, \A[314] );
  and g15315 (n8694, \A[313] , n_8481);
  not g15316 (n_8483, n8694);
  and g15317 (n8695, \A[315] , n_8483);
  not g15318 (n_8484, n8693);
  and g15319 (n8696, n_8484, n8695);
  and g15320 (n8697, n_8484, n_8483);
  not g15321 (n_8485, \A[315] );
  not g15322 (n_8486, n8697);
  and g15323 (n8698, n_8485, n_8486);
  not g15324 (n_8487, n8696);
  not g15325 (n_8488, n8698);
  and g15326 (n8699, n_8487, n_8488);
  not g15327 (n_8490, \A[316] );
  and g15328 (n8700, n_8490, \A[317] );
  not g15329 (n_8492, \A[317] );
  and g15330 (n8701, \A[316] , n_8492);
  not g15331 (n_8494, n8701);
  and g15332 (n8702, \A[318] , n_8494);
  not g15333 (n_8495, n8700);
  and g15334 (n8703, n_8495, n8702);
  and g15335 (n8704, n_8495, n_8494);
  not g15336 (n_8496, \A[318] );
  not g15337 (n_8497, n8704);
  and g15338 (n8705, n_8496, n_8497);
  not g15339 (n_8498, n8703);
  not g15340 (n_8499, n8705);
  and g15341 (n8706, n_8498, n_8499);
  not g15342 (n_8500, n8699);
  and g15343 (n8707, n_8500, n8706);
  not g15344 (n_8501, n8706);
  and g15345 (n8708, n8699, n_8501);
  not g15346 (n_8502, n8707);
  not g15347 (n_8503, n8708);
  and g15348 (n8709, n_8502, n_8503);
  and g15349 (n8710, \A[316] , \A[317] );
  and g15350 (n8711, \A[318] , n_8497);
  not g15351 (n_8504, n8710);
  not g15352 (n_8505, n8711);
  and g15353 (n8712, n_8504, n_8505);
  and g15354 (n8713, \A[313] , \A[314] );
  and g15355 (n8714, \A[315] , n_8486);
  not g15356 (n_8506, n8713);
  not g15357 (n_8507, n8714);
  and g15358 (n8715, n_8506, n_8507);
  not g15359 (n_8508, n8712);
  and g15360 (n8716, n_8508, n8715);
  not g15361 (n_8509, n8715);
  and g15362 (n8717, n8712, n_8509);
  not g15363 (n_8510, n8716);
  not g15364 (n_8511, n8717);
  and g15365 (n8718, n_8510, n_8511);
  and g15366 (n8719, n_8500, n_8501);
  not g15367 (n_8512, n8718);
  and g15368 (n8720, n_8512, n8719);
  and g15369 (n8721, n_8508, n_8509);
  not g15370 (n_8513, n8720);
  not g15371 (n_8514, n8721);
  and g15372 (n8722, n_8513, n_8514);
  and g15373 (n8723, n_8510, n8719);
  and g15374 (n8724, n_8511, n8723);
  not g15375 (n_8515, n8719);
  and g15376 (n8725, n_8512, n_8515);
  not g15377 (n_8516, n8724);
  not g15378 (n_8517, n8725);
  and g15379 (n8726, n_8516, n_8517);
  not g15380 (n_8518, n8722);
  not g15381 (n_8519, n8726);
  and g15382 (n8727, n_8518, n_8519);
  not g15383 (n_8520, n8709);
  not g15384 (n_8521, n8727);
  and g15385 (n8728, n_8520, n_8521);
  not g15386 (n_8523, \A[307] );
  and g15387 (n8729, n_8523, \A[308] );
  not g15388 (n_8525, \A[308] );
  and g15389 (n8730, \A[307] , n_8525);
  not g15390 (n_8527, n8730);
  and g15391 (n8731, \A[309] , n_8527);
  not g15392 (n_8528, n8729);
  and g15393 (n8732, n_8528, n8731);
  and g15394 (n8733, n_8528, n_8527);
  not g15395 (n_8529, \A[309] );
  not g15396 (n_8530, n8733);
  and g15397 (n8734, n_8529, n_8530);
  not g15398 (n_8531, n8732);
  not g15399 (n_8532, n8734);
  and g15400 (n8735, n_8531, n_8532);
  not g15401 (n_8534, \A[310] );
  and g15402 (n8736, n_8534, \A[311] );
  not g15403 (n_8536, \A[311] );
  and g15404 (n8737, \A[310] , n_8536);
  not g15405 (n_8538, n8737);
  and g15406 (n8738, \A[312] , n_8538);
  not g15407 (n_8539, n8736);
  and g15408 (n8739, n_8539, n8738);
  and g15409 (n8740, n_8539, n_8538);
  not g15410 (n_8540, \A[312] );
  not g15411 (n_8541, n8740);
  and g15412 (n8741, n_8540, n_8541);
  not g15413 (n_8542, n8739);
  not g15414 (n_8543, n8741);
  and g15415 (n8742, n_8542, n_8543);
  not g15416 (n_8544, n8735);
  and g15417 (n8743, n_8544, n8742);
  not g15418 (n_8545, n8742);
  and g15419 (n8744, n8735, n_8545);
  not g15420 (n_8546, n8743);
  not g15421 (n_8547, n8744);
  and g15422 (n8745, n_8546, n_8547);
  and g15423 (n8746, \A[310] , \A[311] );
  and g15424 (n8747, \A[312] , n_8541);
  not g15425 (n_8548, n8746);
  not g15426 (n_8549, n8747);
  and g15427 (n8748, n_8548, n_8549);
  and g15428 (n8749, \A[307] , \A[308] );
  and g15429 (n8750, \A[309] , n_8530);
  not g15430 (n_8550, n8749);
  not g15431 (n_8551, n8750);
  and g15432 (n8751, n_8550, n_8551);
  not g15433 (n_8552, n8748);
  and g15434 (n8752, n_8552, n8751);
  not g15435 (n_8553, n8751);
  and g15436 (n8753, n8748, n_8553);
  not g15437 (n_8554, n8752);
  not g15438 (n_8555, n8753);
  and g15439 (n8754, n_8554, n_8555);
  and g15440 (n8755, n_8544, n_8545);
  not g15441 (n_8556, n8754);
  and g15442 (n8756, n_8556, n8755);
  and g15443 (n8757, n_8552, n_8553);
  not g15444 (n_8557, n8756);
  not g15445 (n_8558, n8757);
  and g15446 (n8758, n_8557, n_8558);
  and g15447 (n8759, n_8554, n8755);
  and g15448 (n8760, n_8555, n8759);
  not g15449 (n_8559, n8755);
  and g15450 (n8761, n_8556, n_8559);
  not g15451 (n_8560, n8760);
  not g15452 (n_8561, n8761);
  and g15453 (n8762, n_8560, n_8561);
  not g15454 (n_8562, n8758);
  not g15455 (n_8563, n8762);
  and g15456 (n8763, n_8562, n_8563);
  not g15457 (n_8564, n8745);
  not g15458 (n_8565, n8763);
  and g15459 (n8764, n_8564, n_8565);
  not g15460 (n_8566, n8728);
  and g15461 (n8765, n_8566, n8764);
  not g15462 (n_8567, n8764);
  and g15463 (n8766, n8728, n_8567);
  not g15464 (n_8568, n8765);
  not g15465 (n_8569, n8766);
  and g15466 (n8767, n_8568, n_8569);
  not g15467 (n_8571, \A[301] );
  and g15468 (n8768, n_8571, \A[302] );
  not g15469 (n_8573, \A[302] );
  and g15470 (n8769, \A[301] , n_8573);
  not g15471 (n_8575, n8769);
  and g15472 (n8770, \A[303] , n_8575);
  not g15473 (n_8576, n8768);
  and g15474 (n8771, n_8576, n8770);
  and g15475 (n8772, n_8576, n_8575);
  not g15476 (n_8577, \A[303] );
  not g15477 (n_8578, n8772);
  and g15478 (n8773, n_8577, n_8578);
  not g15479 (n_8579, n8771);
  not g15480 (n_8580, n8773);
  and g15481 (n8774, n_8579, n_8580);
  not g15482 (n_8582, \A[304] );
  and g15483 (n8775, n_8582, \A[305] );
  not g15484 (n_8584, \A[305] );
  and g15485 (n8776, \A[304] , n_8584);
  not g15486 (n_8586, n8776);
  and g15487 (n8777, \A[306] , n_8586);
  not g15488 (n_8587, n8775);
  and g15489 (n8778, n_8587, n8777);
  and g15490 (n8779, n_8587, n_8586);
  not g15491 (n_8588, \A[306] );
  not g15492 (n_8589, n8779);
  and g15493 (n8780, n_8588, n_8589);
  not g15494 (n_8590, n8778);
  not g15495 (n_8591, n8780);
  and g15496 (n8781, n_8590, n_8591);
  not g15497 (n_8592, n8774);
  and g15498 (n8782, n_8592, n8781);
  not g15499 (n_8593, n8781);
  and g15500 (n8783, n8774, n_8593);
  not g15501 (n_8594, n8782);
  not g15502 (n_8595, n8783);
  and g15503 (n8784, n_8594, n_8595);
  and g15504 (n8785, \A[304] , \A[305] );
  and g15505 (n8786, \A[306] , n_8589);
  not g15506 (n_8596, n8785);
  not g15507 (n_8597, n8786);
  and g15508 (n8787, n_8596, n_8597);
  and g15509 (n8788, \A[301] , \A[302] );
  and g15510 (n8789, \A[303] , n_8578);
  not g15511 (n_8598, n8788);
  not g15512 (n_8599, n8789);
  and g15513 (n8790, n_8598, n_8599);
  not g15514 (n_8600, n8787);
  and g15515 (n8791, n_8600, n8790);
  not g15516 (n_8601, n8790);
  and g15517 (n8792, n8787, n_8601);
  not g15518 (n_8602, n8791);
  not g15519 (n_8603, n8792);
  and g15520 (n8793, n_8602, n_8603);
  and g15521 (n8794, n_8592, n_8593);
  not g15522 (n_8604, n8793);
  and g15523 (n8795, n_8604, n8794);
  and g15524 (n8796, n_8600, n_8601);
  not g15525 (n_8605, n8795);
  not g15526 (n_8606, n8796);
  and g15527 (n8797, n_8605, n_8606);
  and g15528 (n8798, n_8602, n8794);
  and g15529 (n8799, n_8603, n8798);
  not g15530 (n_8607, n8794);
  and g15531 (n8800, n_8604, n_8607);
  not g15532 (n_8608, n8799);
  not g15533 (n_8609, n8800);
  and g15534 (n8801, n_8608, n_8609);
  not g15535 (n_8610, n8797);
  not g15536 (n_8611, n8801);
  and g15537 (n8802, n_8610, n_8611);
  not g15538 (n_8612, n8784);
  not g15539 (n_8613, n8802);
  and g15540 (n8803, n_8612, n_8613);
  not g15541 (n_8615, \A[295] );
  and g15542 (n8804, n_8615, \A[296] );
  not g15543 (n_8617, \A[296] );
  and g15544 (n8805, \A[295] , n_8617);
  not g15545 (n_8619, n8805);
  and g15546 (n8806, \A[297] , n_8619);
  not g15547 (n_8620, n8804);
  and g15548 (n8807, n_8620, n8806);
  and g15549 (n8808, n_8620, n_8619);
  not g15550 (n_8621, \A[297] );
  not g15551 (n_8622, n8808);
  and g15552 (n8809, n_8621, n_8622);
  not g15553 (n_8623, n8807);
  not g15554 (n_8624, n8809);
  and g15555 (n8810, n_8623, n_8624);
  not g15556 (n_8626, \A[298] );
  and g15557 (n8811, n_8626, \A[299] );
  not g15558 (n_8628, \A[299] );
  and g15559 (n8812, \A[298] , n_8628);
  not g15560 (n_8630, n8812);
  and g15561 (n8813, \A[300] , n_8630);
  not g15562 (n_8631, n8811);
  and g15563 (n8814, n_8631, n8813);
  and g15564 (n8815, n_8631, n_8630);
  not g15565 (n_8632, \A[300] );
  not g15566 (n_8633, n8815);
  and g15567 (n8816, n_8632, n_8633);
  not g15568 (n_8634, n8814);
  not g15569 (n_8635, n8816);
  and g15570 (n8817, n_8634, n_8635);
  not g15571 (n_8636, n8810);
  and g15572 (n8818, n_8636, n8817);
  not g15573 (n_8637, n8817);
  and g15574 (n8819, n8810, n_8637);
  not g15575 (n_8638, n8818);
  not g15576 (n_8639, n8819);
  and g15577 (n8820, n_8638, n_8639);
  and g15578 (n8821, \A[298] , \A[299] );
  and g15579 (n8822, \A[300] , n_8633);
  not g15580 (n_8640, n8821);
  not g15581 (n_8641, n8822);
  and g15582 (n8823, n_8640, n_8641);
  and g15583 (n8824, \A[295] , \A[296] );
  and g15584 (n8825, \A[297] , n_8622);
  not g15585 (n_8642, n8824);
  not g15586 (n_8643, n8825);
  and g15587 (n8826, n_8642, n_8643);
  not g15588 (n_8644, n8823);
  and g15589 (n8827, n_8644, n8826);
  not g15590 (n_8645, n8826);
  and g15591 (n8828, n8823, n_8645);
  not g15592 (n_8646, n8827);
  not g15593 (n_8647, n8828);
  and g15594 (n8829, n_8646, n_8647);
  and g15595 (n8830, n_8636, n_8637);
  not g15596 (n_8648, n8829);
  and g15597 (n8831, n_8648, n8830);
  and g15598 (n8832, n_8644, n_8645);
  not g15599 (n_8649, n8831);
  not g15600 (n_8650, n8832);
  and g15601 (n8833, n_8649, n_8650);
  and g15602 (n8834, n_8646, n8830);
  and g15603 (n8835, n_8647, n8834);
  not g15604 (n_8651, n8830);
  and g15605 (n8836, n_8648, n_8651);
  not g15606 (n_8652, n8835);
  not g15607 (n_8653, n8836);
  and g15608 (n8837, n_8652, n_8653);
  not g15609 (n_8654, n8833);
  not g15610 (n_8655, n8837);
  and g15611 (n8838, n_8654, n_8655);
  not g15612 (n_8656, n8820);
  not g15613 (n_8657, n8838);
  and g15614 (n8839, n_8656, n_8657);
  not g15615 (n_8658, n8803);
  and g15616 (n8840, n_8658, n8839);
  not g15617 (n_8659, n8839);
  and g15618 (n8841, n8803, n_8659);
  not g15619 (n_8660, n8840);
  not g15620 (n_8661, n8841);
  and g15621 (n8842, n_8660, n_8661);
  not g15622 (n_8662, n8767);
  and g15623 (n8843, n_8662, n8842);
  not g15624 (n_8663, n8842);
  and g15625 (n8844, n8767, n_8663);
  not g15626 (n_8664, n8843);
  not g15627 (n_8665, n8844);
  and g15628 (n8845, n_8664, n_8665);
  not g15629 (n_8667, \A[289] );
  and g15630 (n8846, n_8667, \A[290] );
  not g15631 (n_8669, \A[290] );
  and g15632 (n8847, \A[289] , n_8669);
  not g15633 (n_8671, n8847);
  and g15634 (n8848, \A[291] , n_8671);
  not g15635 (n_8672, n8846);
  and g15636 (n8849, n_8672, n8848);
  and g15637 (n8850, n_8672, n_8671);
  not g15638 (n_8673, \A[291] );
  not g15639 (n_8674, n8850);
  and g15640 (n8851, n_8673, n_8674);
  not g15641 (n_8675, n8849);
  not g15642 (n_8676, n8851);
  and g15643 (n8852, n_8675, n_8676);
  not g15644 (n_8678, \A[292] );
  and g15645 (n8853, n_8678, \A[293] );
  not g15646 (n_8680, \A[293] );
  and g15647 (n8854, \A[292] , n_8680);
  not g15648 (n_8682, n8854);
  and g15649 (n8855, \A[294] , n_8682);
  not g15650 (n_8683, n8853);
  and g15651 (n8856, n_8683, n8855);
  and g15652 (n8857, n_8683, n_8682);
  not g15653 (n_8684, \A[294] );
  not g15654 (n_8685, n8857);
  and g15655 (n8858, n_8684, n_8685);
  not g15656 (n_8686, n8856);
  not g15657 (n_8687, n8858);
  and g15658 (n8859, n_8686, n_8687);
  not g15659 (n_8688, n8852);
  and g15660 (n8860, n_8688, n8859);
  not g15661 (n_8689, n8859);
  and g15662 (n8861, n8852, n_8689);
  not g15663 (n_8690, n8860);
  not g15664 (n_8691, n8861);
  and g15665 (n8862, n_8690, n_8691);
  and g15666 (n8863, \A[292] , \A[293] );
  and g15667 (n8864, \A[294] , n_8685);
  not g15668 (n_8692, n8863);
  not g15669 (n_8693, n8864);
  and g15670 (n8865, n_8692, n_8693);
  and g15671 (n8866, \A[289] , \A[290] );
  and g15672 (n8867, \A[291] , n_8674);
  not g15673 (n_8694, n8866);
  not g15674 (n_8695, n8867);
  and g15675 (n8868, n_8694, n_8695);
  not g15676 (n_8696, n8865);
  and g15677 (n8869, n_8696, n8868);
  not g15678 (n_8697, n8868);
  and g15679 (n8870, n8865, n_8697);
  not g15680 (n_8698, n8869);
  not g15681 (n_8699, n8870);
  and g15682 (n8871, n_8698, n_8699);
  and g15683 (n8872, n_8688, n_8689);
  not g15684 (n_8700, n8871);
  and g15685 (n8873, n_8700, n8872);
  and g15686 (n8874, n_8696, n_8697);
  not g15687 (n_8701, n8873);
  not g15688 (n_8702, n8874);
  and g15689 (n8875, n_8701, n_8702);
  and g15690 (n8876, n_8698, n8872);
  and g15691 (n8877, n_8699, n8876);
  not g15692 (n_8703, n8872);
  and g15693 (n8878, n_8700, n_8703);
  not g15694 (n_8704, n8877);
  not g15695 (n_8705, n8878);
  and g15696 (n8879, n_8704, n_8705);
  not g15697 (n_8706, n8875);
  not g15698 (n_8707, n8879);
  and g15699 (n8880, n_8706, n_8707);
  not g15700 (n_8708, n8862);
  not g15701 (n_8709, n8880);
  and g15702 (n8881, n_8708, n_8709);
  not g15703 (n_8711, \A[283] );
  and g15704 (n8882, n_8711, \A[284] );
  not g15705 (n_8713, \A[284] );
  and g15706 (n8883, \A[283] , n_8713);
  not g15707 (n_8715, n8883);
  and g15708 (n8884, \A[285] , n_8715);
  not g15709 (n_8716, n8882);
  and g15710 (n8885, n_8716, n8884);
  and g15711 (n8886, n_8716, n_8715);
  not g15712 (n_8717, \A[285] );
  not g15713 (n_8718, n8886);
  and g15714 (n8887, n_8717, n_8718);
  not g15715 (n_8719, n8885);
  not g15716 (n_8720, n8887);
  and g15717 (n8888, n_8719, n_8720);
  not g15718 (n_8722, \A[286] );
  and g15719 (n8889, n_8722, \A[287] );
  not g15720 (n_8724, \A[287] );
  and g15721 (n8890, \A[286] , n_8724);
  not g15722 (n_8726, n8890);
  and g15723 (n8891, \A[288] , n_8726);
  not g15724 (n_8727, n8889);
  and g15725 (n8892, n_8727, n8891);
  and g15726 (n8893, n_8727, n_8726);
  not g15727 (n_8728, \A[288] );
  not g15728 (n_8729, n8893);
  and g15729 (n8894, n_8728, n_8729);
  not g15730 (n_8730, n8892);
  not g15731 (n_8731, n8894);
  and g15732 (n8895, n_8730, n_8731);
  not g15733 (n_8732, n8888);
  and g15734 (n8896, n_8732, n8895);
  not g15735 (n_8733, n8895);
  and g15736 (n8897, n8888, n_8733);
  not g15737 (n_8734, n8896);
  not g15738 (n_8735, n8897);
  and g15739 (n8898, n_8734, n_8735);
  and g15740 (n8899, \A[286] , \A[287] );
  and g15741 (n8900, \A[288] , n_8729);
  not g15742 (n_8736, n8899);
  not g15743 (n_8737, n8900);
  and g15744 (n8901, n_8736, n_8737);
  and g15745 (n8902, \A[283] , \A[284] );
  and g15746 (n8903, \A[285] , n_8718);
  not g15747 (n_8738, n8902);
  not g15748 (n_8739, n8903);
  and g15749 (n8904, n_8738, n_8739);
  not g15750 (n_8740, n8901);
  and g15751 (n8905, n_8740, n8904);
  not g15752 (n_8741, n8904);
  and g15753 (n8906, n8901, n_8741);
  not g15754 (n_8742, n8905);
  not g15755 (n_8743, n8906);
  and g15756 (n8907, n_8742, n_8743);
  and g15757 (n8908, n_8732, n_8733);
  not g15758 (n_8744, n8907);
  and g15759 (n8909, n_8744, n8908);
  and g15760 (n8910, n_8740, n_8741);
  not g15761 (n_8745, n8909);
  not g15762 (n_8746, n8910);
  and g15763 (n8911, n_8745, n_8746);
  and g15764 (n8912, n_8742, n8908);
  and g15765 (n8913, n_8743, n8912);
  not g15766 (n_8747, n8908);
  and g15767 (n8914, n_8744, n_8747);
  not g15768 (n_8748, n8913);
  not g15769 (n_8749, n8914);
  and g15770 (n8915, n_8748, n_8749);
  not g15771 (n_8750, n8911);
  not g15772 (n_8751, n8915);
  and g15773 (n8916, n_8750, n_8751);
  not g15774 (n_8752, n8898);
  not g15775 (n_8753, n8916);
  and g15776 (n8917, n_8752, n_8753);
  not g15777 (n_8754, n8881);
  and g15778 (n8918, n_8754, n8917);
  not g15779 (n_8755, n8917);
  and g15780 (n8919, n8881, n_8755);
  not g15781 (n_8756, n8918);
  not g15782 (n_8757, n8919);
  and g15783 (n8920, n_8756, n_8757);
  not g15784 (n_8759, \A[277] );
  and g15785 (n8921, n_8759, \A[278] );
  not g15786 (n_8761, \A[278] );
  and g15787 (n8922, \A[277] , n_8761);
  not g15788 (n_8763, n8922);
  and g15789 (n8923, \A[279] , n_8763);
  not g15790 (n_8764, n8921);
  and g15791 (n8924, n_8764, n8923);
  and g15792 (n8925, n_8764, n_8763);
  not g15793 (n_8765, \A[279] );
  not g15794 (n_8766, n8925);
  and g15795 (n8926, n_8765, n_8766);
  not g15796 (n_8767, n8924);
  not g15797 (n_8768, n8926);
  and g15798 (n8927, n_8767, n_8768);
  not g15799 (n_8770, \A[280] );
  and g15800 (n8928, n_8770, \A[281] );
  not g15801 (n_8772, \A[281] );
  and g15802 (n8929, \A[280] , n_8772);
  not g15803 (n_8774, n8929);
  and g15804 (n8930, \A[282] , n_8774);
  not g15805 (n_8775, n8928);
  and g15806 (n8931, n_8775, n8930);
  and g15807 (n8932, n_8775, n_8774);
  not g15808 (n_8776, \A[282] );
  not g15809 (n_8777, n8932);
  and g15810 (n8933, n_8776, n_8777);
  not g15811 (n_8778, n8931);
  not g15812 (n_8779, n8933);
  and g15813 (n8934, n_8778, n_8779);
  not g15814 (n_8780, n8927);
  and g15815 (n8935, n_8780, n8934);
  not g15816 (n_8781, n8934);
  and g15817 (n8936, n8927, n_8781);
  not g15818 (n_8782, n8935);
  not g15819 (n_8783, n8936);
  and g15820 (n8937, n_8782, n_8783);
  and g15821 (n8938, \A[280] , \A[281] );
  and g15822 (n8939, \A[282] , n_8777);
  not g15823 (n_8784, n8938);
  not g15824 (n_8785, n8939);
  and g15825 (n8940, n_8784, n_8785);
  and g15826 (n8941, \A[277] , \A[278] );
  and g15827 (n8942, \A[279] , n_8766);
  not g15828 (n_8786, n8941);
  not g15829 (n_8787, n8942);
  and g15830 (n8943, n_8786, n_8787);
  not g15831 (n_8788, n8940);
  and g15832 (n8944, n_8788, n8943);
  not g15833 (n_8789, n8943);
  and g15834 (n8945, n8940, n_8789);
  not g15835 (n_8790, n8944);
  not g15836 (n_8791, n8945);
  and g15837 (n8946, n_8790, n_8791);
  and g15838 (n8947, n_8780, n_8781);
  not g15839 (n_8792, n8946);
  and g15840 (n8948, n_8792, n8947);
  and g15841 (n8949, n_8788, n_8789);
  not g15842 (n_8793, n8948);
  not g15843 (n_8794, n8949);
  and g15844 (n8950, n_8793, n_8794);
  and g15845 (n8951, n_8790, n8947);
  and g15846 (n8952, n_8791, n8951);
  not g15847 (n_8795, n8947);
  and g15848 (n8953, n_8792, n_8795);
  not g15849 (n_8796, n8952);
  not g15850 (n_8797, n8953);
  and g15851 (n8954, n_8796, n_8797);
  not g15852 (n_8798, n8950);
  not g15853 (n_8799, n8954);
  and g15854 (n8955, n_8798, n_8799);
  not g15855 (n_8800, n8937);
  not g15856 (n_8801, n8955);
  and g15857 (n8956, n_8800, n_8801);
  not g15858 (n_8803, \A[271] );
  and g15859 (n8957, n_8803, \A[272] );
  not g15860 (n_8805, \A[272] );
  and g15861 (n8958, \A[271] , n_8805);
  not g15862 (n_8807, n8958);
  and g15863 (n8959, \A[273] , n_8807);
  not g15864 (n_8808, n8957);
  and g15865 (n8960, n_8808, n8959);
  and g15866 (n8961, n_8808, n_8807);
  not g15867 (n_8809, \A[273] );
  not g15868 (n_8810, n8961);
  and g15869 (n8962, n_8809, n_8810);
  not g15870 (n_8811, n8960);
  not g15871 (n_8812, n8962);
  and g15872 (n8963, n_8811, n_8812);
  not g15873 (n_8814, \A[274] );
  and g15874 (n8964, n_8814, \A[275] );
  not g15875 (n_8816, \A[275] );
  and g15876 (n8965, \A[274] , n_8816);
  not g15877 (n_8818, n8965);
  and g15878 (n8966, \A[276] , n_8818);
  not g15879 (n_8819, n8964);
  and g15880 (n8967, n_8819, n8966);
  and g15881 (n8968, n_8819, n_8818);
  not g15882 (n_8820, \A[276] );
  not g15883 (n_8821, n8968);
  and g15884 (n8969, n_8820, n_8821);
  not g15885 (n_8822, n8967);
  not g15886 (n_8823, n8969);
  and g15887 (n8970, n_8822, n_8823);
  not g15888 (n_8824, n8963);
  and g15889 (n8971, n_8824, n8970);
  not g15890 (n_8825, n8970);
  and g15891 (n8972, n8963, n_8825);
  not g15892 (n_8826, n8971);
  not g15893 (n_8827, n8972);
  and g15894 (n8973, n_8826, n_8827);
  and g15895 (n8974, \A[274] , \A[275] );
  and g15896 (n8975, \A[276] , n_8821);
  not g15897 (n_8828, n8974);
  not g15898 (n_8829, n8975);
  and g15899 (n8976, n_8828, n_8829);
  and g15900 (n8977, \A[271] , \A[272] );
  and g15901 (n8978, \A[273] , n_8810);
  not g15902 (n_8830, n8977);
  not g15903 (n_8831, n8978);
  and g15904 (n8979, n_8830, n_8831);
  not g15905 (n_8832, n8976);
  and g15906 (n8980, n_8832, n8979);
  not g15907 (n_8833, n8979);
  and g15908 (n8981, n8976, n_8833);
  not g15909 (n_8834, n8980);
  not g15910 (n_8835, n8981);
  and g15911 (n8982, n_8834, n_8835);
  and g15912 (n8983, n_8824, n_8825);
  not g15913 (n_8836, n8982);
  and g15914 (n8984, n_8836, n8983);
  and g15915 (n8985, n_8832, n_8833);
  not g15916 (n_8837, n8984);
  not g15917 (n_8838, n8985);
  and g15918 (n8986, n_8837, n_8838);
  and g15919 (n8987, n_8834, n8983);
  and g15920 (n8988, n_8835, n8987);
  not g15921 (n_8839, n8983);
  and g15922 (n8989, n_8836, n_8839);
  not g15923 (n_8840, n8988);
  not g15924 (n_8841, n8989);
  and g15925 (n8990, n_8840, n_8841);
  not g15926 (n_8842, n8986);
  not g15927 (n_8843, n8990);
  and g15928 (n8991, n_8842, n_8843);
  not g15929 (n_8844, n8973);
  not g15930 (n_8845, n8991);
  and g15931 (n8992, n_8844, n_8845);
  not g15932 (n_8846, n8956);
  and g15933 (n8993, n_8846, n8992);
  not g15934 (n_8847, n8992);
  and g15935 (n8994, n8956, n_8847);
  not g15936 (n_8848, n8993);
  not g15937 (n_8849, n8994);
  and g15938 (n8995, n_8848, n_8849);
  not g15939 (n_8850, n8920);
  and g15940 (n8996, n_8850, n8995);
  not g15941 (n_8851, n8995);
  and g15942 (n8997, n8920, n_8851);
  not g15943 (n_8852, n8996);
  not g15944 (n_8853, n8997);
  and g15945 (n8998, n_8852, n_8853);
  not g15946 (n_8854, n8845);
  and g15947 (n8999, n_8854, n8998);
  not g15948 (n_8855, n8998);
  and g15949 (n9000, n8845, n_8855);
  not g15950 (n_8856, n8999);
  not g15951 (n_8857, n9000);
  and g15952 (n9001, n_8856, n_8857);
  not g15953 (n_8858, n8692);
  not g15954 (n_8859, n9001);
  and g15955 (n9002, n_8858, n_8859);
  not g15956 (n_8860, n8689);
  and g15957 (n9003, n_8860, n9002);
  not g15958 (n_8861, n8684);
  and g15959 (n9004, n_8861, n9003);
  and g15960 (n9005, n_8861, n_8860);
  not g15961 (n_8862, n9002);
  not g15962 (n_8863, n9005);
  and g15963 (n9006, n_8862, n_8863);
  not g15964 (n_8864, n9004);
  not g15965 (n_8865, n9006);
  and g15966 (n9007, n_8864, n_8865);
  and g15967 (n9008, n_8656, n_8654);
  not g15968 (n_8866, n9008);
  and g15969 (n9009, n_8655, n_8866);
  and g15970 (n9010, n_8612, n_8656);
  and g15971 (n9011, n_8613, n9010);
  and g15972 (n9012, n_8657, n9011);
  and g15973 (n9013, n_8612, n_8610);
  not g15974 (n_8867, n9013);
  and g15975 (n9014, n_8611, n_8867);
  not g15976 (n_8868, n9012);
  and g15977 (n9015, n_8868, n9014);
  not g15978 (n_8869, n9014);
  and g15979 (n9016, n9012, n_8869);
  not g15980 (n_8870, n9015);
  not g15981 (n_8871, n9016);
  and g15982 (n9017, n_8870, n_8871);
  not g15983 (n_8872, n9009);
  not g15984 (n_8873, n9017);
  and g15985 (n9018, n_8872, n_8873);
  and g15986 (n9019, n_8868, n_8869);
  not g15991 (n_8874, n9019);
  not g15992 (n_8875, n9023);
  and g15993 (n9024, n_8874, n_8875);
  not g15994 (n_8876, n9024);
  and g15995 (n9025, n9009, n_8876);
  not g15996 (n_8877, n9018);
  not g15997 (n_8878, n9025);
  and g15998 (n9026, n_8877, n_8878);
  and g15999 (n9027, n_8564, n_8562);
  not g16000 (n_8879, n9027);
  and g16001 (n9028, n_8563, n_8879);
  and g16002 (n9029, n_8520, n_8564);
  and g16003 (n9030, n_8521, n9029);
  and g16004 (n9031, n_8565, n9030);
  and g16005 (n9032, n_8520, n_8518);
  not g16006 (n_8880, n9032);
  and g16007 (n9033, n_8519, n_8880);
  not g16008 (n_8881, n9031);
  not g16009 (n_8882, n9033);
  and g16010 (n9034, n_8881, n_8882);
  not g16015 (n_8883, n9034);
  not g16016 (n_8884, n9038);
  and g16017 (n9039, n_8883, n_8884);
  not g16018 (n_8885, n9039);
  and g16019 (n9040, n9028, n_8885);
  and g16020 (n9041, n_8881, n9033);
  and g16021 (n9042, n9031, n_8882);
  not g16022 (n_8886, n9041);
  not g16023 (n_8887, n9042);
  and g16024 (n9043, n_8886, n_8887);
  not g16025 (n_8888, n9028);
  not g16026 (n_8889, n9043);
  and g16027 (n9044, n_8888, n_8889);
  and g16028 (n9045, n_8662, n_8663);
  not g16029 (n_8890, n9044);
  not g16030 (n_8891, n9045);
  and g16031 (n9046, n_8890, n_8891);
  not g16032 (n_8892, n9040);
  and g16033 (n9047, n_8892, n9046);
  and g16034 (n9048, n_8892, n_8890);
  not g16035 (n_8893, n9048);
  and g16036 (n9049, n9045, n_8893);
  not g16037 (n_8894, n9047);
  not g16038 (n_8895, n9049);
  and g16039 (n9050, n_8894, n_8895);
  not g16040 (n_8896, n9026);
  not g16041 (n_8897, n9050);
  and g16042 (n9051, n_8896, n_8897);
  and g16043 (n9052, n_8890, n9045);
  and g16044 (n9053, n_8892, n9052);
  and g16045 (n9054, n_8891, n_8893);
  not g16046 (n_8898, n9053);
  not g16047 (n_8899, n9054);
  and g16048 (n9055, n_8898, n_8899);
  not g16049 (n_8900, n9055);
  and g16050 (n9056, n9026, n_8900);
  and g16051 (n9057, n_8854, n_8855);
  not g16052 (n_8901, n9056);
  and g16053 (n9058, n_8901, n9057);
  not g16054 (n_8902, n9051);
  and g16055 (n9059, n_8902, n9058);
  and g16056 (n9060, n_8902, n_8901);
  not g16057 (n_8903, n9057);
  not g16058 (n_8904, n9060);
  and g16059 (n9061, n_8903, n_8904);
  not g16060 (n_8905, n9059);
  not g16061 (n_8906, n9061);
  and g16062 (n9062, n_8905, n_8906);
  and g16063 (n9063, n_8752, n_8750);
  not g16064 (n_8907, n9063);
  and g16065 (n9064, n_8751, n_8907);
  and g16066 (n9065, n_8708, n_8752);
  and g16067 (n9066, n_8709, n9065);
  and g16068 (n9067, n_8753, n9066);
  and g16069 (n9068, n_8708, n_8706);
  not g16070 (n_8908, n9068);
  and g16071 (n9069, n_8707, n_8908);
  not g16072 (n_8909, n9067);
  not g16073 (n_8910, n9069);
  and g16074 (n9070, n_8909, n_8910);
  not g16079 (n_8911, n9070);
  not g16080 (n_8912, n9074);
  and g16081 (n9075, n_8911, n_8912);
  not g16082 (n_8913, n9075);
  and g16083 (n9076, n9064, n_8913);
  and g16084 (n9077, n_8909, n9069);
  and g16085 (n9078, n9067, n_8910);
  not g16086 (n_8914, n9077);
  not g16087 (n_8915, n9078);
  and g16088 (n9079, n_8914, n_8915);
  not g16089 (n_8916, n9064);
  not g16090 (n_8917, n9079);
  and g16091 (n9080, n_8916, n_8917);
  and g16092 (n9081, n_8850, n_8851);
  not g16093 (n_8918, n9080);
  and g16094 (n9082, n_8918, n9081);
  not g16095 (n_8919, n9076);
  and g16096 (n9083, n_8919, n9082);
  and g16097 (n9084, n_8919, n_8918);
  not g16098 (n_8920, n9081);
  not g16099 (n_8921, n9084);
  and g16100 (n9085, n_8920, n_8921);
  not g16101 (n_8922, n9083);
  not g16102 (n_8923, n9085);
  and g16103 (n9086, n_8922, n_8923);
  and g16104 (n9087, n_8844, n_8842);
  not g16105 (n_8924, n9087);
  and g16106 (n9088, n_8843, n_8924);
  and g16107 (n9089, n_8800, n_8844);
  and g16108 (n9090, n_8801, n9089);
  and g16109 (n9091, n_8845, n9090);
  and g16110 (n9092, n_8800, n_8798);
  not g16111 (n_8925, n9092);
  and g16112 (n9093, n_8799, n_8925);
  not g16113 (n_8926, n9091);
  and g16114 (n9094, n_8926, n9093);
  not g16115 (n_8927, n9093);
  and g16116 (n9095, n9091, n_8927);
  not g16117 (n_8928, n9094);
  not g16118 (n_8929, n9095);
  and g16119 (n9096, n_8928, n_8929);
  not g16120 (n_8930, n9088);
  not g16121 (n_8931, n9096);
  and g16122 (n9097, n_8930, n_8931);
  and g16123 (n9098, n_8926, n_8927);
  not g16128 (n_8932, n9098);
  not g16129 (n_8933, n9102);
  and g16130 (n9103, n_8932, n_8933);
  not g16131 (n_8934, n9103);
  and g16132 (n9104, n9088, n_8934);
  not g16133 (n_8935, n9097);
  not g16134 (n_8936, n9104);
  and g16135 (n9105, n_8935, n_8936);
  not g16136 (n_8937, n9086);
  and g16137 (n9106, n_8937, n9105);
  and g16138 (n9107, n_8918, n_8920);
  and g16139 (n9108, n_8919, n9107);
  and g16140 (n9109, n9081, n_8921);
  not g16141 (n_8938, n9108);
  not g16142 (n_8939, n9109);
  and g16143 (n9110, n_8938, n_8939);
  not g16144 (n_8940, n9105);
  not g16145 (n_8941, n9110);
  and g16146 (n9111, n_8940, n_8941);
  not g16147 (n_8942, n9106);
  not g16148 (n_8943, n9111);
  and g16149 (n9112, n_8942, n_8943);
  not g16150 (n_8944, n9062);
  and g16151 (n9113, n_8944, n9112);
  and g16152 (n9114, n_8901, n_8903);
  and g16153 (n9115, n_8902, n9114);
  and g16154 (n9116, n9057, n_8904);
  not g16155 (n_8945, n9115);
  not g16156 (n_8946, n9116);
  and g16157 (n9117, n_8945, n_8946);
  not g16158 (n_8947, n9112);
  not g16159 (n_8948, n9117);
  and g16160 (n9118, n_8947, n_8948);
  not g16161 (n_8949, n9113);
  not g16162 (n_8950, n9118);
  and g16163 (n9119, n_8949, n_8950);
  not g16164 (n_8951, n9007);
  and g16165 (n9120, n_8951, n9119);
  and g16166 (n9121, n_8860, n_8862);
  and g16167 (n9122, n_8861, n9121);
  and g16168 (n9123, n9002, n_8863);
  not g16169 (n_8952, n9122);
  not g16170 (n_8953, n9123);
  and g16171 (n9124, n_8952, n_8953);
  not g16172 (n_8954, n9119);
  not g16173 (n_8955, n9124);
  and g16174 (n9125, n_8954, n_8955);
  not g16175 (n_8956, n9120);
  not g16176 (n_8957, n9125);
  and g16177 (n9126, n_8956, n_8957);
  and g16178 (n9127, \A[394] , \A[395] );
  not g16179 (n_8960, \A[395] );
  and g16180 (n9128, \A[394] , n_8960);
  not g16181 (n_8961, \A[394] );
  and g16182 (n9129, n_8961, \A[395] );
  not g16183 (n_8962, n9128);
  not g16184 (n_8963, n9129);
  and g16185 (n9130, n_8962, n_8963);
  not g16186 (n_8965, n9130);
  and g16187 (n9131, \A[396] , n_8965);
  not g16188 (n_8966, n9127);
  not g16189 (n_8967, n9131);
  and g16190 (n9132, n_8966, n_8967);
  and g16191 (n9133, \A[391] , \A[392] );
  not g16192 (n_8970, \A[392] );
  and g16193 (n9134, \A[391] , n_8970);
  not g16194 (n_8971, \A[391] );
  and g16195 (n9135, n_8971, \A[392] );
  not g16196 (n_8972, n9134);
  not g16197 (n_8973, n9135);
  and g16198 (n9136, n_8972, n_8973);
  not g16199 (n_8975, n9136);
  and g16200 (n9137, \A[393] , n_8975);
  not g16201 (n_8976, n9133);
  not g16202 (n_8977, n9137);
  and g16203 (n9138, n_8976, n_8977);
  not g16204 (n_8978, n9138);
  and g16205 (n9139, n9132, n_8978);
  not g16206 (n_8979, n9132);
  and g16207 (n9140, n_8979, n9138);
  and g16208 (n9141, \A[393] , n_8972);
  and g16209 (n9142, n_8973, n9141);
  not g16210 (n_8980, \A[393] );
  and g16211 (n9143, n_8980, n_8975);
  not g16212 (n_8981, n9142);
  not g16213 (n_8982, n9143);
  and g16214 (n9144, n_8981, n_8982);
  and g16215 (n9145, \A[396] , n_8962);
  and g16216 (n9146, n_8963, n9145);
  not g16217 (n_8983, \A[396] );
  and g16218 (n9147, n_8983, n_8965);
  not g16219 (n_8984, n9146);
  not g16220 (n_8985, n9147);
  and g16221 (n9148, n_8984, n_8985);
  not g16222 (n_8986, n9144);
  not g16223 (n_8987, n9148);
  and g16224 (n9149, n_8986, n_8987);
  not g16225 (n_8988, n9140);
  and g16226 (n9150, n_8988, n9149);
  not g16227 (n_8989, n9139);
  and g16228 (n9151, n_8989, n9150);
  and g16229 (n9152, n_8989, n_8988);
  not g16230 (n_8990, n9149);
  not g16231 (n_8991, n9152);
  and g16232 (n9153, n_8990, n_8991);
  not g16233 (n_8992, n9151);
  not g16234 (n_8993, n9153);
  and g16235 (n9154, n_8992, n_8993);
  and g16236 (n9155, n_8986, n9148);
  and g16237 (n9156, n9144, n_8987);
  not g16238 (n_8994, n9155);
  not g16239 (n_8995, n9156);
  and g16240 (n9157, n_8994, n_8995);
  and g16241 (n9158, n9149, n_8991);
  and g16242 (n9159, n_8979, n_8978);
  not g16243 (n_8996, n9158);
  not g16244 (n_8997, n9159);
  and g16245 (n9160, n_8996, n_8997);
  not g16246 (n_8998, n9157);
  not g16247 (n_8999, n9160);
  and g16248 (n9161, n_8998, n_8999);
  not g16249 (n_9000, n9154);
  not g16250 (n_9001, n9161);
  and g16251 (n9162, n_9000, n_9001);
  and g16252 (n9163, n_9000, n_8999);
  and g16253 (n9164, \A[400] , \A[401] );
  not g16254 (n_9004, \A[401] );
  and g16255 (n9165, \A[400] , n_9004);
  not g16256 (n_9005, \A[400] );
  and g16257 (n9166, n_9005, \A[401] );
  not g16258 (n_9006, n9165);
  not g16259 (n_9007, n9166);
  and g16260 (n9167, n_9006, n_9007);
  not g16261 (n_9009, n9167);
  and g16262 (n9168, \A[402] , n_9009);
  not g16263 (n_9010, n9164);
  not g16264 (n_9011, n9168);
  and g16265 (n9169, n_9010, n_9011);
  and g16266 (n9170, \A[397] , \A[398] );
  not g16267 (n_9014, \A[398] );
  and g16268 (n9171, \A[397] , n_9014);
  not g16269 (n_9015, \A[397] );
  and g16270 (n9172, n_9015, \A[398] );
  not g16271 (n_9016, n9171);
  not g16272 (n_9017, n9172);
  and g16273 (n9173, n_9016, n_9017);
  not g16274 (n_9019, n9173);
  and g16275 (n9174, \A[399] , n_9019);
  not g16276 (n_9020, n9170);
  not g16277 (n_9021, n9174);
  and g16278 (n9175, n_9020, n_9021);
  not g16279 (n_9022, n9169);
  and g16280 (n9176, n_9022, n9175);
  not g16281 (n_9023, n9175);
  and g16282 (n9177, n9169, n_9023);
  not g16283 (n_9024, n9176);
  not g16284 (n_9025, n9177);
  and g16285 (n9178, n_9024, n_9025);
  and g16286 (n9179, \A[399] , n_9016);
  and g16287 (n9180, n_9017, n9179);
  not g16288 (n_9026, \A[399] );
  and g16289 (n9181, n_9026, n_9019);
  not g16290 (n_9027, n9180);
  not g16291 (n_9028, n9181);
  and g16292 (n9182, n_9027, n_9028);
  and g16293 (n9183, \A[402] , n_9006);
  and g16294 (n9184, n_9007, n9183);
  not g16295 (n_9029, \A[402] );
  and g16296 (n9185, n_9029, n_9009);
  not g16297 (n_9030, n9184);
  not g16298 (n_9031, n9185);
  and g16299 (n9186, n_9030, n_9031);
  not g16300 (n_9032, n9182);
  not g16301 (n_9033, n9186);
  and g16302 (n9187, n_9032, n_9033);
  not g16303 (n_9034, n9178);
  and g16304 (n9188, n_9034, n9187);
  and g16305 (n9189, n_9022, n_9023);
  not g16306 (n_9035, n9188);
  not g16307 (n_9036, n9189);
  and g16308 (n9190, n_9035, n_9036);
  and g16309 (n9191, n_9024, n9187);
  and g16310 (n9192, n_9025, n9191);
  not g16311 (n_9037, n9187);
  and g16312 (n9193, n_9034, n_9037);
  not g16313 (n_9038, n9192);
  not g16314 (n_9039, n9193);
  and g16315 (n9194, n_9038, n_9039);
  not g16316 (n_9040, n9190);
  not g16317 (n_9041, n9194);
  and g16318 (n9195, n_9040, n_9041);
  and g16319 (n9196, n_9032, n9186);
  and g16320 (n9197, n9182, n_9033);
  not g16321 (n_9042, n9196);
  not g16322 (n_9043, n9197);
  and g16323 (n9198, n_9042, n_9043);
  not g16324 (n_9044, n9198);
  and g16325 (n9199, n_8998, n_9044);
  not g16326 (n_9045, n9195);
  and g16327 (n9200, n_9045, n9199);
  not g16328 (n_9046, n9163);
  and g16329 (n9201, n_9046, n9200);
  and g16330 (n9202, n_9040, n_9044);
  not g16331 (n_9047, n9202);
  and g16332 (n9203, n_9041, n_9047);
  not g16333 (n_9048, n9201);
  and g16334 (n9204, n_9048, n9203);
  not g16335 (n_9049, n9203);
  and g16336 (n9205, n9201, n_9049);
  not g16337 (n_9050, n9204);
  not g16338 (n_9051, n9205);
  and g16339 (n9206, n_9050, n_9051);
  not g16340 (n_9052, n9162);
  not g16341 (n_9053, n9206);
  and g16342 (n9207, n_9052, n_9053);
  and g16343 (n9208, n_9048, n_9049);
  not g16348 (n_9054, n9208);
  not g16349 (n_9055, n9212);
  and g16350 (n9213, n_9054, n_9055);
  not g16351 (n_9056, n9213);
  and g16352 (n9214, n9162, n_9056);
  not g16353 (n_9057, n9207);
  not g16354 (n_9058, n9214);
  and g16355 (n9215, n_9057, n_9058);
  and g16356 (n9216, \A[406] , \A[407] );
  not g16357 (n_9061, \A[407] );
  and g16358 (n9217, \A[406] , n_9061);
  not g16359 (n_9062, \A[406] );
  and g16360 (n9218, n_9062, \A[407] );
  not g16361 (n_9063, n9217);
  not g16362 (n_9064, n9218);
  and g16363 (n9219, n_9063, n_9064);
  not g16364 (n_9066, n9219);
  and g16365 (n9220, \A[408] , n_9066);
  not g16366 (n_9067, n9216);
  not g16367 (n_9068, n9220);
  and g16368 (n9221, n_9067, n_9068);
  and g16369 (n9222, \A[403] , \A[404] );
  not g16370 (n_9071, \A[404] );
  and g16371 (n9223, \A[403] , n_9071);
  not g16372 (n_9072, \A[403] );
  and g16373 (n9224, n_9072, \A[404] );
  not g16374 (n_9073, n9223);
  not g16375 (n_9074, n9224);
  and g16376 (n9225, n_9073, n_9074);
  not g16377 (n_9076, n9225);
  and g16378 (n9226, \A[405] , n_9076);
  not g16379 (n_9077, n9222);
  not g16380 (n_9078, n9226);
  and g16381 (n9227, n_9077, n_9078);
  not g16382 (n_9079, n9227);
  and g16383 (n9228, n9221, n_9079);
  not g16384 (n_9080, n9221);
  and g16385 (n9229, n_9080, n9227);
  and g16386 (n9230, \A[405] , n_9073);
  and g16387 (n9231, n_9074, n9230);
  not g16388 (n_9081, \A[405] );
  and g16389 (n9232, n_9081, n_9076);
  not g16390 (n_9082, n9231);
  not g16391 (n_9083, n9232);
  and g16392 (n9233, n_9082, n_9083);
  and g16393 (n9234, \A[408] , n_9063);
  and g16394 (n9235, n_9064, n9234);
  not g16395 (n_9084, \A[408] );
  and g16396 (n9236, n_9084, n_9066);
  not g16397 (n_9085, n9235);
  not g16398 (n_9086, n9236);
  and g16399 (n9237, n_9085, n_9086);
  not g16400 (n_9087, n9233);
  not g16401 (n_9088, n9237);
  and g16402 (n9238, n_9087, n_9088);
  not g16403 (n_9089, n9229);
  and g16404 (n9239, n_9089, n9238);
  not g16405 (n_9090, n9228);
  and g16406 (n9240, n_9090, n9239);
  and g16407 (n9241, n_9090, n_9089);
  not g16408 (n_9091, n9238);
  not g16409 (n_9092, n9241);
  and g16410 (n9242, n_9091, n_9092);
  not g16411 (n_9093, n9240);
  not g16412 (n_9094, n9242);
  and g16413 (n9243, n_9093, n_9094);
  and g16414 (n9244, n_9087, n9237);
  and g16415 (n9245, n9233, n_9088);
  not g16416 (n_9095, n9244);
  not g16417 (n_9096, n9245);
  and g16418 (n9246, n_9095, n_9096);
  and g16419 (n9247, n9238, n_9092);
  and g16420 (n9248, n_9080, n_9079);
  not g16421 (n_9097, n9247);
  not g16422 (n_9098, n9248);
  and g16423 (n9249, n_9097, n_9098);
  not g16424 (n_9099, n9246);
  not g16425 (n_9100, n9249);
  and g16426 (n9250, n_9099, n_9100);
  not g16427 (n_9101, n9243);
  not g16428 (n_9102, n9250);
  and g16429 (n9251, n_9101, n_9102);
  and g16430 (n9252, n_9101, n_9100);
  and g16431 (n9253, \A[412] , \A[413] );
  not g16432 (n_9105, \A[413] );
  and g16433 (n9254, \A[412] , n_9105);
  not g16434 (n_9106, \A[412] );
  and g16435 (n9255, n_9106, \A[413] );
  not g16436 (n_9107, n9254);
  not g16437 (n_9108, n9255);
  and g16438 (n9256, n_9107, n_9108);
  not g16439 (n_9110, n9256);
  and g16440 (n9257, \A[414] , n_9110);
  not g16441 (n_9111, n9253);
  not g16442 (n_9112, n9257);
  and g16443 (n9258, n_9111, n_9112);
  and g16444 (n9259, \A[409] , \A[410] );
  not g16445 (n_9115, \A[410] );
  and g16446 (n9260, \A[409] , n_9115);
  not g16447 (n_9116, \A[409] );
  and g16448 (n9261, n_9116, \A[410] );
  not g16449 (n_9117, n9260);
  not g16450 (n_9118, n9261);
  and g16451 (n9262, n_9117, n_9118);
  not g16452 (n_9120, n9262);
  and g16453 (n9263, \A[411] , n_9120);
  not g16454 (n_9121, n9259);
  not g16455 (n_9122, n9263);
  and g16456 (n9264, n_9121, n_9122);
  not g16457 (n_9123, n9258);
  and g16458 (n9265, n_9123, n9264);
  not g16459 (n_9124, n9264);
  and g16460 (n9266, n9258, n_9124);
  not g16461 (n_9125, n9265);
  not g16462 (n_9126, n9266);
  and g16463 (n9267, n_9125, n_9126);
  and g16464 (n9268, \A[411] , n_9117);
  and g16465 (n9269, n_9118, n9268);
  not g16466 (n_9127, \A[411] );
  and g16467 (n9270, n_9127, n_9120);
  not g16468 (n_9128, n9269);
  not g16469 (n_9129, n9270);
  and g16470 (n9271, n_9128, n_9129);
  and g16471 (n9272, \A[414] , n_9107);
  and g16472 (n9273, n_9108, n9272);
  not g16473 (n_9130, \A[414] );
  and g16474 (n9274, n_9130, n_9110);
  not g16475 (n_9131, n9273);
  not g16476 (n_9132, n9274);
  and g16477 (n9275, n_9131, n_9132);
  not g16478 (n_9133, n9271);
  not g16479 (n_9134, n9275);
  and g16480 (n9276, n_9133, n_9134);
  not g16481 (n_9135, n9267);
  and g16482 (n9277, n_9135, n9276);
  and g16483 (n9278, n_9123, n_9124);
  not g16484 (n_9136, n9277);
  not g16485 (n_9137, n9278);
  and g16486 (n9279, n_9136, n_9137);
  and g16487 (n9280, n_9125, n9276);
  and g16488 (n9281, n_9126, n9280);
  not g16489 (n_9138, n9276);
  and g16490 (n9282, n_9135, n_9138);
  not g16491 (n_9139, n9281);
  not g16492 (n_9140, n9282);
  and g16493 (n9283, n_9139, n_9140);
  not g16494 (n_9141, n9279);
  not g16495 (n_9142, n9283);
  and g16496 (n9284, n_9141, n_9142);
  and g16497 (n9285, n_9133, n9275);
  and g16498 (n9286, n9271, n_9134);
  not g16499 (n_9143, n9285);
  not g16500 (n_9144, n9286);
  and g16501 (n9287, n_9143, n_9144);
  not g16502 (n_9145, n9287);
  and g16503 (n9288, n_9099, n_9145);
  not g16504 (n_9146, n9284);
  and g16505 (n9289, n_9146, n9288);
  not g16506 (n_9147, n9252);
  and g16507 (n9290, n_9147, n9289);
  and g16508 (n9291, n_9141, n_9145);
  not g16509 (n_9148, n9291);
  and g16510 (n9292, n_9142, n_9148);
  not g16511 (n_9149, n9290);
  not g16512 (n_9150, n9292);
  and g16513 (n9293, n_9149, n_9150);
  not g16518 (n_9151, n9293);
  not g16519 (n_9152, n9297);
  and g16520 (n9298, n_9151, n_9152);
  not g16521 (n_9153, n9298);
  and g16522 (n9299, n9251, n_9153);
  and g16523 (n9300, n_9149, n9292);
  and g16524 (n9301, n9290, n_9150);
  not g16525 (n_9154, n9300);
  not g16526 (n_9155, n9301);
  and g16527 (n9302, n_9154, n_9155);
  not g16528 (n_9156, n9251);
  not g16529 (n_9157, n9302);
  and g16530 (n9303, n_9156, n_9157);
  and g16531 (n9304, n_9146, n_9145);
  and g16532 (n9305, n_9099, n_9147);
  not g16533 (n_9158, n9304);
  and g16534 (n9306, n_9158, n9305);
  not g16535 (n_9159, n9305);
  and g16536 (n9307, n9304, n_9159);
  not g16537 (n_9160, n9306);
  not g16538 (n_9161, n9307);
  and g16539 (n9308, n_9160, n_9161);
  and g16540 (n9309, n_9045, n_9044);
  and g16541 (n9310, n_8998, n_9046);
  not g16542 (n_9162, n9309);
  and g16543 (n9311, n_9162, n9310);
  not g16544 (n_9163, n9310);
  and g16545 (n9312, n9309, n_9163);
  not g16546 (n_9164, n9311);
  not g16547 (n_9165, n9312);
  and g16548 (n9313, n_9164, n_9165);
  not g16549 (n_9166, n9308);
  not g16550 (n_9167, n9313);
  and g16551 (n9314, n_9166, n_9167);
  not g16552 (n_9168, n9303);
  not g16553 (n_9169, n9314);
  and g16554 (n9315, n_9168, n_9169);
  not g16555 (n_9170, n9299);
  and g16556 (n9316, n_9170, n9315);
  and g16557 (n9317, n_9170, n_9168);
  not g16558 (n_9171, n9317);
  and g16559 (n9318, n9314, n_9171);
  not g16560 (n_9172, n9316);
  not g16561 (n_9173, n9318);
  and g16562 (n9319, n_9172, n_9173);
  not g16563 (n_9174, n9215);
  not g16564 (n_9175, n9319);
  and g16565 (n9320, n_9174, n_9175);
  and g16566 (n9321, n_9168, n9314);
  and g16567 (n9322, n_9170, n9321);
  and g16568 (n9323, n_9169, n_9171);
  not g16569 (n_9176, n9322);
  not g16570 (n_9177, n9323);
  and g16571 (n9324, n_9176, n_9177);
  not g16572 (n_9178, n9324);
  and g16573 (n9325, n9215, n_9178);
  and g16574 (n9326, n_9166, n9313);
  and g16575 (n9327, n9308, n_9167);
  not g16576 (n_9179, n9326);
  not g16577 (n_9180, n9327);
  and g16578 (n9328, n_9179, n_9180);
  not g16579 (n_9182, \A[385] );
  and g16580 (n9329, n_9182, \A[386] );
  not g16581 (n_9184, \A[386] );
  and g16582 (n9330, \A[385] , n_9184);
  not g16583 (n_9186, n9330);
  and g16584 (n9331, \A[387] , n_9186);
  not g16585 (n_9187, n9329);
  and g16586 (n9332, n_9187, n9331);
  and g16587 (n9333, n_9187, n_9186);
  not g16588 (n_9188, \A[387] );
  not g16589 (n_9189, n9333);
  and g16590 (n9334, n_9188, n_9189);
  not g16591 (n_9190, n9332);
  not g16592 (n_9191, n9334);
  and g16593 (n9335, n_9190, n_9191);
  not g16594 (n_9193, \A[388] );
  and g16595 (n9336, n_9193, \A[389] );
  not g16596 (n_9195, \A[389] );
  and g16597 (n9337, \A[388] , n_9195);
  not g16598 (n_9197, n9337);
  and g16599 (n9338, \A[390] , n_9197);
  not g16600 (n_9198, n9336);
  and g16601 (n9339, n_9198, n9338);
  and g16602 (n9340, n_9198, n_9197);
  not g16603 (n_9199, \A[390] );
  not g16604 (n_9200, n9340);
  and g16605 (n9341, n_9199, n_9200);
  not g16606 (n_9201, n9339);
  not g16607 (n_9202, n9341);
  and g16608 (n9342, n_9201, n_9202);
  not g16609 (n_9203, n9335);
  and g16610 (n9343, n_9203, n9342);
  not g16611 (n_9204, n9342);
  and g16612 (n9344, n9335, n_9204);
  not g16613 (n_9205, n9343);
  not g16614 (n_9206, n9344);
  and g16615 (n9345, n_9205, n_9206);
  and g16616 (n9346, \A[388] , \A[389] );
  and g16617 (n9347, \A[390] , n_9200);
  not g16618 (n_9207, n9346);
  not g16619 (n_9208, n9347);
  and g16620 (n9348, n_9207, n_9208);
  and g16621 (n9349, \A[385] , \A[386] );
  and g16622 (n9350, \A[387] , n_9189);
  not g16623 (n_9209, n9349);
  not g16624 (n_9210, n9350);
  and g16625 (n9351, n_9209, n_9210);
  not g16626 (n_9211, n9348);
  and g16627 (n9352, n_9211, n9351);
  not g16628 (n_9212, n9351);
  and g16629 (n9353, n9348, n_9212);
  not g16630 (n_9213, n9352);
  not g16631 (n_9214, n9353);
  and g16632 (n9354, n_9213, n_9214);
  and g16633 (n9355, n_9203, n_9204);
  not g16634 (n_9215, n9354);
  and g16635 (n9356, n_9215, n9355);
  and g16636 (n9357, n_9211, n_9212);
  not g16637 (n_9216, n9356);
  not g16638 (n_9217, n9357);
  and g16639 (n9358, n_9216, n_9217);
  and g16640 (n9359, n_9213, n9355);
  and g16641 (n9360, n_9214, n9359);
  not g16642 (n_9218, n9355);
  and g16643 (n9361, n_9215, n_9218);
  not g16644 (n_9219, n9360);
  not g16645 (n_9220, n9361);
  and g16646 (n9362, n_9219, n_9220);
  not g16647 (n_9221, n9358);
  not g16648 (n_9222, n9362);
  and g16649 (n9363, n_9221, n_9222);
  not g16650 (n_9223, n9345);
  not g16651 (n_9224, n9363);
  and g16652 (n9364, n_9223, n_9224);
  not g16653 (n_9226, \A[379] );
  and g16654 (n9365, n_9226, \A[380] );
  not g16655 (n_9228, \A[380] );
  and g16656 (n9366, \A[379] , n_9228);
  not g16657 (n_9230, n9366);
  and g16658 (n9367, \A[381] , n_9230);
  not g16659 (n_9231, n9365);
  and g16660 (n9368, n_9231, n9367);
  and g16661 (n9369, n_9231, n_9230);
  not g16662 (n_9232, \A[381] );
  not g16663 (n_9233, n9369);
  and g16664 (n9370, n_9232, n_9233);
  not g16665 (n_9234, n9368);
  not g16666 (n_9235, n9370);
  and g16667 (n9371, n_9234, n_9235);
  not g16668 (n_9237, \A[382] );
  and g16669 (n9372, n_9237, \A[383] );
  not g16670 (n_9239, \A[383] );
  and g16671 (n9373, \A[382] , n_9239);
  not g16672 (n_9241, n9373);
  and g16673 (n9374, \A[384] , n_9241);
  not g16674 (n_9242, n9372);
  and g16675 (n9375, n_9242, n9374);
  and g16676 (n9376, n_9242, n_9241);
  not g16677 (n_9243, \A[384] );
  not g16678 (n_9244, n9376);
  and g16679 (n9377, n_9243, n_9244);
  not g16680 (n_9245, n9375);
  not g16681 (n_9246, n9377);
  and g16682 (n9378, n_9245, n_9246);
  not g16683 (n_9247, n9371);
  and g16684 (n9379, n_9247, n9378);
  not g16685 (n_9248, n9378);
  and g16686 (n9380, n9371, n_9248);
  not g16687 (n_9249, n9379);
  not g16688 (n_9250, n9380);
  and g16689 (n9381, n_9249, n_9250);
  and g16690 (n9382, \A[382] , \A[383] );
  and g16691 (n9383, \A[384] , n_9244);
  not g16692 (n_9251, n9382);
  not g16693 (n_9252, n9383);
  and g16694 (n9384, n_9251, n_9252);
  and g16695 (n9385, \A[379] , \A[380] );
  and g16696 (n9386, \A[381] , n_9233);
  not g16697 (n_9253, n9385);
  not g16698 (n_9254, n9386);
  and g16699 (n9387, n_9253, n_9254);
  not g16700 (n_9255, n9384);
  and g16701 (n9388, n_9255, n9387);
  not g16702 (n_9256, n9387);
  and g16703 (n9389, n9384, n_9256);
  not g16704 (n_9257, n9388);
  not g16705 (n_9258, n9389);
  and g16706 (n9390, n_9257, n_9258);
  and g16707 (n9391, n_9247, n_9248);
  not g16708 (n_9259, n9390);
  and g16709 (n9392, n_9259, n9391);
  and g16710 (n9393, n_9255, n_9256);
  not g16711 (n_9260, n9392);
  not g16712 (n_9261, n9393);
  and g16713 (n9394, n_9260, n_9261);
  and g16714 (n9395, n_9257, n9391);
  and g16715 (n9396, n_9258, n9395);
  not g16716 (n_9262, n9391);
  and g16717 (n9397, n_9259, n_9262);
  not g16718 (n_9263, n9396);
  not g16719 (n_9264, n9397);
  and g16720 (n9398, n_9263, n_9264);
  not g16721 (n_9265, n9394);
  not g16722 (n_9266, n9398);
  and g16723 (n9399, n_9265, n_9266);
  not g16724 (n_9267, n9381);
  not g16725 (n_9268, n9399);
  and g16726 (n9400, n_9267, n_9268);
  not g16727 (n_9269, n9364);
  and g16728 (n9401, n_9269, n9400);
  not g16729 (n_9270, n9400);
  and g16730 (n9402, n9364, n_9270);
  not g16731 (n_9271, n9401);
  not g16732 (n_9272, n9402);
  and g16733 (n9403, n_9271, n_9272);
  not g16734 (n_9274, \A[373] );
  and g16735 (n9404, n_9274, \A[374] );
  not g16736 (n_9276, \A[374] );
  and g16737 (n9405, \A[373] , n_9276);
  not g16738 (n_9278, n9405);
  and g16739 (n9406, \A[375] , n_9278);
  not g16740 (n_9279, n9404);
  and g16741 (n9407, n_9279, n9406);
  and g16742 (n9408, n_9279, n_9278);
  not g16743 (n_9280, \A[375] );
  not g16744 (n_9281, n9408);
  and g16745 (n9409, n_9280, n_9281);
  not g16746 (n_9282, n9407);
  not g16747 (n_9283, n9409);
  and g16748 (n9410, n_9282, n_9283);
  not g16749 (n_9285, \A[376] );
  and g16750 (n9411, n_9285, \A[377] );
  not g16751 (n_9287, \A[377] );
  and g16752 (n9412, \A[376] , n_9287);
  not g16753 (n_9289, n9412);
  and g16754 (n9413, \A[378] , n_9289);
  not g16755 (n_9290, n9411);
  and g16756 (n9414, n_9290, n9413);
  and g16757 (n9415, n_9290, n_9289);
  not g16758 (n_9291, \A[378] );
  not g16759 (n_9292, n9415);
  and g16760 (n9416, n_9291, n_9292);
  not g16761 (n_9293, n9414);
  not g16762 (n_9294, n9416);
  and g16763 (n9417, n_9293, n_9294);
  not g16764 (n_9295, n9410);
  and g16765 (n9418, n_9295, n9417);
  not g16766 (n_9296, n9417);
  and g16767 (n9419, n9410, n_9296);
  not g16768 (n_9297, n9418);
  not g16769 (n_9298, n9419);
  and g16770 (n9420, n_9297, n_9298);
  and g16771 (n9421, \A[376] , \A[377] );
  and g16772 (n9422, \A[378] , n_9292);
  not g16773 (n_9299, n9421);
  not g16774 (n_9300, n9422);
  and g16775 (n9423, n_9299, n_9300);
  and g16776 (n9424, \A[373] , \A[374] );
  and g16777 (n9425, \A[375] , n_9281);
  not g16778 (n_9301, n9424);
  not g16779 (n_9302, n9425);
  and g16780 (n9426, n_9301, n_9302);
  not g16781 (n_9303, n9423);
  and g16782 (n9427, n_9303, n9426);
  not g16783 (n_9304, n9426);
  and g16784 (n9428, n9423, n_9304);
  not g16785 (n_9305, n9427);
  not g16786 (n_9306, n9428);
  and g16787 (n9429, n_9305, n_9306);
  and g16788 (n9430, n_9295, n_9296);
  not g16789 (n_9307, n9429);
  and g16790 (n9431, n_9307, n9430);
  and g16791 (n9432, n_9303, n_9304);
  not g16792 (n_9308, n9431);
  not g16793 (n_9309, n9432);
  and g16794 (n9433, n_9308, n_9309);
  and g16795 (n9434, n_9305, n9430);
  and g16796 (n9435, n_9306, n9434);
  not g16797 (n_9310, n9430);
  and g16798 (n9436, n_9307, n_9310);
  not g16799 (n_9311, n9435);
  not g16800 (n_9312, n9436);
  and g16801 (n9437, n_9311, n_9312);
  not g16802 (n_9313, n9433);
  not g16803 (n_9314, n9437);
  and g16804 (n9438, n_9313, n_9314);
  not g16805 (n_9315, n9420);
  not g16806 (n_9316, n9438);
  and g16807 (n9439, n_9315, n_9316);
  not g16808 (n_9318, \A[367] );
  and g16809 (n9440, n_9318, \A[368] );
  not g16810 (n_9320, \A[368] );
  and g16811 (n9441, \A[367] , n_9320);
  not g16812 (n_9322, n9441);
  and g16813 (n9442, \A[369] , n_9322);
  not g16814 (n_9323, n9440);
  and g16815 (n9443, n_9323, n9442);
  and g16816 (n9444, n_9323, n_9322);
  not g16817 (n_9324, \A[369] );
  not g16818 (n_9325, n9444);
  and g16819 (n9445, n_9324, n_9325);
  not g16820 (n_9326, n9443);
  not g16821 (n_9327, n9445);
  and g16822 (n9446, n_9326, n_9327);
  not g16823 (n_9329, \A[370] );
  and g16824 (n9447, n_9329, \A[371] );
  not g16825 (n_9331, \A[371] );
  and g16826 (n9448, \A[370] , n_9331);
  not g16827 (n_9333, n9448);
  and g16828 (n9449, \A[372] , n_9333);
  not g16829 (n_9334, n9447);
  and g16830 (n9450, n_9334, n9449);
  and g16831 (n9451, n_9334, n_9333);
  not g16832 (n_9335, \A[372] );
  not g16833 (n_9336, n9451);
  and g16834 (n9452, n_9335, n_9336);
  not g16835 (n_9337, n9450);
  not g16836 (n_9338, n9452);
  and g16837 (n9453, n_9337, n_9338);
  not g16838 (n_9339, n9446);
  and g16839 (n9454, n_9339, n9453);
  not g16840 (n_9340, n9453);
  and g16841 (n9455, n9446, n_9340);
  not g16842 (n_9341, n9454);
  not g16843 (n_9342, n9455);
  and g16844 (n9456, n_9341, n_9342);
  and g16845 (n9457, \A[370] , \A[371] );
  and g16846 (n9458, \A[372] , n_9336);
  not g16847 (n_9343, n9457);
  not g16848 (n_9344, n9458);
  and g16849 (n9459, n_9343, n_9344);
  and g16850 (n9460, \A[367] , \A[368] );
  and g16851 (n9461, \A[369] , n_9325);
  not g16852 (n_9345, n9460);
  not g16853 (n_9346, n9461);
  and g16854 (n9462, n_9345, n_9346);
  not g16855 (n_9347, n9459);
  and g16856 (n9463, n_9347, n9462);
  not g16857 (n_9348, n9462);
  and g16858 (n9464, n9459, n_9348);
  not g16859 (n_9349, n9463);
  not g16860 (n_9350, n9464);
  and g16861 (n9465, n_9349, n_9350);
  and g16862 (n9466, n_9339, n_9340);
  not g16863 (n_9351, n9465);
  and g16864 (n9467, n_9351, n9466);
  and g16865 (n9468, n_9347, n_9348);
  not g16866 (n_9352, n9467);
  not g16867 (n_9353, n9468);
  and g16868 (n9469, n_9352, n_9353);
  and g16869 (n9470, n_9349, n9466);
  and g16870 (n9471, n_9350, n9470);
  not g16871 (n_9354, n9466);
  and g16872 (n9472, n_9351, n_9354);
  not g16873 (n_9355, n9471);
  not g16874 (n_9356, n9472);
  and g16875 (n9473, n_9355, n_9356);
  not g16876 (n_9357, n9469);
  not g16877 (n_9358, n9473);
  and g16878 (n9474, n_9357, n_9358);
  not g16879 (n_9359, n9456);
  not g16880 (n_9360, n9474);
  and g16881 (n9475, n_9359, n_9360);
  not g16882 (n_9361, n9439);
  and g16883 (n9476, n_9361, n9475);
  not g16884 (n_9362, n9475);
  and g16885 (n9477, n9439, n_9362);
  not g16886 (n_9363, n9476);
  not g16887 (n_9364, n9477);
  and g16888 (n9478, n_9363, n_9364);
  not g16889 (n_9365, n9403);
  and g16890 (n9479, n_9365, n9478);
  not g16891 (n_9366, n9478);
  and g16892 (n9480, n9403, n_9366);
  not g16893 (n_9367, n9479);
  not g16894 (n_9368, n9480);
  and g16895 (n9481, n_9367, n_9368);
  not g16896 (n_9369, n9328);
  not g16897 (n_9370, n9481);
  and g16898 (n9482, n_9369, n_9370);
  not g16899 (n_9371, n9325);
  and g16900 (n9483, n_9371, n9482);
  not g16901 (n_9372, n9320);
  and g16902 (n9484, n_9372, n9483);
  and g16903 (n9485, n_9372, n_9371);
  not g16904 (n_9373, n9482);
  not g16905 (n_9374, n9485);
  and g16906 (n9486, n_9373, n_9374);
  not g16907 (n_9375, n9484);
  not g16908 (n_9376, n9486);
  and g16909 (n9487, n_9375, n_9376);
  and g16910 (n9488, n_9267, n_9265);
  not g16911 (n_9377, n9488);
  and g16912 (n9489, n_9266, n_9377);
  and g16913 (n9490, n_9223, n_9267);
  and g16914 (n9491, n_9224, n9490);
  and g16915 (n9492, n_9268, n9491);
  and g16916 (n9493, n_9223, n_9221);
  not g16917 (n_9378, n9493);
  and g16918 (n9494, n_9222, n_9378);
  not g16919 (n_9379, n9492);
  not g16920 (n_9380, n9494);
  and g16921 (n9495, n_9379, n_9380);
  not g16926 (n_9381, n9495);
  not g16927 (n_9382, n9499);
  and g16928 (n9500, n_9381, n_9382);
  not g16929 (n_9383, n9500);
  and g16930 (n9501, n9489, n_9383);
  and g16931 (n9502, n_9379, n9494);
  and g16932 (n9503, n9492, n_9380);
  not g16933 (n_9384, n9502);
  not g16934 (n_9385, n9503);
  and g16935 (n9504, n_9384, n_9385);
  not g16936 (n_9386, n9489);
  not g16937 (n_9387, n9504);
  and g16938 (n9505, n_9386, n_9387);
  and g16939 (n9506, n_9365, n_9366);
  not g16940 (n_9388, n9505);
  and g16941 (n9507, n_9388, n9506);
  not g16942 (n_9389, n9501);
  and g16943 (n9508, n_9389, n9507);
  and g16944 (n9509, n_9389, n_9388);
  not g16945 (n_9390, n9506);
  not g16946 (n_9391, n9509);
  and g16947 (n9510, n_9390, n_9391);
  not g16948 (n_9392, n9508);
  not g16949 (n_9393, n9510);
  and g16950 (n9511, n_9392, n_9393);
  and g16951 (n9512, n_9359, n_9357);
  not g16952 (n_9394, n9512);
  and g16953 (n9513, n_9358, n_9394);
  and g16954 (n9514, n_9315, n_9359);
  and g16955 (n9515, n_9316, n9514);
  and g16956 (n9516, n_9360, n9515);
  and g16957 (n9517, n_9315, n_9313);
  not g16958 (n_9395, n9517);
  and g16959 (n9518, n_9314, n_9395);
  not g16960 (n_9396, n9516);
  and g16961 (n9519, n_9396, n9518);
  not g16962 (n_9397, n9518);
  and g16963 (n9520, n9516, n_9397);
  not g16964 (n_9398, n9519);
  not g16965 (n_9399, n9520);
  and g16966 (n9521, n_9398, n_9399);
  not g16967 (n_9400, n9513);
  not g16968 (n_9401, n9521);
  and g16969 (n9522, n_9400, n_9401);
  and g16970 (n9523, n_9396, n_9397);
  not g16975 (n_9402, n9523);
  not g16976 (n_9403, n9527);
  and g16977 (n9528, n_9402, n_9403);
  not g16978 (n_9404, n9528);
  and g16979 (n9529, n9513, n_9404);
  not g16980 (n_9405, n9522);
  not g16981 (n_9406, n9529);
  and g16982 (n9530, n_9405, n_9406);
  not g16983 (n_9407, n9511);
  and g16984 (n9531, n_9407, n9530);
  and g16985 (n9532, n_9388, n_9390);
  and g16986 (n9533, n_9389, n9532);
  and g16987 (n9534, n9506, n_9391);
  not g16988 (n_9408, n9533);
  not g16989 (n_9409, n9534);
  and g16990 (n9535, n_9408, n_9409);
  not g16991 (n_9410, n9530);
  not g16992 (n_9411, n9535);
  and g16993 (n9536, n_9410, n_9411);
  not g16994 (n_9412, n9531);
  not g16995 (n_9413, n9536);
  and g16996 (n9537, n_9412, n_9413);
  not g16997 (n_9414, n9487);
  and g16998 (n9538, n_9414, n9537);
  and g16999 (n9539, n_9371, n_9373);
  and g17000 (n9540, n_9372, n9539);
  and g17001 (n9541, n9482, n_9374);
  not g17002 (n_9415, n9540);
  not g17003 (n_9416, n9541);
  and g17004 (n9542, n_9415, n_9416);
  not g17005 (n_9417, n9537);
  not g17006 (n_9418, n9542);
  and g17007 (n9543, n_9417, n_9418);
  not g17008 (n_9419, n9538);
  not g17009 (n_9420, n9543);
  and g17010 (n9544, n_9419, n_9420);
  and g17011 (n9545, \A[430] , \A[431] );
  not g17012 (n_9423, \A[431] );
  and g17013 (n9546, \A[430] , n_9423);
  not g17014 (n_9424, \A[430] );
  and g17015 (n9547, n_9424, \A[431] );
  not g17016 (n_9425, n9546);
  not g17017 (n_9426, n9547);
  and g17018 (n9548, n_9425, n_9426);
  not g17019 (n_9428, n9548);
  and g17020 (n9549, \A[432] , n_9428);
  not g17021 (n_9429, n9545);
  not g17022 (n_9430, n9549);
  and g17023 (n9550, n_9429, n_9430);
  and g17024 (n9551, \A[427] , \A[428] );
  not g17025 (n_9433, \A[428] );
  and g17026 (n9552, \A[427] , n_9433);
  not g17027 (n_9434, \A[427] );
  and g17028 (n9553, n_9434, \A[428] );
  not g17029 (n_9435, n9552);
  not g17030 (n_9436, n9553);
  and g17031 (n9554, n_9435, n_9436);
  not g17032 (n_9438, n9554);
  and g17033 (n9555, \A[429] , n_9438);
  not g17034 (n_9439, n9551);
  not g17035 (n_9440, n9555);
  and g17036 (n9556, n_9439, n_9440);
  not g17037 (n_9441, n9556);
  and g17038 (n9557, n9550, n_9441);
  not g17039 (n_9442, n9550);
  and g17040 (n9558, n_9442, n9556);
  and g17041 (n9559, \A[429] , n_9435);
  and g17042 (n9560, n_9436, n9559);
  not g17043 (n_9443, \A[429] );
  and g17044 (n9561, n_9443, n_9438);
  not g17045 (n_9444, n9560);
  not g17046 (n_9445, n9561);
  and g17047 (n9562, n_9444, n_9445);
  and g17048 (n9563, \A[432] , n_9425);
  and g17049 (n9564, n_9426, n9563);
  not g17050 (n_9446, \A[432] );
  and g17051 (n9565, n_9446, n_9428);
  not g17052 (n_9447, n9564);
  not g17053 (n_9448, n9565);
  and g17054 (n9566, n_9447, n_9448);
  not g17055 (n_9449, n9562);
  not g17056 (n_9450, n9566);
  and g17057 (n9567, n_9449, n_9450);
  not g17058 (n_9451, n9558);
  and g17059 (n9568, n_9451, n9567);
  not g17060 (n_9452, n9557);
  and g17061 (n9569, n_9452, n9568);
  and g17062 (n9570, n_9452, n_9451);
  not g17063 (n_9453, n9567);
  not g17064 (n_9454, n9570);
  and g17065 (n9571, n_9453, n_9454);
  not g17066 (n_9455, n9569);
  not g17067 (n_9456, n9571);
  and g17068 (n9572, n_9455, n_9456);
  and g17069 (n9573, n_9449, n9566);
  and g17070 (n9574, n9562, n_9450);
  not g17071 (n_9457, n9573);
  not g17072 (n_9458, n9574);
  and g17073 (n9575, n_9457, n_9458);
  and g17074 (n9576, n9567, n_9454);
  and g17075 (n9577, n_9442, n_9441);
  not g17076 (n_9459, n9576);
  not g17077 (n_9460, n9577);
  and g17078 (n9578, n_9459, n_9460);
  not g17079 (n_9461, n9575);
  not g17080 (n_9462, n9578);
  and g17081 (n9579, n_9461, n_9462);
  not g17082 (n_9463, n9572);
  not g17083 (n_9464, n9579);
  and g17084 (n9580, n_9463, n_9464);
  and g17085 (n9581, n_9463, n_9462);
  and g17086 (n9582, \A[436] , \A[437] );
  not g17087 (n_9467, \A[437] );
  and g17088 (n9583, \A[436] , n_9467);
  not g17089 (n_9468, \A[436] );
  and g17090 (n9584, n_9468, \A[437] );
  not g17091 (n_9469, n9583);
  not g17092 (n_9470, n9584);
  and g17093 (n9585, n_9469, n_9470);
  not g17094 (n_9472, n9585);
  and g17095 (n9586, \A[438] , n_9472);
  not g17096 (n_9473, n9582);
  not g17097 (n_9474, n9586);
  and g17098 (n9587, n_9473, n_9474);
  and g17099 (n9588, \A[433] , \A[434] );
  not g17100 (n_9477, \A[434] );
  and g17101 (n9589, \A[433] , n_9477);
  not g17102 (n_9478, \A[433] );
  and g17103 (n9590, n_9478, \A[434] );
  not g17104 (n_9479, n9589);
  not g17105 (n_9480, n9590);
  and g17106 (n9591, n_9479, n_9480);
  not g17107 (n_9482, n9591);
  and g17108 (n9592, \A[435] , n_9482);
  not g17109 (n_9483, n9588);
  not g17110 (n_9484, n9592);
  and g17111 (n9593, n_9483, n_9484);
  not g17112 (n_9485, n9587);
  and g17113 (n9594, n_9485, n9593);
  not g17114 (n_9486, n9593);
  and g17115 (n9595, n9587, n_9486);
  not g17116 (n_9487, n9594);
  not g17117 (n_9488, n9595);
  and g17118 (n9596, n_9487, n_9488);
  and g17119 (n9597, \A[435] , n_9479);
  and g17120 (n9598, n_9480, n9597);
  not g17121 (n_9489, \A[435] );
  and g17122 (n9599, n_9489, n_9482);
  not g17123 (n_9490, n9598);
  not g17124 (n_9491, n9599);
  and g17125 (n9600, n_9490, n_9491);
  and g17126 (n9601, \A[438] , n_9469);
  and g17127 (n9602, n_9470, n9601);
  not g17128 (n_9492, \A[438] );
  and g17129 (n9603, n_9492, n_9472);
  not g17130 (n_9493, n9602);
  not g17131 (n_9494, n9603);
  and g17132 (n9604, n_9493, n_9494);
  not g17133 (n_9495, n9600);
  not g17134 (n_9496, n9604);
  and g17135 (n9605, n_9495, n_9496);
  not g17136 (n_9497, n9596);
  and g17137 (n9606, n_9497, n9605);
  and g17138 (n9607, n_9485, n_9486);
  not g17139 (n_9498, n9606);
  not g17140 (n_9499, n9607);
  and g17141 (n9608, n_9498, n_9499);
  and g17142 (n9609, n_9487, n9605);
  and g17143 (n9610, n_9488, n9609);
  not g17144 (n_9500, n9605);
  and g17145 (n9611, n_9497, n_9500);
  not g17146 (n_9501, n9610);
  not g17147 (n_9502, n9611);
  and g17148 (n9612, n_9501, n_9502);
  not g17149 (n_9503, n9608);
  not g17150 (n_9504, n9612);
  and g17151 (n9613, n_9503, n_9504);
  and g17152 (n9614, n_9495, n9604);
  and g17153 (n9615, n9600, n_9496);
  not g17154 (n_9505, n9614);
  not g17155 (n_9506, n9615);
  and g17156 (n9616, n_9505, n_9506);
  not g17157 (n_9507, n9616);
  and g17158 (n9617, n_9461, n_9507);
  not g17159 (n_9508, n9613);
  and g17160 (n9618, n_9508, n9617);
  not g17161 (n_9509, n9581);
  and g17162 (n9619, n_9509, n9618);
  and g17163 (n9620, n_9503, n_9507);
  not g17164 (n_9510, n9620);
  and g17165 (n9621, n_9504, n_9510);
  not g17166 (n_9511, n9619);
  not g17167 (n_9512, n9621);
  and g17168 (n9622, n_9511, n_9512);
  not g17173 (n_9513, n9622);
  not g17174 (n_9514, n9626);
  and g17175 (n9627, n_9513, n_9514);
  not g17176 (n_9515, n9627);
  and g17177 (n9628, n9580, n_9515);
  and g17178 (n9629, n_9511, n9621);
  and g17179 (n9630, n9619, n_9512);
  not g17180 (n_9516, n9629);
  not g17181 (n_9517, n9630);
  and g17182 (n9631, n_9516, n_9517);
  not g17183 (n_9518, n9580);
  not g17184 (n_9519, n9631);
  and g17185 (n9632, n_9518, n_9519);
  and g17186 (n9633, n_9508, n_9507);
  and g17187 (n9634, n_9461, n_9509);
  not g17188 (n_9520, n9633);
  and g17189 (n9635, n_9520, n9634);
  not g17190 (n_9521, n9634);
  and g17191 (n9636, n9633, n_9521);
  not g17192 (n_9522, n9635);
  not g17193 (n_9523, n9636);
  and g17194 (n9637, n_9522, n_9523);
  not g17195 (n_9525, \A[421] );
  and g17196 (n9638, n_9525, \A[422] );
  not g17197 (n_9527, \A[422] );
  and g17198 (n9639, \A[421] , n_9527);
  not g17199 (n_9529, n9639);
  and g17200 (n9640, \A[423] , n_9529);
  not g17201 (n_9530, n9638);
  and g17202 (n9641, n_9530, n9640);
  and g17203 (n9642, n_9530, n_9529);
  not g17204 (n_9531, \A[423] );
  not g17205 (n_9532, n9642);
  and g17206 (n9643, n_9531, n_9532);
  not g17207 (n_9533, n9641);
  not g17208 (n_9534, n9643);
  and g17209 (n9644, n_9533, n_9534);
  not g17210 (n_9536, \A[424] );
  and g17211 (n9645, n_9536, \A[425] );
  not g17212 (n_9538, \A[425] );
  and g17213 (n9646, \A[424] , n_9538);
  not g17214 (n_9540, n9646);
  and g17215 (n9647, \A[426] , n_9540);
  not g17216 (n_9541, n9645);
  and g17217 (n9648, n_9541, n9647);
  and g17218 (n9649, n_9541, n_9540);
  not g17219 (n_9542, \A[426] );
  not g17220 (n_9543, n9649);
  and g17221 (n9650, n_9542, n_9543);
  not g17222 (n_9544, n9648);
  not g17223 (n_9545, n9650);
  and g17224 (n9651, n_9544, n_9545);
  not g17225 (n_9546, n9644);
  and g17226 (n9652, n_9546, n9651);
  not g17227 (n_9547, n9651);
  and g17228 (n9653, n9644, n_9547);
  not g17229 (n_9548, n9652);
  not g17230 (n_9549, n9653);
  and g17231 (n9654, n_9548, n_9549);
  and g17232 (n9655, \A[424] , \A[425] );
  and g17233 (n9656, \A[426] , n_9543);
  not g17234 (n_9550, n9655);
  not g17235 (n_9551, n9656);
  and g17236 (n9657, n_9550, n_9551);
  and g17237 (n9658, \A[421] , \A[422] );
  and g17238 (n9659, \A[423] , n_9532);
  not g17239 (n_9552, n9658);
  not g17240 (n_9553, n9659);
  and g17241 (n9660, n_9552, n_9553);
  not g17242 (n_9554, n9657);
  and g17243 (n9661, n_9554, n9660);
  not g17244 (n_9555, n9660);
  and g17245 (n9662, n9657, n_9555);
  not g17246 (n_9556, n9661);
  not g17247 (n_9557, n9662);
  and g17248 (n9663, n_9556, n_9557);
  and g17249 (n9664, n_9546, n_9547);
  not g17250 (n_9558, n9663);
  and g17251 (n9665, n_9558, n9664);
  and g17252 (n9666, n_9554, n_9555);
  not g17253 (n_9559, n9665);
  not g17254 (n_9560, n9666);
  and g17255 (n9667, n_9559, n_9560);
  and g17256 (n9668, n_9556, n9664);
  and g17257 (n9669, n_9557, n9668);
  not g17258 (n_9561, n9664);
  and g17259 (n9670, n_9558, n_9561);
  not g17260 (n_9562, n9669);
  not g17261 (n_9563, n9670);
  and g17262 (n9671, n_9562, n_9563);
  not g17263 (n_9564, n9667);
  not g17264 (n_9565, n9671);
  and g17265 (n9672, n_9564, n_9565);
  not g17266 (n_9566, n9654);
  not g17267 (n_9567, n9672);
  and g17268 (n9673, n_9566, n_9567);
  not g17269 (n_9569, \A[415] );
  and g17270 (n9674, n_9569, \A[416] );
  not g17271 (n_9571, \A[416] );
  and g17272 (n9675, \A[415] , n_9571);
  not g17273 (n_9573, n9675);
  and g17274 (n9676, \A[417] , n_9573);
  not g17275 (n_9574, n9674);
  and g17276 (n9677, n_9574, n9676);
  and g17277 (n9678, n_9574, n_9573);
  not g17278 (n_9575, \A[417] );
  not g17279 (n_9576, n9678);
  and g17280 (n9679, n_9575, n_9576);
  not g17281 (n_9577, n9677);
  not g17282 (n_9578, n9679);
  and g17283 (n9680, n_9577, n_9578);
  not g17284 (n_9580, \A[418] );
  and g17285 (n9681, n_9580, \A[419] );
  not g17286 (n_9582, \A[419] );
  and g17287 (n9682, \A[418] , n_9582);
  not g17288 (n_9584, n9682);
  and g17289 (n9683, \A[420] , n_9584);
  not g17290 (n_9585, n9681);
  and g17291 (n9684, n_9585, n9683);
  and g17292 (n9685, n_9585, n_9584);
  not g17293 (n_9586, \A[420] );
  not g17294 (n_9587, n9685);
  and g17295 (n9686, n_9586, n_9587);
  not g17296 (n_9588, n9684);
  not g17297 (n_9589, n9686);
  and g17298 (n9687, n_9588, n_9589);
  not g17299 (n_9590, n9680);
  and g17300 (n9688, n_9590, n9687);
  not g17301 (n_9591, n9687);
  and g17302 (n9689, n9680, n_9591);
  not g17303 (n_9592, n9688);
  not g17304 (n_9593, n9689);
  and g17305 (n9690, n_9592, n_9593);
  and g17306 (n9691, \A[418] , \A[419] );
  and g17307 (n9692, \A[420] , n_9587);
  not g17308 (n_9594, n9691);
  not g17309 (n_9595, n9692);
  and g17310 (n9693, n_9594, n_9595);
  and g17311 (n9694, \A[415] , \A[416] );
  and g17312 (n9695, \A[417] , n_9576);
  not g17313 (n_9596, n9694);
  not g17314 (n_9597, n9695);
  and g17315 (n9696, n_9596, n_9597);
  not g17316 (n_9598, n9693);
  and g17317 (n9697, n_9598, n9696);
  not g17318 (n_9599, n9696);
  and g17319 (n9698, n9693, n_9599);
  not g17320 (n_9600, n9697);
  not g17321 (n_9601, n9698);
  and g17322 (n9699, n_9600, n_9601);
  and g17323 (n9700, n_9590, n_9591);
  not g17324 (n_9602, n9699);
  and g17325 (n9701, n_9602, n9700);
  and g17326 (n9702, n_9598, n_9599);
  not g17327 (n_9603, n9701);
  not g17328 (n_9604, n9702);
  and g17329 (n9703, n_9603, n_9604);
  and g17330 (n9704, n_9600, n9700);
  and g17331 (n9705, n_9601, n9704);
  not g17332 (n_9605, n9700);
  and g17333 (n9706, n_9602, n_9605);
  not g17334 (n_9606, n9705);
  not g17335 (n_9607, n9706);
  and g17336 (n9707, n_9606, n_9607);
  not g17337 (n_9608, n9703);
  not g17338 (n_9609, n9707);
  and g17339 (n9708, n_9608, n_9609);
  not g17340 (n_9610, n9690);
  not g17341 (n_9611, n9708);
  and g17342 (n9709, n_9610, n_9611);
  not g17343 (n_9612, n9673);
  and g17344 (n9710, n_9612, n9709);
  not g17345 (n_9613, n9709);
  and g17346 (n9711, n9673, n_9613);
  not g17347 (n_9614, n9710);
  not g17348 (n_9615, n9711);
  and g17349 (n9712, n_9614, n_9615);
  not g17350 (n_9616, n9637);
  not g17351 (n_9617, n9712);
  and g17352 (n9713, n_9616, n_9617);
  not g17353 (n_9618, n9632);
  and g17354 (n9714, n_9618, n9713);
  not g17355 (n_9619, n9628);
  and g17356 (n9715, n_9619, n9714);
  and g17357 (n9716, n_9619, n_9618);
  not g17358 (n_9620, n9713);
  not g17359 (n_9621, n9716);
  and g17360 (n9717, n_9620, n_9621);
  not g17361 (n_9622, n9715);
  not g17362 (n_9623, n9717);
  and g17363 (n9718, n_9622, n_9623);
  and g17364 (n9719, n_9610, n_9608);
  not g17365 (n_9624, n9719);
  and g17366 (n9720, n_9609, n_9624);
  and g17367 (n9721, n_9566, n_9610);
  and g17368 (n9722, n_9567, n9721);
  and g17369 (n9723, n_9611, n9722);
  and g17370 (n9724, n_9566, n_9564);
  not g17371 (n_9625, n9724);
  and g17372 (n9725, n_9565, n_9625);
  not g17373 (n_9626, n9723);
  and g17374 (n9726, n_9626, n9725);
  not g17375 (n_9627, n9725);
  and g17376 (n9727, n9723, n_9627);
  not g17377 (n_9628, n9726);
  not g17378 (n_9629, n9727);
  and g17379 (n9728, n_9628, n_9629);
  not g17380 (n_9630, n9720);
  not g17381 (n_9631, n9728);
  and g17382 (n9729, n_9630, n_9631);
  and g17383 (n9730, n_9626, n_9627);
  not g17388 (n_9632, n9730);
  not g17389 (n_9633, n9734);
  and g17390 (n9735, n_9632, n_9633);
  not g17391 (n_9634, n9735);
  and g17392 (n9736, n9720, n_9634);
  not g17393 (n_9635, n9729);
  not g17394 (n_9636, n9736);
  and g17395 (n9737, n_9635, n_9636);
  not g17396 (n_9637, n9718);
  and g17397 (n9738, n_9637, n9737);
  and g17398 (n9739, n_9618, n_9620);
  and g17399 (n9740, n_9619, n9739);
  and g17400 (n9741, n9713, n_9621);
  not g17401 (n_9638, n9740);
  not g17402 (n_9639, n9741);
  and g17403 (n9742, n_9638, n_9639);
  not g17404 (n_9640, n9737);
  not g17405 (n_9641, n9742);
  and g17406 (n9743, n_9640, n_9641);
  not g17407 (n_9642, n9738);
  not g17408 (n_9643, n9743);
  and g17409 (n9744, n_9642, n_9643);
  and g17410 (n9745, \A[442] , \A[443] );
  not g17411 (n_9646, \A[443] );
  and g17412 (n9746, \A[442] , n_9646);
  not g17413 (n_9647, \A[442] );
  and g17414 (n9747, n_9647, \A[443] );
  not g17415 (n_9648, n9746);
  not g17416 (n_9649, n9747);
  and g17417 (n9748, n_9648, n_9649);
  not g17418 (n_9651, n9748);
  and g17419 (n9749, \A[444] , n_9651);
  not g17420 (n_9652, n9745);
  not g17421 (n_9653, n9749);
  and g17422 (n9750, n_9652, n_9653);
  and g17423 (n9751, \A[439] , \A[440] );
  not g17424 (n_9656, \A[440] );
  and g17425 (n9752, \A[439] , n_9656);
  not g17426 (n_9657, \A[439] );
  and g17427 (n9753, n_9657, \A[440] );
  not g17428 (n_9658, n9752);
  not g17429 (n_9659, n9753);
  and g17430 (n9754, n_9658, n_9659);
  not g17431 (n_9661, n9754);
  and g17432 (n9755, \A[441] , n_9661);
  not g17433 (n_9662, n9751);
  not g17434 (n_9663, n9755);
  and g17435 (n9756, n_9662, n_9663);
  not g17436 (n_9664, n9756);
  and g17437 (n9757, n9750, n_9664);
  not g17438 (n_9665, n9750);
  and g17439 (n9758, n_9665, n9756);
  and g17440 (n9759, \A[441] , n_9658);
  and g17441 (n9760, n_9659, n9759);
  not g17442 (n_9666, \A[441] );
  and g17443 (n9761, n_9666, n_9661);
  not g17444 (n_9667, n9760);
  not g17445 (n_9668, n9761);
  and g17446 (n9762, n_9667, n_9668);
  and g17447 (n9763, \A[444] , n_9648);
  and g17448 (n9764, n_9649, n9763);
  not g17449 (n_9669, \A[444] );
  and g17450 (n9765, n_9669, n_9651);
  not g17451 (n_9670, n9764);
  not g17452 (n_9671, n9765);
  and g17453 (n9766, n_9670, n_9671);
  not g17454 (n_9672, n9762);
  not g17455 (n_9673, n9766);
  and g17456 (n9767, n_9672, n_9673);
  not g17457 (n_9674, n9758);
  and g17458 (n9768, n_9674, n9767);
  not g17459 (n_9675, n9757);
  and g17460 (n9769, n_9675, n9768);
  and g17461 (n9770, n_9675, n_9674);
  not g17462 (n_9676, n9767);
  not g17463 (n_9677, n9770);
  and g17464 (n9771, n_9676, n_9677);
  not g17465 (n_9678, n9769);
  not g17466 (n_9679, n9771);
  and g17467 (n9772, n_9678, n_9679);
  and g17468 (n9773, n_9672, n9766);
  and g17469 (n9774, n9762, n_9673);
  not g17470 (n_9680, n9773);
  not g17471 (n_9681, n9774);
  and g17472 (n9775, n_9680, n_9681);
  and g17473 (n9776, n9767, n_9677);
  and g17474 (n9777, n_9665, n_9664);
  not g17475 (n_9682, n9776);
  not g17476 (n_9683, n9777);
  and g17477 (n9778, n_9682, n_9683);
  not g17478 (n_9684, n9775);
  not g17479 (n_9685, n9778);
  and g17480 (n9779, n_9684, n_9685);
  not g17481 (n_9686, n9772);
  not g17482 (n_9687, n9779);
  and g17483 (n9780, n_9686, n_9687);
  and g17484 (n9781, n_9686, n_9685);
  and g17485 (n9782, \A[448] , \A[449] );
  not g17486 (n_9690, \A[449] );
  and g17487 (n9783, \A[448] , n_9690);
  not g17488 (n_9691, \A[448] );
  and g17489 (n9784, n_9691, \A[449] );
  not g17490 (n_9692, n9783);
  not g17491 (n_9693, n9784);
  and g17492 (n9785, n_9692, n_9693);
  not g17493 (n_9695, n9785);
  and g17494 (n9786, \A[450] , n_9695);
  not g17495 (n_9696, n9782);
  not g17496 (n_9697, n9786);
  and g17497 (n9787, n_9696, n_9697);
  and g17498 (n9788, \A[445] , \A[446] );
  not g17499 (n_9700, \A[446] );
  and g17500 (n9789, \A[445] , n_9700);
  not g17501 (n_9701, \A[445] );
  and g17502 (n9790, n_9701, \A[446] );
  not g17503 (n_9702, n9789);
  not g17504 (n_9703, n9790);
  and g17505 (n9791, n_9702, n_9703);
  not g17506 (n_9705, n9791);
  and g17507 (n9792, \A[447] , n_9705);
  not g17508 (n_9706, n9788);
  not g17509 (n_9707, n9792);
  and g17510 (n9793, n_9706, n_9707);
  not g17511 (n_9708, n9787);
  and g17512 (n9794, n_9708, n9793);
  not g17513 (n_9709, n9793);
  and g17514 (n9795, n9787, n_9709);
  not g17515 (n_9710, n9794);
  not g17516 (n_9711, n9795);
  and g17517 (n9796, n_9710, n_9711);
  and g17518 (n9797, \A[447] , n_9702);
  and g17519 (n9798, n_9703, n9797);
  not g17520 (n_9712, \A[447] );
  and g17521 (n9799, n_9712, n_9705);
  not g17522 (n_9713, n9798);
  not g17523 (n_9714, n9799);
  and g17524 (n9800, n_9713, n_9714);
  and g17525 (n9801, \A[450] , n_9692);
  and g17526 (n9802, n_9693, n9801);
  not g17527 (n_9715, \A[450] );
  and g17528 (n9803, n_9715, n_9695);
  not g17529 (n_9716, n9802);
  not g17530 (n_9717, n9803);
  and g17531 (n9804, n_9716, n_9717);
  not g17532 (n_9718, n9800);
  not g17533 (n_9719, n9804);
  and g17534 (n9805, n_9718, n_9719);
  not g17535 (n_9720, n9796);
  and g17536 (n9806, n_9720, n9805);
  and g17537 (n9807, n_9708, n_9709);
  not g17538 (n_9721, n9806);
  not g17539 (n_9722, n9807);
  and g17540 (n9808, n_9721, n_9722);
  and g17541 (n9809, n_9710, n9805);
  and g17542 (n9810, n_9711, n9809);
  not g17543 (n_9723, n9805);
  and g17544 (n9811, n_9720, n_9723);
  not g17545 (n_9724, n9810);
  not g17546 (n_9725, n9811);
  and g17547 (n9812, n_9724, n_9725);
  not g17548 (n_9726, n9808);
  not g17549 (n_9727, n9812);
  and g17550 (n9813, n_9726, n_9727);
  and g17551 (n9814, n_9718, n9804);
  and g17552 (n9815, n9800, n_9719);
  not g17553 (n_9728, n9814);
  not g17554 (n_9729, n9815);
  and g17555 (n9816, n_9728, n_9729);
  not g17556 (n_9730, n9816);
  and g17557 (n9817, n_9684, n_9730);
  not g17558 (n_9731, n9813);
  and g17559 (n9818, n_9731, n9817);
  not g17560 (n_9732, n9781);
  and g17561 (n9819, n_9732, n9818);
  and g17562 (n9820, n_9726, n_9730);
  not g17563 (n_9733, n9820);
  and g17564 (n9821, n_9727, n_9733);
  not g17565 (n_9734, n9819);
  and g17566 (n9822, n_9734, n9821);
  not g17567 (n_9735, n9821);
  and g17568 (n9823, n9819, n_9735);
  not g17569 (n_9736, n9822);
  not g17570 (n_9737, n9823);
  and g17571 (n9824, n_9736, n_9737);
  not g17572 (n_9738, n9780);
  not g17573 (n_9739, n9824);
  and g17574 (n9825, n_9738, n_9739);
  and g17575 (n9826, n_9734, n_9735);
  not g17580 (n_9740, n9826);
  not g17581 (n_9741, n9830);
  and g17582 (n9831, n_9740, n_9741);
  not g17583 (n_9742, n9831);
  and g17584 (n9832, n9780, n_9742);
  not g17585 (n_9743, n9825);
  not g17586 (n_9744, n9832);
  and g17587 (n9833, n_9743, n_9744);
  and g17588 (n9834, \A[454] , \A[455] );
  not g17589 (n_9747, \A[455] );
  and g17590 (n9835, \A[454] , n_9747);
  not g17591 (n_9748, \A[454] );
  and g17592 (n9836, n_9748, \A[455] );
  not g17593 (n_9749, n9835);
  not g17594 (n_9750, n9836);
  and g17595 (n9837, n_9749, n_9750);
  not g17596 (n_9752, n9837);
  and g17597 (n9838, \A[456] , n_9752);
  not g17598 (n_9753, n9834);
  not g17599 (n_9754, n9838);
  and g17600 (n9839, n_9753, n_9754);
  and g17601 (n9840, \A[451] , \A[452] );
  not g17602 (n_9757, \A[452] );
  and g17603 (n9841, \A[451] , n_9757);
  not g17604 (n_9758, \A[451] );
  and g17605 (n9842, n_9758, \A[452] );
  not g17606 (n_9759, n9841);
  not g17607 (n_9760, n9842);
  and g17608 (n9843, n_9759, n_9760);
  not g17609 (n_9762, n9843);
  and g17610 (n9844, \A[453] , n_9762);
  not g17611 (n_9763, n9840);
  not g17612 (n_9764, n9844);
  and g17613 (n9845, n_9763, n_9764);
  not g17614 (n_9765, n9845);
  and g17615 (n9846, n9839, n_9765);
  not g17616 (n_9766, n9839);
  and g17617 (n9847, n_9766, n9845);
  and g17618 (n9848, \A[453] , n_9759);
  and g17619 (n9849, n_9760, n9848);
  not g17620 (n_9767, \A[453] );
  and g17621 (n9850, n_9767, n_9762);
  not g17622 (n_9768, n9849);
  not g17623 (n_9769, n9850);
  and g17624 (n9851, n_9768, n_9769);
  and g17625 (n9852, \A[456] , n_9749);
  and g17626 (n9853, n_9750, n9852);
  not g17627 (n_9770, \A[456] );
  and g17628 (n9854, n_9770, n_9752);
  not g17629 (n_9771, n9853);
  not g17630 (n_9772, n9854);
  and g17631 (n9855, n_9771, n_9772);
  not g17632 (n_9773, n9851);
  not g17633 (n_9774, n9855);
  and g17634 (n9856, n_9773, n_9774);
  not g17635 (n_9775, n9847);
  and g17636 (n9857, n_9775, n9856);
  not g17637 (n_9776, n9846);
  and g17638 (n9858, n_9776, n9857);
  and g17639 (n9859, n_9776, n_9775);
  not g17640 (n_9777, n9856);
  not g17641 (n_9778, n9859);
  and g17642 (n9860, n_9777, n_9778);
  not g17643 (n_9779, n9858);
  not g17644 (n_9780, n9860);
  and g17645 (n9861, n_9779, n_9780);
  and g17646 (n9862, n_9773, n9855);
  and g17647 (n9863, n9851, n_9774);
  not g17648 (n_9781, n9862);
  not g17649 (n_9782, n9863);
  and g17650 (n9864, n_9781, n_9782);
  and g17651 (n9865, n9856, n_9778);
  and g17652 (n9866, n_9766, n_9765);
  not g17653 (n_9783, n9865);
  not g17654 (n_9784, n9866);
  and g17655 (n9867, n_9783, n_9784);
  not g17656 (n_9785, n9864);
  not g17657 (n_9786, n9867);
  and g17658 (n9868, n_9785, n_9786);
  not g17659 (n_9787, n9861);
  not g17660 (n_9788, n9868);
  and g17661 (n9869, n_9787, n_9788);
  and g17662 (n9870, n_9787, n_9786);
  and g17663 (n9871, \A[460] , \A[461] );
  not g17664 (n_9791, \A[461] );
  and g17665 (n9872, \A[460] , n_9791);
  not g17666 (n_9792, \A[460] );
  and g17667 (n9873, n_9792, \A[461] );
  not g17668 (n_9793, n9872);
  not g17669 (n_9794, n9873);
  and g17670 (n9874, n_9793, n_9794);
  not g17671 (n_9796, n9874);
  and g17672 (n9875, \A[462] , n_9796);
  not g17673 (n_9797, n9871);
  not g17674 (n_9798, n9875);
  and g17675 (n9876, n_9797, n_9798);
  and g17676 (n9877, \A[457] , \A[458] );
  not g17677 (n_9801, \A[458] );
  and g17678 (n9878, \A[457] , n_9801);
  not g17679 (n_9802, \A[457] );
  and g17680 (n9879, n_9802, \A[458] );
  not g17681 (n_9803, n9878);
  not g17682 (n_9804, n9879);
  and g17683 (n9880, n_9803, n_9804);
  not g17684 (n_9806, n9880);
  and g17685 (n9881, \A[459] , n_9806);
  not g17686 (n_9807, n9877);
  not g17687 (n_9808, n9881);
  and g17688 (n9882, n_9807, n_9808);
  not g17689 (n_9809, n9876);
  and g17690 (n9883, n_9809, n9882);
  not g17691 (n_9810, n9882);
  and g17692 (n9884, n9876, n_9810);
  not g17693 (n_9811, n9883);
  not g17694 (n_9812, n9884);
  and g17695 (n9885, n_9811, n_9812);
  and g17696 (n9886, \A[459] , n_9803);
  and g17697 (n9887, n_9804, n9886);
  not g17698 (n_9813, \A[459] );
  and g17699 (n9888, n_9813, n_9806);
  not g17700 (n_9814, n9887);
  not g17701 (n_9815, n9888);
  and g17702 (n9889, n_9814, n_9815);
  and g17703 (n9890, \A[462] , n_9793);
  and g17704 (n9891, n_9794, n9890);
  not g17705 (n_9816, \A[462] );
  and g17706 (n9892, n_9816, n_9796);
  not g17707 (n_9817, n9891);
  not g17708 (n_9818, n9892);
  and g17709 (n9893, n_9817, n_9818);
  not g17710 (n_9819, n9889);
  not g17711 (n_9820, n9893);
  and g17712 (n9894, n_9819, n_9820);
  not g17713 (n_9821, n9885);
  and g17714 (n9895, n_9821, n9894);
  and g17715 (n9896, n_9809, n_9810);
  not g17716 (n_9822, n9895);
  not g17717 (n_9823, n9896);
  and g17718 (n9897, n_9822, n_9823);
  and g17719 (n9898, n_9811, n9894);
  and g17720 (n9899, n_9812, n9898);
  not g17721 (n_9824, n9894);
  and g17722 (n9900, n_9821, n_9824);
  not g17723 (n_9825, n9899);
  not g17724 (n_9826, n9900);
  and g17725 (n9901, n_9825, n_9826);
  not g17726 (n_9827, n9897);
  not g17727 (n_9828, n9901);
  and g17728 (n9902, n_9827, n_9828);
  and g17729 (n9903, n_9819, n9893);
  and g17730 (n9904, n9889, n_9820);
  not g17731 (n_9829, n9903);
  not g17732 (n_9830, n9904);
  and g17733 (n9905, n_9829, n_9830);
  not g17734 (n_9831, n9905);
  and g17735 (n9906, n_9785, n_9831);
  not g17736 (n_9832, n9902);
  and g17737 (n9907, n_9832, n9906);
  not g17738 (n_9833, n9870);
  and g17739 (n9908, n_9833, n9907);
  and g17740 (n9909, n_9827, n_9831);
  not g17741 (n_9834, n9909);
  and g17742 (n9910, n_9828, n_9834);
  not g17743 (n_9835, n9908);
  not g17744 (n_9836, n9910);
  and g17745 (n9911, n_9835, n_9836);
  not g17750 (n_9837, n9911);
  not g17751 (n_9838, n9915);
  and g17752 (n9916, n_9837, n_9838);
  not g17753 (n_9839, n9916);
  and g17754 (n9917, n9869, n_9839);
  and g17755 (n9918, n_9835, n9910);
  and g17756 (n9919, n9908, n_9836);
  not g17757 (n_9840, n9918);
  not g17758 (n_9841, n9919);
  and g17759 (n9920, n_9840, n_9841);
  not g17760 (n_9842, n9869);
  not g17761 (n_9843, n9920);
  and g17762 (n9921, n_9842, n_9843);
  and g17763 (n9922, n_9832, n_9831);
  and g17764 (n9923, n_9785, n_9833);
  not g17765 (n_9844, n9922);
  and g17766 (n9924, n_9844, n9923);
  not g17767 (n_9845, n9923);
  and g17768 (n9925, n9922, n_9845);
  not g17769 (n_9846, n9924);
  not g17770 (n_9847, n9925);
  and g17771 (n9926, n_9846, n_9847);
  and g17772 (n9927, n_9731, n_9730);
  and g17773 (n9928, n_9684, n_9732);
  not g17774 (n_9848, n9927);
  and g17775 (n9929, n_9848, n9928);
  not g17776 (n_9849, n9928);
  and g17777 (n9930, n9927, n_9849);
  not g17778 (n_9850, n9929);
  not g17779 (n_9851, n9930);
  and g17780 (n9931, n_9850, n_9851);
  not g17781 (n_9852, n9926);
  not g17782 (n_9853, n9931);
  and g17783 (n9932, n_9852, n_9853);
  not g17784 (n_9854, n9921);
  not g17785 (n_9855, n9932);
  and g17786 (n9933, n_9854, n_9855);
  not g17787 (n_9856, n9917);
  and g17788 (n9934, n_9856, n9933);
  and g17789 (n9935, n_9856, n_9854);
  not g17790 (n_9857, n9935);
  and g17791 (n9936, n9932, n_9857);
  not g17792 (n_9858, n9934);
  not g17793 (n_9859, n9936);
  and g17794 (n9937, n_9858, n_9859);
  not g17795 (n_9860, n9833);
  not g17796 (n_9861, n9937);
  and g17797 (n9938, n_9860, n_9861);
  and g17798 (n9939, n_9854, n9932);
  and g17799 (n9940, n_9856, n9939);
  and g17800 (n9941, n_9855, n_9857);
  not g17801 (n_9862, n9940);
  not g17802 (n_9863, n9941);
  and g17803 (n9942, n_9862, n_9863);
  not g17804 (n_9864, n9942);
  and g17805 (n9943, n9833, n_9864);
  and g17806 (n9944, n_9852, n9931);
  and g17807 (n9945, n9926, n_9853);
  not g17808 (n_9865, n9944);
  not g17809 (n_9866, n9945);
  and g17810 (n9946, n_9865, n_9866);
  and g17811 (n9947, n_9616, n9712);
  and g17812 (n9948, n9637, n_9617);
  not g17813 (n_9867, n9947);
  not g17814 (n_9868, n9948);
  and g17815 (n9949, n_9867, n_9868);
  not g17816 (n_9869, n9946);
  not g17817 (n_9870, n9949);
  and g17818 (n9950, n_9869, n_9870);
  not g17819 (n_9871, n9943);
  not g17820 (n_9872, n9950);
  and g17821 (n9951, n_9871, n_9872);
  not g17822 (n_9873, n9938);
  and g17823 (n9952, n_9873, n9951);
  and g17824 (n9953, n_9873, n_9871);
  not g17825 (n_9874, n9953);
  and g17826 (n9954, n9950, n_9874);
  not g17827 (n_9875, n9952);
  not g17828 (n_9876, n9954);
  and g17829 (n9955, n_9875, n_9876);
  not g17830 (n_9877, n9744);
  not g17831 (n_9878, n9955);
  and g17832 (n9956, n_9877, n_9878);
  and g17833 (n9957, n_9871, n9950);
  and g17834 (n9958, n_9873, n9957);
  and g17835 (n9959, n_9872, n_9874);
  not g17836 (n_9879, n9958);
  not g17837 (n_9880, n9959);
  and g17838 (n9960, n_9879, n_9880);
  not g17839 (n_9881, n9960);
  and g17840 (n9961, n9744, n_9881);
  and g17841 (n9962, n_9869, n9949);
  and g17842 (n9963, n9946, n_9870);
  not g17843 (n_9882, n9962);
  not g17844 (n_9883, n9963);
  and g17845 (n9964, n_9882, n_9883);
  and g17846 (n9965, n_9369, n9481);
  and g17847 (n9966, n9328, n_9370);
  not g17848 (n_9884, n9965);
  not g17849 (n_9885, n9966);
  and g17850 (n9967, n_9884, n_9885);
  not g17851 (n_9886, n9964);
  not g17852 (n_9887, n9967);
  and g17853 (n9968, n_9886, n_9887);
  not g17854 (n_9888, n9961);
  not g17855 (n_9889, n9968);
  and g17856 (n9969, n_9888, n_9889);
  not g17857 (n_9890, n9956);
  and g17858 (n9970, n_9890, n9969);
  and g17859 (n9971, n_9890, n_9888);
  not g17860 (n_9891, n9971);
  and g17861 (n9972, n9968, n_9891);
  not g17862 (n_9892, n9970);
  not g17863 (n_9893, n9972);
  and g17864 (n9973, n_9892, n_9893);
  not g17865 (n_9894, n9544);
  not g17866 (n_9895, n9973);
  and g17867 (n9974, n_9894, n_9895);
  and g17868 (n9975, n_9888, n9968);
  and g17869 (n9976, n_9890, n9975);
  and g17870 (n9977, n_9889, n_9891);
  not g17871 (n_9896, n9976);
  not g17872 (n_9897, n9977);
  and g17873 (n9978, n_9896, n_9897);
  not g17874 (n_9898, n9978);
  and g17875 (n9979, n9544, n_9898);
  and g17876 (n9980, n_9886, n9967);
  and g17877 (n9981, n9964, n_9887);
  not g17878 (n_9899, n9980);
  not g17879 (n_9900, n9981);
  and g17880 (n9982, n_9899, n_9900);
  and g17881 (n9983, n_8858, n9001);
  and g17882 (n9984, n8692, n_8859);
  not g17883 (n_9901, n9983);
  not g17884 (n_9902, n9984);
  and g17885 (n9985, n_9901, n_9902);
  not g17886 (n_9903, n9982);
  not g17887 (n_9904, n9985);
  and g17888 (n9986, n_9903, n_9904);
  not g17889 (n_9905, n9979);
  not g17890 (n_9906, n9986);
  and g17891 (n9987, n_9905, n_9906);
  not g17892 (n_9907, n9974);
  and g17893 (n9988, n_9907, n9987);
  and g17894 (n9989, n_9907, n_9905);
  not g17895 (n_9908, n9989);
  and g17896 (n9990, n9986, n_9908);
  not g17897 (n_9909, n9988);
  not g17898 (n_9910, n9990);
  and g17899 (n9991, n_9909, n_9910);
  not g17900 (n_9911, n9126);
  not g17901 (n_9912, n9991);
  and g17902 (n9992, n_9911, n_9912);
  and g17903 (n9993, n_9905, n9986);
  and g17904 (n9994, n_9907, n9993);
  and g17905 (n9995, n_9906, n_9908);
  not g17906 (n_9913, n9994);
  not g17907 (n_9914, n9995);
  and g17908 (n9996, n_9913, n_9914);
  not g17909 (n_9915, n9996);
  and g17910 (n9997, n9126, n_9915);
  and g17911 (n9998, n_9903, n9985);
  and g17912 (n9999, n9982, n_9904);
  not g17913 (n_9916, n9998);
  not g17914 (n_9917, n9999);
  and g17915 (n10000, n_9916, n_9917);
  and g17916 (n10001, n_7819, n8023);
  and g17917 (n10002, n7402, n_7820);
  not g17918 (n_9918, n10001);
  not g17919 (n_9919, n10002);
  and g17920 (n10003, n_9918, n_9919);
  not g17921 (n_9920, n10000);
  not g17922 (n_9921, n10003);
  and g17923 (n10004, n_9920, n_9921);
  not g17924 (n_9922, n9997);
  not g17925 (n_9923, n10004);
  and g17926 (n10005, n_9922, n_9923);
  not g17927 (n_9924, n9992);
  and g17928 (n10006, n_9924, n10005);
  and g17929 (n10007, n_9924, n_9922);
  not g17930 (n_9925, n10007);
  and g17931 (n10008, n10004, n_9925);
  not g17932 (n_9926, n10006);
  not g17933 (n_9927, n10008);
  and g17934 (n10009, n_9926, n_9927);
  not g17935 (n_9928, n8272);
  not g17936 (n_9929, n10009);
  and g17937 (n10010, n_9928, n_9929);
  and g17938 (n10011, n_9922, n10004);
  and g17939 (n10012, n_9924, n10011);
  and g17940 (n10013, n_9923, n_9925);
  not g17941 (n_9930, n10012);
  not g17942 (n_9931, n10013);
  and g17943 (n10014, n_9930, n_9931);
  not g17944 (n_9932, n10014);
  and g17945 (n10015, n8272, n_9932);
  and g17946 (n10016, n_9920, n10003);
  and g17947 (n10017, n10000, n_9921);
  not g17948 (n_9933, n10016);
  not g17949 (n_9934, n10017);
  and g17950 (n10018, n_9933, n_9934);
  and g17951 (n10019, n_5916, n6297);
  and g17952 (n10020, n_5150, n_5917);
  and g17953 (n10021, n_5151, n10020);
  not g17954 (n_9935, n10019);
  not g17955 (n_9936, n10021);
  and g17956 (n10022, n_9935, n_9936);
  not g17957 (n_9937, n10018);
  not g17958 (n_9938, n10022);
  and g17959 (n10023, n_9937, n_9938);
  not g17960 (n_9939, n10015);
  not g17961 (n_9940, n10023);
  and g17962 (n10024, n_9939, n_9940);
  not g17963 (n_9941, n10010);
  and g17964 (n10025, n_9941, n10024);
  and g17965 (n10026, n_9941, n_9939);
  not g17966 (n_9942, n10026);
  and g17967 (n10027, n10023, n_9942);
  not g17968 (n_9943, n10025);
  not g17969 (n_9944, n10027);
  and g17970 (n10028, n_9943, n_9944);
  not g17971 (n_9945, n6546);
  not g17972 (n_9946, n10028);
  and g17973 (n10029, n_9945, n_9946);
  and g17974 (n10030, n_3436, n3975);
  and g17975 (n10031, n3972, n_3437);
  not g17976 (n_9947, n10030);
  not g17977 (n_9948, n10031);
  and g17978 (n10032, n_9947, n_9948);
  and g17979 (n10033, n_9937, n10022);
  and g17980 (n10034, n10018, n_9938);
  not g17981 (n_9949, n10033);
  not g17982 (n_9950, n10034);
  and g17983 (n10035, n_9949, n_9950);
  not g17984 (n_9951, n10032);
  not g17985 (n_9952, n10035);
  and g17986 (n10036, n_9951, n_9952);
  and g17987 (n10037, n_9939, n10023);
  and g17988 (n10038, n_9941, n10037);
  and g17989 (n10039, n_9940, n_9942);
  not g17990 (n_9953, n10038);
  not g17991 (n_9954, n10039);
  and g17992 (n10040, n_9953, n_9954);
  not g17993 (n_9955, n10040);
  and g17994 (n10041, n6546, n_9955);
  not g17995 (n_9956, n10036);
  not g17996 (n_9957, n10041);
  and g17997 (n10042, n_9956, n_9957);
  not g17998 (n_9958, n10029);
  and g17999 (n10043, n_9958, n10042);
  not g18000 (n_9959, n4472);
  not g18001 (n_9960, n10043);
  and g18002 (n10044, n_9959, n_9960);
  and g18003 (n10045, n_9958, n_9957);
  not g18004 (n_9961, n10045);
  and g18005 (n10046, n10036, n_9961);
  not g18006 (n_9962, n10044);
  not g18007 (n_9963, n10046);
  and g18008 (n10047, n_9962, n_9963);
  and g18009 (n10048, n_9945, n_9943);
  not g18010 (n_9964, n10048);
  and g18011 (n10049, n_9944, n_9964);
  and g18012 (n10050, n_6108, n_6106);
  not g18013 (n_9965, n10050);
  and g18014 (n10051, n_6107, n_9965);
  and g18015 (n10052, n_5145, n_5143);
  not g18016 (n_9966, n10052);
  and g18017 (n10053, n_5144, n_9966);
  and g18018 (n10054, n_5128, n_5126);
  not g18019 (n_9967, n10054);
  and g18020 (n10055, n_5127, n_9967);
  and g18021 (n10056, n_4651, n_4649);
  not g18022 (n_9968, n10056);
  and g18023 (n10057, n_4650, n_9968);
  and g18024 (n10058, n5172, n_4643);
  not g18025 (n_9969, n10058);
  and g18026 (n10059, n_4644, n_9969);
  and g18027 (n10060, n_4633, n_4631);
  not g18028 (n_9970, n10060);
  and g18029 (n10061, n_4632, n_9970);
  and g18030 (n10062, n_4617, n_4618);
  not g18031 (n_9971, n10062);
  and g18032 (n10063, n_4626, n_9971);
  not g18033 (n_9972, n10061);
  and g18034 (n10064, n_9972, n10063);
  not g18035 (n_9973, n10063);
  and g18036 (n10065, n_4632, n_9973);
  and g18037 (n10066, n_9970, n10065);
  and g18038 (n10067, n_4552, n_4551);
  not g18039 (n_9974, n10067);
  and g18040 (n10068, n_4550, n_9974);
  not g18041 (n_9975, n10066);
  and g18042 (n10069, n_9975, n10068);
  not g18043 (n_9976, n10064);
  and g18044 (n10070, n_9976, n10069);
  and g18045 (n10071, n_9976, n_9975);
  not g18046 (n_9977, n10068);
  not g18047 (n_9978, n10071);
  and g18048 (n10072, n_9977, n_9978);
  not g18049 (n_9979, n10070);
  not g18050 (n_9980, n10072);
  and g18051 (n10073, n_9979, n_9980);
  not g18052 (n_9981, n10059);
  not g18053 (n_9982, n10073);
  and g18054 (n10074, n_9981, n_9982);
  not g18058 (n_9983, n10074);
  not g18059 (n_9984, n10077);
  and g18060 (n10078, n_9983, n_9984);
  and g18061 (n10079, n_4503, n_4501);
  not g18062 (n_9985, n10079);
  and g18063 (n10080, n_4502, n_9985);
  and g18064 (n10081, n4926, n_4383);
  not g18065 (n_9986, n10081);
  and g18066 (n10082, n_4384, n_9986);
  and g18067 (n10083, n_4370, n_4373);
  not g18068 (n_9987, n10083);
  and g18069 (n10084, n_4369, n_9987);
  and g18070 (n10085, n_4329, n_4327);
  not g18071 (n_9988, n10085);
  and g18072 (n10086, n_4328, n_9988);
  not g18073 (n_9989, n10084);
  and g18074 (n10087, n_9989, n10086);
  not g18075 (n_9990, n10086);
  and g18076 (n10088, n10084, n_9990);
  not g18077 (n_9991, n10087);
  not g18078 (n_9992, n10088);
  and g18079 (n10089, n_9991, n_9992);
  not g18080 (n_9993, n10082);
  not g18081 (n_9994, n10089);
  and g18082 (n10090, n_9993, n_9994);
  not g18086 (n_9995, n10090);
  not g18087 (n_9996, n10093);
  and g18088 (n10094, n_9995, n_9996);
  and g18089 (n10095, n5015, n_4480);
  not g18090 (n_9997, n10095);
  and g18091 (n10096, n_4481, n_9997);
  and g18092 (n10097, n_4471, n_4474);
  not g18093 (n_9998, n10097);
  and g18094 (n10098, n_4470, n_9998);
  and g18095 (n10099, n_4430, n_4428);
  not g18096 (n_9999, n10099);
  and g18097 (n10100, n_4429, n_9999);
  not g18098 (n_10000, n10098);
  and g18099 (n10101, n_10000, n10100);
  not g18100 (n_10001, n10100);
  and g18101 (n10102, n10098, n_10001);
  not g18102 (n_10002, n10101);
  not g18103 (n_10003, n10102);
  and g18104 (n10103, n_10002, n_10003);
  not g18105 (n_10004, n10096);
  not g18106 (n_10005, n10103);
  and g18107 (n10104, n_10004, n_10005);
  not g18111 (n_10006, n10104);
  not g18112 (n_10007, n10107);
  and g18113 (n10108, n_10006, n_10007);
  not g18114 (n_10008, n10094);
  and g18115 (n10109, n_10008, n10108);
  not g18116 (n_10009, n10108);
  and g18117 (n10110, n10094, n_10009);
  not g18118 (n_10010, n10109);
  not g18119 (n_10011, n10110);
  and g18120 (n10111, n_10010, n_10011);
  not g18121 (n_10012, n10080);
  not g18122 (n_10013, n10111);
  and g18123 (n10112, n_10012, n_10013);
  and g18124 (n10113, n10080, n10111);
  not g18125 (n_10014, n10112);
  not g18126 (n_10015, n10113);
  and g18127 (n10114, n_10014, n_10015);
  not g18128 (n_10016, n10078);
  and g18129 (n10115, n_10016, n10114);
  not g18130 (n_10017, n10114);
  and g18131 (n10116, n10078, n_10017);
  not g18132 (n_10018, n10115);
  not g18133 (n_10019, n10116);
  and g18134 (n10117, n_10018, n_10019);
  not g18135 (n_10020, n10057);
  not g18136 (n_10021, n10117);
  and g18137 (n10118, n_10020, n_10021);
  and g18138 (n10119, n10057, n10117);
  not g18139 (n_10022, n10118);
  not g18140 (n_10023, n10119);
  and g18141 (n10120, n_10022, n_10023);
  and g18142 (n10121, n_5111, n_5109);
  not g18143 (n_10024, n10121);
  and g18144 (n10122, n_5110, n_10024);
  and g18145 (n10123, n_4874, n_4872);
  not g18146 (n_10025, n10123);
  and g18147 (n10124, n_4873, n_10025);
  and g18148 (n10125, n5394, n_4866);
  not g18149 (n_10026, n10125);
  and g18150 (n10126, n_4867, n_10026);
  and g18151 (n10127, n_4800, n_4799);
  not g18152 (n_10027, n10127);
  and g18153 (n10128, n_4798, n_10027);
  and g18154 (n10129, n_4844, n_4843);
  not g18155 (n_10028, n10129);
  and g18156 (n10130, n_4842, n_10028);
  not g18157 (n_10029, n10128);
  and g18158 (n10131, n_10029, n10130);
  not g18159 (n_10030, n10130);
  and g18160 (n10132, n10128, n_10030);
  not g18161 (n_10031, n10131);
  not g18162 (n_10032, n10132);
  and g18163 (n10133, n_10031, n_10032);
  not g18164 (n_10033, n10126);
  not g18165 (n_10034, n10133);
  and g18166 (n10134, n_10033, n_10034);
  not g18170 (n_10035, n10134);
  not g18171 (n_10036, n10137);
  and g18172 (n10138, n_10035, n_10036);
  and g18173 (n10139, n5254, n_4747);
  not g18174 (n_10037, n10139);
  and g18175 (n10140, n_4748, n_10037);
  and g18176 (n10141, n_4738, n_4741);
  not g18177 (n_10038, n10141);
  and g18178 (n10142, n_4737, n_10038);
  and g18179 (n10143, n_4697, n_4695);
  not g18180 (n_10039, n10143);
  and g18181 (n10144, n_4696, n_10039);
  not g18182 (n_10040, n10142);
  and g18183 (n10145, n_10040, n10144);
  not g18184 (n_10041, n10144);
  and g18185 (n10146, n10142, n_10041);
  not g18186 (n_10042, n10145);
  not g18187 (n_10043, n10146);
  and g18188 (n10147, n_10042, n_10043);
  not g18189 (n_10044, n10140);
  not g18190 (n_10045, n10147);
  and g18191 (n10148, n_10044, n_10045);
  not g18195 (n_10046, n10148);
  not g18196 (n_10047, n10151);
  and g18197 (n10152, n_10046, n_10047);
  not g18198 (n_10048, n10138);
  and g18199 (n10153, n_10048, n10152);
  not g18200 (n_10049, n10152);
  and g18201 (n10154, n10138, n_10049);
  not g18202 (n_10050, n10153);
  not g18203 (n_10051, n10154);
  and g18204 (n10155, n_10050, n_10051);
  not g18205 (n_10052, n10124);
  not g18206 (n_10053, n10155);
  and g18207 (n10156, n_10052, n_10053);
  and g18208 (n10157, n10124, n10155);
  not g18209 (n_10054, n10156);
  not g18210 (n_10055, n10157);
  and g18211 (n10158, n_10054, n_10055);
  and g18212 (n10159, n_5094, n_5092);
  not g18213 (n_10056, n10159);
  and g18214 (n10160, n_5093, n_10056);
  and g18215 (n10161, n5454, n_4974);
  not g18216 (n_10057, n10161);
  and g18217 (n10162, n_4975, n_10057);
  and g18218 (n10163, n_4961, n_4964);
  not g18219 (n_10058, n10163);
  and g18220 (n10164, n_4960, n_10058);
  and g18221 (n10165, n_4920, n_4918);
  not g18222 (n_10059, n10165);
  and g18223 (n10166, n_4919, n_10059);
  not g18224 (n_10060, n10164);
  and g18225 (n10167, n_10060, n10166);
  not g18226 (n_10061, n10166);
  and g18227 (n10168, n10164, n_10061);
  not g18228 (n_10062, n10167);
  not g18229 (n_10063, n10168);
  and g18230 (n10169, n_10062, n_10063);
  not g18231 (n_10064, n10162);
  not g18232 (n_10065, n10169);
  and g18233 (n10170, n_10064, n_10065);
  not g18237 (n_10066, n10170);
  not g18238 (n_10067, n10173);
  and g18239 (n10174, n_10066, n_10067);
  and g18240 (n10175, n5543, n_5071);
  not g18241 (n_10068, n10175);
  and g18242 (n10176, n_5072, n_10068);
  and g18243 (n10177, n_5062, n_5065);
  not g18244 (n_10069, n10177);
  and g18245 (n10178, n_5061, n_10069);
  and g18246 (n10179, n_5021, n_5019);
  not g18247 (n_10070, n10179);
  and g18248 (n10180, n_5020, n_10070);
  not g18249 (n_10071, n10178);
  and g18250 (n10181, n_10071, n10180);
  not g18251 (n_10072, n10180);
  and g18252 (n10182, n10178, n_10072);
  not g18253 (n_10073, n10181);
  not g18254 (n_10074, n10182);
  and g18255 (n10183, n_10073, n_10074);
  not g18256 (n_10075, n10176);
  not g18257 (n_10076, n10183);
  and g18258 (n10184, n_10075, n_10076);
  not g18262 (n_10077, n10184);
  not g18263 (n_10078, n10187);
  and g18264 (n10188, n_10077, n_10078);
  not g18265 (n_10079, n10174);
  and g18266 (n10189, n_10079, n10188);
  not g18267 (n_10080, n10188);
  and g18268 (n10190, n10174, n_10080);
  not g18269 (n_10081, n10189);
  not g18270 (n_10082, n10190);
  and g18271 (n10191, n_10081, n_10082);
  not g18272 (n_10083, n10160);
  not g18273 (n_10084, n10191);
  and g18274 (n10192, n_10083, n_10084);
  and g18275 (n10193, n10160, n10191);
  not g18276 (n_10085, n10192);
  not g18277 (n_10086, n10193);
  and g18278 (n10194, n_10085, n_10086);
  not g18279 (n_10087, n10158);
  and g18280 (n10195, n_10087, n10194);
  not g18281 (n_10088, n10194);
  and g18282 (n10196, n10158, n_10088);
  not g18283 (n_10089, n10195);
  not g18284 (n_10090, n10196);
  and g18285 (n10197, n_10089, n_10090);
  not g18286 (n_10091, n10122);
  not g18287 (n_10092, n10197);
  and g18288 (n10198, n_10091, n_10092);
  and g18289 (n10199, n10122, n10197);
  not g18290 (n_10093, n10198);
  not g18291 (n_10094, n10199);
  and g18292 (n10200, n_10093, n_10094);
  not g18293 (n_10095, n10120);
  and g18294 (n10201, n_10095, n10200);
  not g18295 (n_10096, n10200);
  and g18296 (n10202, n10120, n_10096);
  not g18297 (n_10097, n10201);
  not g18298 (n_10098, n10202);
  and g18299 (n10203, n_10097, n_10098);
  and g18300 (n10204, n10055, n10203);
  not g18301 (n_10099, n10055);
  not g18302 (n_10100, n10203);
  and g18303 (n10205, n_10099, n_10100);
  and g18304 (n10206, n_4283, n_4281);
  not g18305 (n_10101, n10206);
  and g18306 (n10207, n_4282, n_10101);
  and g18307 (n10208, n_4276, n_4274);
  not g18308 (n_10102, n10208);
  and g18309 (n10209, n_4275, n_10102);
  and g18310 (n10210, n4859, n_4268);
  not g18311 (n_10103, n10210);
  and g18312 (n10211, n_4269, n_10103);
  and g18313 (n10212, n_4181, n_4180);
  not g18314 (n_10104, n10212);
  and g18315 (n10213, n_4179, n_10104);
  and g18316 (n10214, n_4225, n_4224);
  not g18317 (n_10105, n10214);
  and g18318 (n10215, n_4223, n_10105);
  not g18319 (n_10106, n10213);
  and g18320 (n10216, n_10106, n10215);
  not g18321 (n_10107, n10215);
  and g18322 (n10217, n10213, n_10107);
  not g18323 (n_10108, n10216);
  not g18324 (n_10109, n10217);
  and g18325 (n10218, n_10108, n_10109);
  not g18326 (n_10110, n10211);
  not g18327 (n_10111, n10218);
  and g18328 (n10219, n_10110, n_10111);
  not g18332 (n_10112, n10219);
  not g18333 (n_10113, n10222);
  and g18334 (n10223, n_10112, n_10113);
  and g18335 (n10224, n4835, n_4247);
  not g18336 (n_10114, n10224);
  and g18337 (n10225, n_4248, n_10114);
  and g18338 (n10226, n_4089, n_4088);
  not g18339 (n_10115, n10226);
  and g18340 (n10227, n_4087, n_10115);
  and g18341 (n10228, n_4133, n_4132);
  not g18342 (n_10116, n10228);
  and g18343 (n10229, n_4131, n_10116);
  not g18344 (n_10117, n10227);
  and g18345 (n10230, n_10117, n10229);
  not g18346 (n_10118, n10229);
  and g18347 (n10231, n10227, n_10118);
  not g18348 (n_10119, n10230);
  not g18349 (n_10120, n10231);
  and g18350 (n10232, n_10119, n_10120);
  not g18351 (n_10121, n10225);
  not g18352 (n_10122, n10232);
  and g18353 (n10233, n_10121, n_10122);
  not g18357 (n_10123, n10233);
  not g18358 (n_10124, n10236);
  and g18359 (n10237, n_10123, n_10124);
  not g18360 (n_10125, n10223);
  and g18361 (n10238, n_10125, n10237);
  not g18362 (n_10126, n10237);
  and g18363 (n10239, n10223, n_10126);
  not g18364 (n_10127, n10238);
  not g18365 (n_10128, n10239);
  and g18366 (n10240, n_10127, n_10128);
  not g18367 (n_10129, n10209);
  not g18368 (n_10130, n10240);
  and g18369 (n10241, n_10129, n_10130);
  and g18370 (n10242, n10209, n10240);
  not g18371 (n_10131, n10241);
  not g18372 (n_10132, n10242);
  and g18373 (n10243, n_10131, n_10132);
  and g18374 (n10244, n_4040, n_4038);
  not g18375 (n_10133, n10244);
  and g18376 (n10245, n_4039, n_10133);
  and g18377 (n10246, n4508, n_3920);
  not g18378 (n_10134, n10246);
  and g18379 (n10247, n_3921, n_10134);
  and g18380 (n10248, n_3907, n_3910);
  not g18381 (n_10135, n10248);
  and g18382 (n10249, n_3906, n_10135);
  and g18383 (n10250, n_3866, n_3864);
  not g18384 (n_10136, n10250);
  and g18385 (n10251, n_3865, n_10136);
  not g18386 (n_10137, n10249);
  and g18387 (n10252, n_10137, n10251);
  not g18388 (n_10138, n10251);
  and g18389 (n10253, n10249, n_10138);
  not g18390 (n_10139, n10252);
  not g18391 (n_10140, n10253);
  and g18392 (n10254, n_10139, n_10140);
  not g18393 (n_10141, n10247);
  not g18394 (n_10142, n10254);
  and g18395 (n10255, n_10141, n_10142);
  not g18399 (n_10143, n10255);
  not g18400 (n_10144, n10258);
  and g18401 (n10259, n_10143, n_10144);
  and g18402 (n10260, n4597, n_4017);
  not g18403 (n_10145, n10260);
  and g18404 (n10261, n_4018, n_10145);
  and g18405 (n10262, n_4008, n_4011);
  not g18406 (n_10146, n10262);
  and g18407 (n10263, n_4007, n_10146);
  and g18408 (n10264, n_3967, n_3965);
  not g18409 (n_10147, n10264);
  and g18410 (n10265, n_3966, n_10147);
  not g18411 (n_10148, n10263);
  and g18412 (n10266, n_10148, n10265);
  not g18413 (n_10149, n10265);
  and g18414 (n10267, n10263, n_10149);
  not g18415 (n_10150, n10266);
  not g18416 (n_10151, n10267);
  and g18417 (n10268, n_10150, n_10151);
  not g18418 (n_10152, n10261);
  not g18419 (n_10153, n10268);
  and g18420 (n10269, n_10152, n_10153);
  not g18424 (n_10154, n10269);
  not g18425 (n_10155, n10272);
  and g18426 (n10273, n_10154, n_10155);
  not g18427 (n_10156, n10259);
  and g18428 (n10274, n_10156, n10273);
  not g18429 (n_10157, n10273);
  and g18430 (n10275, n10259, n_10157);
  not g18431 (n_10158, n10274);
  not g18432 (n_10159, n10275);
  and g18433 (n10276, n_10158, n_10159);
  not g18434 (n_10160, n10245);
  not g18435 (n_10161, n10276);
  and g18436 (n10277, n_10160, n_10161);
  and g18437 (n10278, n10245, n10276);
  not g18438 (n_10162, n10277);
  not g18439 (n_10163, n10278);
  and g18440 (n10279, n_10162, n_10163);
  not g18441 (n_10164, n10243);
  and g18442 (n10280, n_10164, n10279);
  not g18443 (n_10165, n10279);
  and g18444 (n10281, n10243, n_10165);
  not g18445 (n_10166, n10280);
  not g18446 (n_10167, n10281);
  and g18447 (n10282, n_10166, n_10167);
  not g18448 (n_10168, n10207);
  not g18449 (n_10169, n10282);
  and g18450 (n10283, n_10168, n_10169);
  and g18451 (n10284, n10207, n10282);
  not g18452 (n_10170, n10283);
  not g18453 (n_10171, n10284);
  and g18454 (n10285, n_10170, n_10171);
  not g18455 (n_10172, n10205);
  not g18456 (n_10173, n10285);
  and g18457 (n10286, n_10172, n_10173);
  not g18458 (n_10174, n10204);
  and g18459 (n10287, n_10174, n10286);
  and g18460 (n10288, n_10174, n_10172);
  not g18461 (n_10175, n10288);
  and g18462 (n10289, n10285, n_10175);
  not g18463 (n_10176, n10287);
  not g18464 (n_10177, n10289);
  and g18465 (n10290, n_10176, n_10177);
  and g18466 (n10291, n10053, n10290);
  not g18467 (n_10178, n10053);
  not g18468 (n_10179, n10290);
  and g18469 (n10292, n_10178, n_10179);
  and g18470 (n10293, n_6101, n_6099);
  not g18471 (n_10180, n10293);
  and g18472 (n10294, n_6100, n_10180);
  and g18473 (n10295, n_6094, n_6092);
  not g18474 (n_10181, n10295);
  and g18475 (n10296, n_6093, n_10181);
  and g18476 (n10297, n_6087, n_6085);
  not g18477 (n_10182, n10297);
  and g18478 (n10298, n_6086, n_10182);
  and g18479 (n10299, n6501, n_6079);
  not g18480 (n_10183, n10299);
  and g18481 (n10300, n_6080, n_10183);
  and g18482 (n10301, n_5854, n_5853);
  not g18483 (n_10184, n10301);
  and g18484 (n10302, n_5852, n_10184);
  and g18485 (n10303, n_5898, n_5897);
  not g18486 (n_10185, n10303);
  and g18487 (n10304, n_5896, n_10185);
  not g18488 (n_10186, n10302);
  and g18489 (n10305, n_10186, n10304);
  not g18490 (n_10187, n10304);
  and g18491 (n10306, n10302, n_10187);
  not g18492 (n_10188, n10305);
  not g18493 (n_10189, n10306);
  and g18494 (n10307, n_10188, n_10189);
  not g18495 (n_10190, n10300);
  not g18496 (n_10191, n10307);
  and g18497 (n10308, n_10190, n_10191);
  not g18501 (n_10192, n10308);
  not g18502 (n_10193, n10311);
  and g18503 (n10312, n_10192, n_10193);
  and g18504 (n10313, n6477, n_6058);
  not g18505 (n_10194, n10313);
  and g18506 (n10314, n_6059, n_10194);
  and g18507 (n10315, n_5762, n_5761);
  not g18508 (n_10195, n10315);
  and g18509 (n10316, n_5760, n_10195);
  and g18510 (n10317, n_5806, n_5805);
  not g18511 (n_10196, n10317);
  and g18512 (n10318, n_5804, n_10196);
  not g18513 (n_10197, n10316);
  and g18514 (n10319, n_10197, n10318);
  not g18515 (n_10198, n10318);
  and g18516 (n10320, n10316, n_10198);
  not g18517 (n_10199, n10319);
  not g18518 (n_10200, n10320);
  and g18519 (n10321, n_10199, n_10200);
  not g18520 (n_10201, n10314);
  not g18521 (n_10202, n10321);
  and g18522 (n10322, n_10201, n_10202);
  not g18526 (n_10203, n10322);
  not g18527 (n_10204, n10325);
  and g18528 (n10326, n_10203, n_10204);
  not g18529 (n_10205, n10312);
  and g18530 (n10327, n_10205, n10326);
  not g18531 (n_10206, n10326);
  and g18532 (n10328, n10312, n_10206);
  not g18533 (n_10207, n10327);
  not g18534 (n_10208, n10328);
  and g18535 (n10329, n_10207, n_10208);
  not g18536 (n_10209, n10298);
  not g18537 (n_10210, n10329);
  and g18538 (n10330, n_10209, n_10210);
  and g18539 (n10331, n10298, n10329);
  not g18540 (n_10211, n10330);
  not g18541 (n_10212, n10331);
  and g18542 (n10332, n_10211, n_10212);
  and g18543 (n10333, n_6043, n_6041);
  not g18544 (n_10213, n10333);
  and g18545 (n10334, n_6042, n_10213);
  and g18546 (n10335, n6422, n_6021);
  not g18547 (n_10214, n10335);
  and g18548 (n10336, n_6022, n_10214);
  and g18549 (n10337, n_5666, n_5665);
  not g18550 (n_10215, n10337);
  and g18551 (n10338, n_5664, n_10215);
  and g18552 (n10339, n_5710, n_5709);
  not g18553 (n_10216, n10339);
  and g18554 (n10340, n_5708, n_10216);
  not g18555 (n_10217, n10338);
  and g18556 (n10341, n_10217, n10340);
  not g18557 (n_10218, n10340);
  and g18558 (n10342, n10338, n_10218);
  not g18559 (n_10219, n10341);
  not g18560 (n_10220, n10342);
  and g18561 (n10343, n_10219, n_10220);
  not g18562 (n_10221, n10336);
  not g18563 (n_10222, n10343);
  and g18564 (n10344, n_10221, n_10222);
  not g18568 (n_10223, n10344);
  not g18569 (n_10224, n10347);
  and g18570 (n10348, n_10223, n_10224);
  and g18571 (n10349, n6441, n_6030);
  not g18572 (n_10225, n10349);
  and g18573 (n10350, n_6031, n_10225);
  and g18574 (n10351, n_5574, n_5573);
  not g18575 (n_10226, n10351);
  and g18576 (n10352, n_5572, n_10226);
  and g18577 (n10353, n_5618, n_5617);
  not g18578 (n_10227, n10353);
  and g18579 (n10354, n_5616, n_10227);
  not g18580 (n_10228, n10352);
  and g18581 (n10355, n_10228, n10354);
  not g18582 (n_10229, n10354);
  and g18583 (n10356, n10352, n_10229);
  not g18584 (n_10230, n10355);
  not g18585 (n_10231, n10356);
  and g18586 (n10357, n_10230, n_10231);
  not g18587 (n_10232, n10350);
  not g18588 (n_10233, n10357);
  and g18589 (n10358, n_10232, n_10233);
  not g18593 (n_10234, n10358);
  not g18594 (n_10235, n10361);
  and g18595 (n10362, n_10234, n_10235);
  not g18596 (n_10236, n10348);
  and g18597 (n10363, n_10236, n10362);
  not g18598 (n_10237, n10362);
  and g18599 (n10364, n10348, n_10237);
  not g18600 (n_10238, n10363);
  not g18601 (n_10239, n10364);
  and g18602 (n10365, n_10238, n_10239);
  not g18603 (n_10240, n10334);
  not g18604 (n_10241, n10365);
  and g18605 (n10366, n_10240, n_10241);
  and g18606 (n10367, n10334, n10365);
  not g18607 (n_10242, n10366);
  not g18608 (n_10243, n10367);
  and g18609 (n10368, n_10242, n_10243);
  not g18610 (n_10244, n10332);
  and g18611 (n10369, n_10244, n10368);
  not g18612 (n_10245, n10368);
  and g18613 (n10370, n10332, n_10245);
  not g18614 (n_10246, n10369);
  not g18615 (n_10247, n10370);
  and g18616 (n10371, n_10246, n_10247);
  not g18617 (n_10248, n10296);
  not g18618 (n_10249, n10371);
  and g18619 (n10372, n_10248, n_10249);
  and g18620 (n10373, n10296, n10371);
  not g18621 (n_10250, n10372);
  not g18622 (n_10251, n10373);
  and g18623 (n10374, n_10250, n_10251);
  and g18624 (n10375, n_6002, n_6000);
  not g18625 (n_10252, n10375);
  and g18626 (n10376, n_6001, n_10252);
  and g18627 (n10377, n_5957, n_5955);
  not g18628 (n_10253, n10377);
  and g18629 (n10378, n_5956, n_10253);
  and g18630 (n10379, n6329, n_5949);
  not g18631 (n_10254, n10379);
  and g18632 (n10380, n_5950, n_10254);
  and g18633 (n10381, n_5474, n_5473);
  not g18634 (n_10255, n10381);
  and g18635 (n10382, n_5472, n_10255);
  and g18636 (n10383, n_5518, n_5517);
  not g18637 (n_10256, n10383);
  and g18638 (n10384, n_5516, n_10256);
  not g18639 (n_10257, n10382);
  and g18640 (n10385, n_10257, n10384);
  not g18641 (n_10258, n10384);
  and g18642 (n10386, n10382, n_10258);
  not g18643 (n_10259, n10385);
  not g18644 (n_10260, n10386);
  and g18645 (n10387, n_10259, n_10260);
  not g18646 (n_10261, n10380);
  not g18647 (n_10262, n10387);
  and g18648 (n10388, n_10261, n_10262);
  not g18652 (n_10263, n10388);
  not g18653 (n_10264, n10391);
  and g18654 (n10392, n_10263, n_10264);
  and g18655 (n10393, n6305, n_5928);
  not g18656 (n_10265, n10393);
  and g18657 (n10394, n_5929, n_10265);
  and g18658 (n10395, n_5382, n_5381);
  not g18659 (n_10266, n10395);
  and g18660 (n10396, n_5380, n_10266);
  and g18661 (n10397, n_5426, n_5425);
  not g18662 (n_10267, n10397);
  and g18663 (n10398, n_5424, n_10267);
  not g18664 (n_10268, n10396);
  and g18665 (n10399, n_10268, n10398);
  not g18666 (n_10269, n10398);
  and g18667 (n10400, n10396, n_10269);
  not g18668 (n_10270, n10399);
  not g18669 (n_10271, n10400);
  and g18670 (n10401, n_10270, n_10271);
  not g18671 (n_10272, n10394);
  not g18672 (n_10273, n10401);
  and g18673 (n10402, n_10272, n_10273);
  not g18677 (n_10274, n10402);
  not g18678 (n_10275, n10405);
  and g18679 (n10406, n_10274, n_10275);
  not g18680 (n_10276, n10392);
  and g18681 (n10407, n_10276, n10406);
  not g18682 (n_10277, n10406);
  and g18683 (n10408, n10392, n_10277);
  not g18684 (n_10278, n10407);
  not g18685 (n_10279, n10408);
  and g18686 (n10409, n_10278, n_10279);
  not g18687 (n_10280, n10378);
  not g18688 (n_10281, n10409);
  and g18689 (n10410, n_10280, n_10281);
  and g18690 (n10411, n10378, n10409);
  not g18691 (n_10282, n10410);
  not g18692 (n_10283, n10411);
  and g18693 (n10412, n_10282, n_10283);
  and g18694 (n10413, n_5991, n_5989);
  not g18695 (n_10284, n10413);
  and g18696 (n10414, n_5990, n_10284);
  and g18697 (n10415, n6355, n_5969);
  not g18698 (n_10285, n10415);
  and g18699 (n10416, n_5970, n_10285);
  and g18700 (n10417, n_5286, n_5285);
  not g18701 (n_10286, n10417);
  and g18702 (n10418, n_5284, n_10286);
  and g18703 (n10419, n_5330, n_5329);
  not g18704 (n_10287, n10419);
  and g18705 (n10420, n_5328, n_10287);
  not g18706 (n_10288, n10418);
  and g18707 (n10421, n_10288, n10420);
  not g18708 (n_10289, n10420);
  and g18709 (n10422, n10418, n_10289);
  not g18710 (n_10290, n10421);
  not g18711 (n_10291, n10422);
  and g18712 (n10423, n_10290, n_10291);
  not g18713 (n_10292, n10416);
  not g18714 (n_10293, n10423);
  and g18715 (n10424, n_10292, n_10293);
  not g18719 (n_10294, n10424);
  not g18720 (n_10295, n10427);
  and g18721 (n10428, n_10294, n_10295);
  and g18722 (n10429, n6374, n_5978);
  not g18723 (n_10296, n10429);
  and g18724 (n10430, n_5979, n_10296);
  and g18725 (n10431, n_5194, n_5193);
  not g18726 (n_10297, n10431);
  and g18727 (n10432, n_5192, n_10297);
  and g18728 (n10433, n_5238, n_5237);
  not g18729 (n_10298, n10433);
  and g18730 (n10434, n_5236, n_10298);
  not g18731 (n_10299, n10432);
  and g18732 (n10435, n_10299, n10434);
  not g18733 (n_10300, n10434);
  and g18734 (n10436, n10432, n_10300);
  not g18735 (n_10301, n10435);
  not g18736 (n_10302, n10436);
  and g18737 (n10437, n_10301, n_10302);
  not g18738 (n_10303, n10430);
  not g18739 (n_10304, n10437);
  and g18740 (n10438, n_10303, n_10304);
  not g18744 (n_10305, n10438);
  not g18745 (n_10306, n10441);
  and g18746 (n10442, n_10305, n_10306);
  not g18747 (n_10307, n10428);
  and g18748 (n10443, n_10307, n10442);
  not g18749 (n_10308, n10442);
  and g18750 (n10444, n10428, n_10308);
  not g18751 (n_10309, n10443);
  not g18752 (n_10310, n10444);
  and g18753 (n10445, n_10309, n_10310);
  not g18754 (n_10311, n10414);
  not g18755 (n_10312, n10445);
  and g18756 (n10446, n_10311, n_10312);
  and g18757 (n10447, n10414, n10445);
  not g18758 (n_10313, n10446);
  not g18759 (n_10314, n10447);
  and g18760 (n10448, n_10313, n_10314);
  not g18761 (n_10315, n10412);
  and g18762 (n10449, n_10315, n10448);
  not g18763 (n_10316, n10448);
  and g18764 (n10450, n10412, n_10316);
  not g18765 (n_10317, n10449);
  not g18766 (n_10318, n10450);
  and g18767 (n10451, n_10317, n_10318);
  not g18768 (n_10319, n10376);
  not g18769 (n_10320, n10451);
  and g18770 (n10452, n_10319, n_10320);
  and g18771 (n10453, n10376, n10451);
  not g18772 (n_10321, n10452);
  not g18773 (n_10322, n10453);
  and g18774 (n10454, n_10321, n_10322);
  not g18775 (n_10323, n10374);
  and g18776 (n10455, n_10323, n10454);
  not g18777 (n_10324, n10454);
  and g18778 (n10456, n10374, n_10324);
  not g18779 (n_10325, n10455);
  not g18780 (n_10326, n10456);
  and g18781 (n10457, n_10325, n_10326);
  not g18782 (n_10327, n10294);
  not g18783 (n_10328, n10457);
  and g18784 (n10458, n_10327, n_10328);
  and g18785 (n10459, n10294, n10457);
  not g18786 (n_10329, n10458);
  not g18787 (n_10330, n10459);
  and g18788 (n10460, n_10329, n_10330);
  not g18789 (n_10331, n10292);
  not g18790 (n_10332, n10460);
  and g18791 (n10461, n_10331, n_10332);
  not g18792 (n_10333, n10291);
  and g18793 (n10462, n_10333, n10461);
  and g18794 (n10463, n_10333, n_10331);
  not g18795 (n_10334, n10463);
  and g18796 (n10464, n10460, n_10334);
  not g18797 (n_10335, n10462);
  not g18798 (n_10336, n10464);
  and g18799 (n10465, n_10335, n_10336);
  not g18800 (n_10337, n10051);
  not g18801 (n_10338, n10465);
  and g18802 (n10466, n_10337, n_10338);
  and g18803 (n10467, n10051, n10465);
  not g18804 (n_10339, n10466);
  not g18805 (n_10340, n10467);
  and g18806 (n10468, n_10339, n_10340);
  and g18807 (n10469, n_9928, n_9926);
  not g18808 (n_10341, n10469);
  and g18809 (n10470, n_9927, n_10341);
  and g18810 (n10471, n_8011, n_8009);
  not g18811 (n_10342, n10471);
  and g18812 (n10472, n_8010, n_10342);
  and g18813 (n10473, n_8004, n_8002);
  not g18814 (n_10343, n10473);
  and g18815 (n10474, n_8003, n_10343);
  and g18816 (n10475, n_7997, n_7995);
  not g18817 (n_10344, n10475);
  and g18818 (n10476, n_7996, n_10344);
  and g18819 (n10477, n_7990, n_7988);
  not g18820 (n_10345, n10477);
  and g18821 (n10478, n_7989, n_10345);
  and g18822 (n10479, n8227, n_7982);
  not g18823 (n_10346, n10479);
  and g18824 (n10480, n_7983, n_10346);
  and g18825 (n10481, n_7757, n_7756);
  not g18826 (n_10347, n10481);
  and g18827 (n10482, n_7755, n_10347);
  and g18828 (n10483, n_7801, n_7800);
  not g18829 (n_10348, n10483);
  and g18830 (n10484, n_7799, n_10348);
  not g18831 (n_10349, n10482);
  and g18832 (n10485, n_10349, n10484);
  not g18833 (n_10350, n10484);
  and g18834 (n10486, n10482, n_10350);
  not g18835 (n_10351, n10485);
  not g18836 (n_10352, n10486);
  and g18837 (n10487, n_10351, n_10352);
  not g18838 (n_10353, n10480);
  not g18839 (n_10354, n10487);
  and g18840 (n10488, n_10353, n_10354);
  not g18844 (n_10355, n10488);
  not g18845 (n_10356, n10491);
  and g18846 (n10492, n_10355, n_10356);
  and g18847 (n10493, n8203, n_7961);
  not g18848 (n_10357, n10493);
  and g18849 (n10494, n_7962, n_10357);
  and g18850 (n10495, n_7665, n_7664);
  not g18851 (n_10358, n10495);
  and g18852 (n10496, n_7663, n_10358);
  and g18853 (n10497, n_7709, n_7708);
  not g18854 (n_10359, n10497);
  and g18855 (n10498, n_7707, n_10359);
  not g18856 (n_10360, n10496);
  and g18857 (n10499, n_10360, n10498);
  not g18858 (n_10361, n10498);
  and g18859 (n10500, n10496, n_10361);
  not g18860 (n_10362, n10499);
  not g18861 (n_10363, n10500);
  and g18862 (n10501, n_10362, n_10363);
  not g18863 (n_10364, n10494);
  not g18864 (n_10365, n10501);
  and g18865 (n10502, n_10364, n_10365);
  not g18869 (n_10366, n10502);
  not g18870 (n_10367, n10505);
  and g18871 (n10506, n_10366, n_10367);
  not g18872 (n_10368, n10492);
  and g18873 (n10507, n_10368, n10506);
  not g18874 (n_10369, n10506);
  and g18875 (n10508, n10492, n_10369);
  not g18876 (n_10370, n10507);
  not g18877 (n_10371, n10508);
  and g18878 (n10509, n_10370, n_10371);
  not g18879 (n_10372, n10478);
  not g18880 (n_10373, n10509);
  and g18881 (n10510, n_10372, n_10373);
  and g18882 (n10511, n10478, n10509);
  not g18883 (n_10374, n10510);
  not g18884 (n_10375, n10511);
  and g18885 (n10512, n_10374, n_10375);
  and g18886 (n10513, n_7946, n_7944);
  not g18887 (n_10376, n10513);
  and g18888 (n10514, n_7945, n_10376);
  and g18889 (n10515, n8148, n_7924);
  not g18890 (n_10377, n10515);
  and g18891 (n10516, n_7925, n_10377);
  and g18892 (n10517, n_7569, n_7568);
  not g18893 (n_10378, n10517);
  and g18894 (n10518, n_7567, n_10378);
  and g18895 (n10519, n_7613, n_7612);
  not g18896 (n_10379, n10519);
  and g18897 (n10520, n_7611, n_10379);
  not g18898 (n_10380, n10518);
  and g18899 (n10521, n_10380, n10520);
  not g18900 (n_10381, n10520);
  and g18901 (n10522, n10518, n_10381);
  not g18902 (n_10382, n10521);
  not g18903 (n_10383, n10522);
  and g18904 (n10523, n_10382, n_10383);
  not g18905 (n_10384, n10516);
  not g18906 (n_10385, n10523);
  and g18907 (n10524, n_10384, n_10385);
  not g18911 (n_10386, n10524);
  not g18912 (n_10387, n10527);
  and g18913 (n10528, n_10386, n_10387);
  and g18914 (n10529, n8167, n_7933);
  not g18915 (n_10388, n10529);
  and g18916 (n10530, n_7934, n_10388);
  and g18917 (n10531, n_7477, n_7476);
  not g18918 (n_10389, n10531);
  and g18919 (n10532, n_7475, n_10389);
  and g18920 (n10533, n_7521, n_7520);
  not g18921 (n_10390, n10533);
  and g18922 (n10534, n_7519, n_10390);
  not g18923 (n_10391, n10532);
  and g18924 (n10535, n_10391, n10534);
  not g18925 (n_10392, n10534);
  and g18926 (n10536, n10532, n_10392);
  not g18927 (n_10393, n10535);
  not g18928 (n_10394, n10536);
  and g18929 (n10537, n_10393, n_10394);
  not g18930 (n_10395, n10530);
  not g18931 (n_10396, n10537);
  and g18932 (n10538, n_10395, n_10396);
  not g18936 (n_10397, n10538);
  not g18937 (n_10398, n10541);
  and g18938 (n10542, n_10397, n_10398);
  not g18939 (n_10399, n10528);
  and g18940 (n10543, n_10399, n10542);
  not g18941 (n_10400, n10542);
  and g18942 (n10544, n10528, n_10400);
  not g18943 (n_10401, n10543);
  not g18944 (n_10402, n10544);
  and g18945 (n10545, n_10401, n_10402);
  not g18946 (n_10403, n10514);
  not g18947 (n_10404, n10545);
  and g18948 (n10546, n_10403, n_10404);
  and g18949 (n10547, n10514, n10545);
  not g18950 (n_10405, n10546);
  not g18951 (n_10406, n10547);
  and g18952 (n10548, n_10405, n_10406);
  not g18953 (n_10407, n10512);
  and g18954 (n10549, n_10407, n10548);
  not g18955 (n_10408, n10548);
  and g18956 (n10550, n10512, n_10408);
  not g18957 (n_10409, n10549);
  not g18958 (n_10410, n10550);
  and g18959 (n10551, n_10409, n_10410);
  not g18960 (n_10411, n10476);
  not g18961 (n_10412, n10551);
  and g18962 (n10552, n_10411, n_10412);
  and g18963 (n10553, n10476, n10551);
  not g18964 (n_10413, n10552);
  not g18965 (n_10414, n10553);
  and g18966 (n10554, n_10413, n_10414);
  and g18967 (n10555, n_7905, n_7903);
  not g18968 (n_10415, n10555);
  and g18969 (n10556, n_7904, n_10415);
  and g18970 (n10557, n_7860, n_7858);
  not g18971 (n_10416, n10557);
  and g18972 (n10558, n_7859, n_10416);
  and g18973 (n10559, n8055, n_7852);
  not g18974 (n_10417, n10559);
  and g18975 (n10560, n_7853, n_10417);
  and g18976 (n10561, n_7377, n_7376);
  not g18977 (n_10418, n10561);
  and g18978 (n10562, n_7375, n_10418);
  and g18979 (n10563, n_7421, n_7420);
  not g18980 (n_10419, n10563);
  and g18981 (n10564, n_7419, n_10419);
  not g18982 (n_10420, n10562);
  and g18983 (n10565, n_10420, n10564);
  not g18984 (n_10421, n10564);
  and g18985 (n10566, n10562, n_10421);
  not g18986 (n_10422, n10565);
  not g18987 (n_10423, n10566);
  and g18988 (n10567, n_10422, n_10423);
  not g18989 (n_10424, n10560);
  not g18990 (n_10425, n10567);
  and g18991 (n10568, n_10424, n_10425);
  not g18995 (n_10426, n10568);
  not g18996 (n_10427, n10571);
  and g18997 (n10572, n_10426, n_10427);
  and g18998 (n10573, n8031, n_7831);
  not g18999 (n_10428, n10573);
  and g19000 (n10574, n_7832, n_10428);
  and g19001 (n10575, n_7285, n_7284);
  not g19002 (n_10429, n10575);
  and g19003 (n10576, n_7283, n_10429);
  and g19004 (n10577, n_7329, n_7328);
  not g19005 (n_10430, n10577);
  and g19006 (n10578, n_7327, n_10430);
  not g19007 (n_10431, n10576);
  and g19008 (n10579, n_10431, n10578);
  not g19009 (n_10432, n10578);
  and g19010 (n10580, n10576, n_10432);
  not g19011 (n_10433, n10579);
  not g19012 (n_10434, n10580);
  and g19013 (n10581, n_10433, n_10434);
  not g19014 (n_10435, n10574);
  not g19015 (n_10436, n10581);
  and g19016 (n10582, n_10435, n_10436);
  not g19020 (n_10437, n10582);
  not g19021 (n_10438, n10585);
  and g19022 (n10586, n_10437, n_10438);
  not g19023 (n_10439, n10572);
  and g19024 (n10587, n_10439, n10586);
  not g19025 (n_10440, n10586);
  and g19026 (n10588, n10572, n_10440);
  not g19027 (n_10441, n10587);
  not g19028 (n_10442, n10588);
  and g19029 (n10589, n_10441, n_10442);
  not g19030 (n_10443, n10558);
  not g19031 (n_10444, n10589);
  and g19032 (n10590, n_10443, n_10444);
  and g19033 (n10591, n10558, n10589);
  not g19034 (n_10445, n10590);
  not g19035 (n_10446, n10591);
  and g19036 (n10592, n_10445, n_10446);
  and g19037 (n10593, n_7894, n_7892);
  not g19038 (n_10447, n10593);
  and g19039 (n10594, n_7893, n_10447);
  and g19040 (n10595, n8081, n_7872);
  not g19041 (n_10448, n10595);
  and g19042 (n10596, n_7873, n_10448);
  and g19043 (n10597, n_7189, n_7188);
  not g19044 (n_10449, n10597);
  and g19045 (n10598, n_7187, n_10449);
  and g19046 (n10599, n_7233, n_7232);
  not g19047 (n_10450, n10599);
  and g19048 (n10600, n_7231, n_10450);
  not g19049 (n_10451, n10598);
  and g19050 (n10601, n_10451, n10600);
  not g19051 (n_10452, n10600);
  and g19052 (n10602, n10598, n_10452);
  not g19053 (n_10453, n10601);
  not g19054 (n_10454, n10602);
  and g19055 (n10603, n_10453, n_10454);
  not g19056 (n_10455, n10596);
  not g19057 (n_10456, n10603);
  and g19058 (n10604, n_10455, n_10456);
  not g19062 (n_10457, n10604);
  not g19063 (n_10458, n10607);
  and g19064 (n10608, n_10457, n_10458);
  and g19065 (n10609, n8100, n_7881);
  not g19066 (n_10459, n10609);
  and g19067 (n10610, n_7882, n_10459);
  and g19068 (n10611, n_7097, n_7096);
  not g19069 (n_10460, n10611);
  and g19070 (n10612, n_7095, n_10460);
  and g19071 (n10613, n_7141, n_7140);
  not g19072 (n_10461, n10613);
  and g19073 (n10614, n_7139, n_10461);
  not g19074 (n_10462, n10612);
  and g19075 (n10615, n_10462, n10614);
  not g19076 (n_10463, n10614);
  and g19077 (n10616, n10612, n_10463);
  not g19078 (n_10464, n10615);
  not g19079 (n_10465, n10616);
  and g19080 (n10617, n_10464, n_10465);
  not g19081 (n_10466, n10610);
  not g19082 (n_10467, n10617);
  and g19083 (n10618, n_10466, n_10467);
  not g19087 (n_10468, n10618);
  not g19088 (n_10469, n10621);
  and g19089 (n10622, n_10468, n_10469);
  not g19090 (n_10470, n10608);
  and g19091 (n10623, n_10470, n10622);
  not g19092 (n_10471, n10622);
  and g19093 (n10624, n10608, n_10471);
  not g19094 (n_10472, n10623);
  not g19095 (n_10473, n10624);
  and g19096 (n10625, n_10472, n_10473);
  not g19097 (n_10474, n10594);
  not g19098 (n_10475, n10625);
  and g19099 (n10626, n_10474, n_10475);
  and g19100 (n10627, n10594, n10625);
  not g19101 (n_10476, n10626);
  not g19102 (n_10477, n10627);
  and g19103 (n10628, n_10476, n_10477);
  not g19104 (n_10478, n10592);
  and g19105 (n10629, n_10478, n10628);
  not g19106 (n_10479, n10628);
  and g19107 (n10630, n10592, n_10479);
  not g19108 (n_10480, n10629);
  not g19109 (n_10481, n10630);
  and g19110 (n10631, n_10480, n_10481);
  not g19111 (n_10482, n10556);
  not g19112 (n_10483, n10631);
  and g19113 (n10632, n_10482, n_10483);
  and g19114 (n10633, n10556, n10631);
  not g19115 (n_10484, n10632);
  not g19116 (n_10485, n10633);
  and g19117 (n10634, n_10484, n_10485);
  not g19118 (n_10486, n10554);
  and g19119 (n10635, n_10486, n10634);
  not g19120 (n_10487, n10634);
  and g19121 (n10636, n10554, n_10487);
  not g19122 (n_10488, n10635);
  not g19123 (n_10489, n10636);
  and g19124 (n10637, n_10488, n_10489);
  not g19125 (n_10490, n10474);
  not g19126 (n_10491, n10637);
  and g19127 (n10638, n_10490, n_10491);
  and g19128 (n10639, n10474, n10637);
  not g19129 (n_10492, n10638);
  not g19130 (n_10493, n10639);
  and g19131 (n10640, n_10492, n_10493);
  and g19132 (n10641, n_7048, n_7046);
  not g19133 (n_10494, n10641);
  and g19134 (n10642, n_7047, n_10494);
  and g19135 (n10643, n_6571, n_6569);
  not g19136 (n_10495, n10643);
  and g19137 (n10644, n_6570, n_10495);
  and g19138 (n10645, n_6564, n_6562);
  not g19139 (n_10496, n10645);
  and g19140 (n10646, n_6563, n_10496);
  and g19141 (n10647, n6933, n_6556);
  not g19142 (n_10497, n10647);
  and g19143 (n10648, n_6557, n_10497);
  and g19144 (n10649, n_6469, n_6468);
  not g19145 (n_10498, n10649);
  and g19146 (n10650, n_6467, n_10498);
  and g19147 (n10651, n_6513, n_6512);
  not g19148 (n_10499, n10651);
  and g19149 (n10652, n_6511, n_10499);
  not g19150 (n_10500, n10650);
  and g19151 (n10653, n_10500, n10652);
  not g19152 (n_10501, n10652);
  and g19153 (n10654, n10650, n_10501);
  not g19154 (n_10502, n10653);
  not g19155 (n_10503, n10654);
  and g19156 (n10655, n_10502, n_10503);
  not g19157 (n_10504, n10648);
  not g19158 (n_10505, n10655);
  and g19159 (n10656, n_10504, n_10505);
  not g19163 (n_10506, n10656);
  not g19164 (n_10507, n10659);
  and g19165 (n10660, n_10506, n_10507);
  and g19166 (n10661, n6909, n_6535);
  not g19167 (n_10508, n10661);
  and g19168 (n10662, n_6536, n_10508);
  and g19169 (n10663, n_6377, n_6376);
  not g19170 (n_10509, n10663);
  and g19171 (n10664, n_6375, n_10509);
  and g19172 (n10665, n_6421, n_6420);
  not g19173 (n_10510, n10665);
  and g19174 (n10666, n_6419, n_10510);
  not g19175 (n_10511, n10664);
  and g19176 (n10667, n_10511, n10666);
  not g19177 (n_10512, n10666);
  and g19178 (n10668, n10664, n_10512);
  not g19179 (n_10513, n10667);
  not g19180 (n_10514, n10668);
  and g19181 (n10669, n_10513, n_10514);
  not g19182 (n_10515, n10662);
  not g19183 (n_10516, n10669);
  and g19184 (n10670, n_10515, n_10516);
  not g19188 (n_10517, n10670);
  not g19189 (n_10518, n10673);
  and g19190 (n10674, n_10517, n_10518);
  not g19191 (n_10519, n10660);
  and g19192 (n10675, n_10519, n10674);
  not g19193 (n_10520, n10674);
  and g19194 (n10676, n10660, n_10520);
  not g19195 (n_10521, n10675);
  not g19196 (n_10522, n10676);
  and g19197 (n10677, n_10521, n_10522);
  not g19198 (n_10523, n10646);
  not g19199 (n_10524, n10677);
  and g19200 (n10678, n_10523, n_10524);
  and g19201 (n10679, n10646, n10677);
  not g19202 (n_10525, n10678);
  not g19203 (n_10526, n10679);
  and g19204 (n10680, n_10525, n_10526);
  and g19205 (n10681, n_6328, n_6326);
  not g19206 (n_10527, n10681);
  and g19207 (n10682, n_6327, n_10527);
  and g19208 (n10683, n6582, n_6208);
  not g19209 (n_10528, n10683);
  and g19210 (n10684, n_6209, n_10528);
  and g19211 (n10685, n_6195, n_6198);
  not g19212 (n_10529, n10685);
  and g19213 (n10686, n_6194, n_10529);
  and g19214 (n10687, n_6154, n_6152);
  not g19215 (n_10530, n10687);
  and g19216 (n10688, n_6153, n_10530);
  not g19217 (n_10531, n10686);
  and g19218 (n10689, n_10531, n10688);
  not g19219 (n_10532, n10688);
  and g19220 (n10690, n10686, n_10532);
  not g19221 (n_10533, n10689);
  not g19222 (n_10534, n10690);
  and g19223 (n10691, n_10533, n_10534);
  not g19224 (n_10535, n10684);
  not g19225 (n_10536, n10691);
  and g19226 (n10692, n_10535, n_10536);
  not g19230 (n_10537, n10692);
  not g19231 (n_10538, n10695);
  and g19232 (n10696, n_10537, n_10538);
  and g19233 (n10697, n6671, n_6305);
  not g19234 (n_10539, n10697);
  and g19235 (n10698, n_6306, n_10539);
  and g19236 (n10699, n_6296, n_6299);
  not g19237 (n_10540, n10699);
  and g19238 (n10700, n_6295, n_10540);
  and g19239 (n10701, n_6255, n_6253);
  not g19240 (n_10541, n10701);
  and g19241 (n10702, n_6254, n_10541);
  not g19242 (n_10542, n10700);
  and g19243 (n10703, n_10542, n10702);
  not g19244 (n_10543, n10702);
  and g19245 (n10704, n10700, n_10543);
  not g19246 (n_10544, n10703);
  not g19247 (n_10545, n10704);
  and g19248 (n10705, n_10544, n_10545);
  not g19249 (n_10546, n10698);
  not g19250 (n_10547, n10705);
  and g19251 (n10706, n_10546, n_10547);
  not g19255 (n_10548, n10706);
  not g19256 (n_10549, n10709);
  and g19257 (n10710, n_10548, n_10549);
  not g19258 (n_10550, n10696);
  and g19259 (n10711, n_10550, n10710);
  not g19260 (n_10551, n10710);
  and g19261 (n10712, n10696, n_10551);
  not g19262 (n_10552, n10711);
  not g19263 (n_10553, n10712);
  and g19264 (n10713, n_10552, n_10553);
  not g19265 (n_10554, n10682);
  not g19266 (n_10555, n10713);
  and g19267 (n10714, n_10554, n_10555);
  and g19268 (n10715, n10682, n10713);
  not g19269 (n_10556, n10714);
  not g19270 (n_10557, n10715);
  and g19271 (n10716, n_10556, n_10557);
  not g19272 (n_10558, n10680);
  and g19273 (n10717, n_10558, n10716);
  not g19274 (n_10559, n10716);
  and g19275 (n10718, n10680, n_10559);
  not g19276 (n_10560, n10717);
  not g19277 (n_10561, n10718);
  and g19278 (n10719, n_10560, n_10561);
  not g19279 (n_10562, n10644);
  not g19280 (n_10563, n10719);
  and g19281 (n10720, n_10562, n_10563);
  and g19282 (n10721, n10644, n10719);
  not g19283 (n_10564, n10720);
  not g19284 (n_10565, n10721);
  and g19285 (n10722, n_10564, n_10565);
  and g19286 (n10723, n_7031, n_7029);
  not g19287 (n_10566, n10723);
  and g19288 (n10724, n_7030, n_10566);
  and g19289 (n10725, n_6794, n_6792);
  not g19290 (n_10567, n10725);
  and g19291 (n10726, n_6793, n_10567);
  and g19292 (n10727, n7140, n_6786);
  not g19293 (n_10568, n10727);
  and g19294 (n10728, n_6787, n_10568);
  and g19295 (n10729, n_6720, n_6719);
  not g19296 (n_10569, n10729);
  and g19297 (n10730, n_6718, n_10569);
  and g19298 (n10731, n_6764, n_6763);
  not g19299 (n_10570, n10731);
  and g19300 (n10732, n_6762, n_10570);
  not g19301 (n_10571, n10730);
  and g19302 (n10733, n_10571, n10732);
  not g19303 (n_10572, n10732);
  and g19304 (n10734, n10730, n_10572);
  not g19305 (n_10573, n10733);
  not g19306 (n_10574, n10734);
  and g19307 (n10735, n_10573, n_10574);
  not g19308 (n_10575, n10728);
  not g19309 (n_10576, n10735);
  and g19310 (n10736, n_10575, n_10576);
  not g19314 (n_10577, n10736);
  not g19315 (n_10578, n10739);
  and g19316 (n10740, n_10577, n_10578);
  and g19317 (n10741, n7000, n_6667);
  not g19318 (n_10579, n10741);
  and g19319 (n10742, n_6668, n_10579);
  and g19320 (n10743, n_6658, n_6661);
  not g19321 (n_10580, n10743);
  and g19322 (n10744, n_6657, n_10580);
  and g19323 (n10745, n_6617, n_6615);
  not g19324 (n_10581, n10745);
  and g19325 (n10746, n_6616, n_10581);
  not g19326 (n_10582, n10744);
  and g19327 (n10747, n_10582, n10746);
  not g19328 (n_10583, n10746);
  and g19329 (n10748, n10744, n_10583);
  not g19330 (n_10584, n10747);
  not g19331 (n_10585, n10748);
  and g19332 (n10749, n_10584, n_10585);
  not g19333 (n_10586, n10742);
  not g19334 (n_10587, n10749);
  and g19335 (n10750, n_10586, n_10587);
  not g19339 (n_10588, n10750);
  not g19340 (n_10589, n10753);
  and g19341 (n10754, n_10588, n_10589);
  not g19342 (n_10590, n10740);
  and g19343 (n10755, n_10590, n10754);
  not g19344 (n_10591, n10754);
  and g19345 (n10756, n10740, n_10591);
  not g19346 (n_10592, n10755);
  not g19347 (n_10593, n10756);
  and g19348 (n10757, n_10592, n_10593);
  not g19349 (n_10594, n10726);
  not g19350 (n_10595, n10757);
  and g19351 (n10758, n_10594, n_10595);
  and g19352 (n10759, n10726, n10757);
  not g19353 (n_10596, n10758);
  not g19354 (n_10597, n10759);
  and g19355 (n10760, n_10596, n_10597);
  and g19356 (n10761, n_7014, n_7012);
  not g19357 (n_10598, n10761);
  and g19358 (n10762, n_7013, n_10598);
  and g19359 (n10763, n7200, n_6894);
  not g19360 (n_10599, n10763);
  and g19361 (n10764, n_6895, n_10599);
  and g19362 (n10765, n_6881, n_6884);
  not g19363 (n_10600, n10765);
  and g19364 (n10766, n_6880, n_10600);
  and g19365 (n10767, n_6840, n_6838);
  not g19366 (n_10601, n10767);
  and g19367 (n10768, n_6839, n_10601);
  not g19368 (n_10602, n10766);
  and g19369 (n10769, n_10602, n10768);
  not g19370 (n_10603, n10768);
  and g19371 (n10770, n10766, n_10603);
  not g19372 (n_10604, n10769);
  not g19373 (n_10605, n10770);
  and g19374 (n10771, n_10604, n_10605);
  not g19375 (n_10606, n10764);
  not g19376 (n_10607, n10771);
  and g19377 (n10772, n_10606, n_10607);
  not g19381 (n_10608, n10772);
  not g19382 (n_10609, n10775);
  and g19383 (n10776, n_10608, n_10609);
  and g19384 (n10777, n7289, n_6991);
  not g19385 (n_10610, n10777);
  and g19386 (n10778, n_6992, n_10610);
  and g19387 (n10779, n_6982, n_6985);
  not g19388 (n_10611, n10779);
  and g19389 (n10780, n_6981, n_10611);
  and g19390 (n10781, n_6941, n_6939);
  not g19391 (n_10612, n10781);
  and g19392 (n10782, n_6940, n_10612);
  not g19393 (n_10613, n10780);
  and g19394 (n10783, n_10613, n10782);
  not g19395 (n_10614, n10782);
  and g19396 (n10784, n10780, n_10614);
  not g19397 (n_10615, n10783);
  not g19398 (n_10616, n10784);
  and g19399 (n10785, n_10615, n_10616);
  not g19400 (n_10617, n10778);
  not g19401 (n_10618, n10785);
  and g19402 (n10786, n_10617, n_10618);
  not g19406 (n_10619, n10786);
  not g19407 (n_10620, n10789);
  and g19408 (n10790, n_10619, n_10620);
  not g19409 (n_10621, n10776);
  and g19410 (n10791, n_10621, n10790);
  not g19411 (n_10622, n10790);
  and g19412 (n10792, n10776, n_10622);
  not g19413 (n_10623, n10791);
  not g19414 (n_10624, n10792);
  and g19415 (n10793, n_10623, n_10624);
  not g19416 (n_10625, n10762);
  not g19417 (n_10626, n10793);
  and g19418 (n10794, n_10625, n_10626);
  and g19419 (n10795, n10762, n10793);
  not g19420 (n_10627, n10794);
  not g19421 (n_10628, n10795);
  and g19422 (n10796, n_10627, n_10628);
  not g19423 (n_10629, n10760);
  and g19424 (n10797, n_10629, n10796);
  not g19425 (n_10630, n10796);
  and g19426 (n10798, n10760, n_10630);
  not g19427 (n_10631, n10797);
  not g19428 (n_10632, n10798);
  and g19429 (n10799, n_10631, n_10632);
  not g19430 (n_10633, n10724);
  not g19431 (n_10634, n10799);
  and g19432 (n10800, n_10633, n_10634);
  and g19433 (n10801, n10724, n10799);
  not g19434 (n_10635, n10800);
  not g19435 (n_10636, n10801);
  and g19436 (n10802, n_10635, n_10636);
  not g19437 (n_10637, n10722);
  and g19438 (n10803, n_10637, n10802);
  not g19439 (n_10638, n10802);
  and g19440 (n10804, n10722, n_10638);
  not g19441 (n_10639, n10803);
  not g19442 (n_10640, n10804);
  and g19443 (n10805, n_10639, n_10640);
  not g19444 (n_10641, n10642);
  not g19445 (n_10642, n10805);
  and g19446 (n10806, n_10641, n_10642);
  and g19447 (n10807, n10642, n10805);
  not g19448 (n_10643, n10806);
  not g19449 (n_10644, n10807);
  and g19450 (n10808, n_10643, n_10644);
  not g19451 (n_10645, n10640);
  and g19452 (n10809, n_10645, n10808);
  not g19453 (n_10646, n10808);
  and g19454 (n10810, n10640, n_10646);
  not g19455 (n_10647, n10809);
  not g19456 (n_10648, n10810);
  and g19457 (n10811, n_10647, n_10648);
  not g19458 (n_10649, n10472);
  not g19459 (n_10650, n10811);
  and g19460 (n10812, n_10649, n_10650);
  and g19461 (n10813, n10472, n10811);
  not g19462 (n_10651, n10812);
  not g19463 (n_10652, n10813);
  and g19464 (n10814, n_10651, n_10652);
  and g19465 (n10815, n_9911, n_9909);
  not g19466 (n_10653, n10815);
  and g19467 (n10816, n_9910, n_10653);
  and g19468 (n10817, n_8954, n_8952);
  not g19469 (n_10654, n10817);
  and g19470 (n10818, n_8953, n_10654);
  and g19471 (n10819, n_8947, n_8945);
  not g19472 (n_10655, n10819);
  and g19473 (n10820, n_8946, n_10655);
  and g19474 (n10821, n_8940, n_8938);
  not g19475 (n_10656, n10821);
  and g19476 (n10822, n_8939, n_10656);
  and g19477 (n10823, n9088, n_8932);
  not g19478 (n_10657, n10823);
  and g19479 (n10824, n_8933, n_10657);
  and g19480 (n10825, n_8800, n_8799);
  not g19481 (n_10658, n10825);
  and g19482 (n10826, n_8798, n_10658);
  and g19483 (n10827, n_8844, n_8843);
  not g19484 (n_10659, n10827);
  and g19485 (n10828, n_8842, n_10659);
  not g19486 (n_10660, n10826);
  and g19487 (n10829, n_10660, n10828);
  not g19488 (n_10661, n10828);
  and g19489 (n10830, n10826, n_10661);
  not g19490 (n_10662, n10829);
  not g19491 (n_10663, n10830);
  and g19492 (n10831, n_10662, n_10663);
  not g19493 (n_10664, n10824);
  not g19494 (n_10665, n10831);
  and g19495 (n10832, n_10664, n_10665);
  not g19499 (n_10666, n10832);
  not g19500 (n_10667, n10835);
  and g19501 (n10836, n_10666, n_10667);
  and g19502 (n10837, n9064, n_8911);
  not g19503 (n_10668, n10837);
  and g19504 (n10838, n_8912, n_10668);
  and g19505 (n10839, n_8708, n_8707);
  not g19506 (n_10669, n10839);
  and g19507 (n10840, n_8706, n_10669);
  and g19508 (n10841, n_8752, n_8751);
  not g19509 (n_10670, n10841);
  and g19510 (n10842, n_8750, n_10670);
  not g19511 (n_10671, n10840);
  and g19512 (n10843, n_10671, n10842);
  not g19513 (n_10672, n10842);
  and g19514 (n10844, n10840, n_10672);
  not g19515 (n_10673, n10843);
  not g19516 (n_10674, n10844);
  and g19517 (n10845, n_10673, n_10674);
  not g19518 (n_10675, n10838);
  not g19519 (n_10676, n10845);
  and g19520 (n10846, n_10675, n_10676);
  not g19524 (n_10677, n10846);
  not g19525 (n_10678, n10849);
  and g19526 (n10850, n_10677, n_10678);
  not g19527 (n_10679, n10836);
  and g19528 (n10851, n_10679, n10850);
  not g19529 (n_10680, n10850);
  and g19530 (n10852, n10836, n_10680);
  not g19531 (n_10681, n10851);
  not g19532 (n_10682, n10852);
  and g19533 (n10853, n_10681, n_10682);
  not g19534 (n_10683, n10822);
  not g19535 (n_10684, n10853);
  and g19536 (n10854, n_10683, n_10684);
  and g19537 (n10855, n10822, n10853);
  not g19538 (n_10685, n10854);
  not g19539 (n_10686, n10855);
  and g19540 (n10856, n_10685, n_10686);
  and g19541 (n10857, n_8896, n_8894);
  not g19542 (n_10687, n10857);
  and g19543 (n10858, n_8895, n_10687);
  and g19544 (n10859, n9009, n_8874);
  not g19545 (n_10688, n10859);
  and g19546 (n10860, n_8875, n_10688);
  and g19547 (n10861, n_8612, n_8611);
  not g19548 (n_10689, n10861);
  and g19549 (n10862, n_8610, n_10689);
  and g19550 (n10863, n_8656, n_8655);
  not g19551 (n_10690, n10863);
  and g19552 (n10864, n_8654, n_10690);
  not g19553 (n_10691, n10862);
  and g19554 (n10865, n_10691, n10864);
  not g19555 (n_10692, n10864);
  and g19556 (n10866, n10862, n_10692);
  not g19557 (n_10693, n10865);
  not g19558 (n_10694, n10866);
  and g19559 (n10867, n_10693, n_10694);
  not g19560 (n_10695, n10860);
  not g19561 (n_10696, n10867);
  and g19562 (n10868, n_10695, n_10696);
  not g19566 (n_10697, n10868);
  not g19567 (n_10698, n10871);
  and g19568 (n10872, n_10697, n_10698);
  and g19569 (n10873, n9028, n_8883);
  not g19570 (n_10699, n10873);
  and g19571 (n10874, n_8884, n_10699);
  and g19572 (n10875, n_8520, n_8519);
  not g19573 (n_10700, n10875);
  and g19574 (n10876, n_8518, n_10700);
  and g19575 (n10877, n_8564, n_8563);
  not g19576 (n_10701, n10877);
  and g19577 (n10878, n_8562, n_10701);
  not g19578 (n_10702, n10876);
  and g19579 (n10879, n_10702, n10878);
  not g19580 (n_10703, n10878);
  and g19581 (n10880, n10876, n_10703);
  not g19582 (n_10704, n10879);
  not g19583 (n_10705, n10880);
  and g19584 (n10881, n_10704, n_10705);
  not g19585 (n_10706, n10874);
  not g19586 (n_10707, n10881);
  and g19587 (n10882, n_10706, n_10707);
  not g19591 (n_10708, n10882);
  not g19592 (n_10709, n10885);
  and g19593 (n10886, n_10708, n_10709);
  not g19594 (n_10710, n10872);
  and g19595 (n10887, n_10710, n10886);
  not g19596 (n_10711, n10886);
  and g19597 (n10888, n10872, n_10711);
  not g19598 (n_10712, n10887);
  not g19599 (n_10713, n10888);
  and g19600 (n10889, n_10712, n_10713);
  not g19601 (n_10714, n10858);
  not g19602 (n_10715, n10889);
  and g19603 (n10890, n_10714, n_10715);
  and g19604 (n10891, n10858, n10889);
  not g19605 (n_10716, n10890);
  not g19606 (n_10717, n10891);
  and g19607 (n10892, n_10716, n_10717);
  not g19608 (n_10718, n10856);
  and g19609 (n10893, n_10718, n10892);
  not g19610 (n_10719, n10892);
  and g19611 (n10894, n10856, n_10719);
  not g19612 (n_10720, n10893);
  not g19613 (n_10721, n10894);
  and g19614 (n10895, n_10720, n_10721);
  not g19615 (n_10722, n10820);
  not g19616 (n_10723, n10895);
  and g19617 (n10896, n_10722, n_10723);
  and g19618 (n10897, n10820, n10895);
  not g19619 (n_10724, n10896);
  not g19620 (n_10725, n10897);
  and g19621 (n10898, n_10724, n_10725);
  and g19622 (n10899, n_8471, n_8469);
  not g19623 (n_10726, n10899);
  and g19624 (n10900, n_8470, n_10726);
  and g19625 (n10901, n_8234, n_8232);
  not g19626 (n_10727, n10901);
  and g19627 (n10902, n_8233, n_10727);
  and g19628 (n10903, n8448, n_8226);
  not g19629 (n_10728, n10903);
  and g19630 (n10904, n_8227, n_10728);
  and g19631 (n10905, n_8160, n_8159);
  not g19632 (n_10729, n10905);
  and g19633 (n10906, n_8158, n_10729);
  and g19634 (n10907, n_8204, n_8203);
  not g19635 (n_10730, n10907);
  and g19636 (n10908, n_8202, n_10730);
  not g19637 (n_10731, n10906);
  and g19638 (n10909, n_10731, n10908);
  not g19639 (n_10732, n10908);
  and g19640 (n10910, n10906, n_10732);
  not g19641 (n_10733, n10909);
  not g19642 (n_10734, n10910);
  and g19643 (n10911, n_10733, n_10734);
  not g19644 (n_10735, n10904);
  not g19645 (n_10736, n10911);
  and g19646 (n10912, n_10735, n_10736);
  not g19650 (n_10737, n10912);
  not g19651 (n_10738, n10915);
  and g19652 (n10916, n_10737, n_10738);
  and g19653 (n10917, n8308, n_8107);
  not g19654 (n_10739, n10917);
  and g19655 (n10918, n_8108, n_10739);
  and g19656 (n10919, n_8098, n_8101);
  not g19657 (n_10740, n10919);
  and g19658 (n10920, n_8097, n_10740);
  and g19659 (n10921, n_8057, n_8055);
  not g19660 (n_10741, n10921);
  and g19661 (n10922, n_8056, n_10741);
  not g19662 (n_10742, n10920);
  and g19663 (n10923, n_10742, n10922);
  not g19664 (n_10743, n10922);
  and g19665 (n10924, n10920, n_10743);
  not g19666 (n_10744, n10923);
  not g19667 (n_10745, n10924);
  and g19668 (n10925, n_10744, n_10745);
  not g19669 (n_10746, n10918);
  not g19670 (n_10747, n10925);
  and g19671 (n10926, n_10746, n_10747);
  not g19675 (n_10748, n10926);
  not g19676 (n_10749, n10929);
  and g19677 (n10930, n_10748, n_10749);
  not g19678 (n_10750, n10916);
  and g19679 (n10931, n_10750, n10930);
  not g19680 (n_10751, n10930);
  and g19681 (n10932, n10916, n_10751);
  not g19682 (n_10752, n10931);
  not g19683 (n_10753, n10932);
  and g19684 (n10933, n_10752, n_10753);
  not g19685 (n_10754, n10902);
  not g19686 (n_10755, n10933);
  and g19687 (n10934, n_10754, n_10755);
  and g19688 (n10935, n10902, n10933);
  not g19689 (n_10756, n10934);
  not g19690 (n_10757, n10935);
  and g19691 (n10936, n_10756, n_10757);
  and g19692 (n10937, n_8454, n_8452);
  not g19693 (n_10758, n10937);
  and g19694 (n10938, n_8453, n_10758);
  and g19695 (n10939, n8508, n_8334);
  not g19696 (n_10759, n10939);
  and g19697 (n10940, n_8335, n_10759);
  and g19698 (n10941, n_8321, n_8324);
  not g19699 (n_10760, n10941);
  and g19700 (n10942, n_8320, n_10760);
  and g19701 (n10943, n_8280, n_8278);
  not g19702 (n_10761, n10943);
  and g19703 (n10944, n_8279, n_10761);
  not g19704 (n_10762, n10942);
  and g19705 (n10945, n_10762, n10944);
  not g19706 (n_10763, n10944);
  and g19707 (n10946, n10942, n_10763);
  not g19708 (n_10764, n10945);
  not g19709 (n_10765, n10946);
  and g19710 (n10947, n_10764, n_10765);
  not g19711 (n_10766, n10940);
  not g19712 (n_10767, n10947);
  and g19713 (n10948, n_10766, n_10767);
  not g19717 (n_10768, n10948);
  not g19718 (n_10769, n10951);
  and g19719 (n10952, n_10768, n_10769);
  and g19720 (n10953, n8597, n_8431);
  not g19721 (n_10770, n10953);
  and g19722 (n10954, n_8432, n_10770);
  and g19723 (n10955, n_8422, n_8425);
  not g19724 (n_10771, n10955);
  and g19725 (n10956, n_8421, n_10771);
  and g19726 (n10957, n_8381, n_8379);
  not g19727 (n_10772, n10957);
  and g19728 (n10958, n_8380, n_10772);
  not g19729 (n_10773, n10956);
  and g19730 (n10959, n_10773, n10958);
  not g19731 (n_10774, n10958);
  and g19732 (n10960, n10956, n_10774);
  not g19733 (n_10775, n10959);
  not g19734 (n_10776, n10960);
  and g19735 (n10961, n_10775, n_10776);
  not g19736 (n_10777, n10954);
  not g19737 (n_10778, n10961);
  and g19738 (n10962, n_10777, n_10778);
  not g19742 (n_10779, n10962);
  not g19743 (n_10780, n10965);
  and g19744 (n10966, n_10779, n_10780);
  not g19745 (n_10781, n10952);
  and g19746 (n10967, n_10781, n10966);
  not g19747 (n_10782, n10966);
  and g19748 (n10968, n10952, n_10782);
  not g19749 (n_10783, n10967);
  not g19750 (n_10784, n10968);
  and g19751 (n10969, n_10783, n_10784);
  not g19752 (n_10785, n10938);
  not g19753 (n_10786, n10969);
  and g19754 (n10970, n_10785, n_10786);
  and g19755 (n10971, n10938, n10969);
  not g19756 (n_10787, n10970);
  not g19757 (n_10788, n10971);
  and g19758 (n10972, n_10787, n_10788);
  not g19759 (n_10789, n10936);
  and g19760 (n10973, n_10789, n10972);
  not g19761 (n_10790, n10972);
  and g19762 (n10974, n10936, n_10790);
  not g19763 (n_10791, n10973);
  not g19764 (n_10792, n10974);
  and g19765 (n10975, n_10791, n_10792);
  not g19766 (n_10793, n10900);
  not g19767 (n_10794, n10975);
  and g19768 (n10976, n_10793, n_10794);
  and g19769 (n10977, n10900, n10975);
  not g19770 (n_10795, n10976);
  not g19771 (n_10796, n10977);
  and g19772 (n10978, n_10795, n_10796);
  not g19773 (n_10797, n10898);
  and g19774 (n10979, n_10797, n10978);
  not g19775 (n_10798, n10978);
  and g19776 (n10980, n10898, n_10798);
  not g19777 (n_10799, n10979);
  not g19778 (n_10800, n10980);
  and g19779 (n10981, n_10799, n_10800);
  not g19780 (n_10801, n10818);
  not g19781 (n_10802, n10981);
  and g19782 (n10982, n_10801, n_10802);
  and g19783 (n10983, n10818, n10981);
  not g19784 (n_10803, n10982);
  not g19785 (n_10804, n10983);
  and g19786 (n10984, n_10803, n_10804);
  and g19787 (n10985, n_9894, n_9892);
  not g19788 (n_10805, n10985);
  and g19789 (n10986, n_9893, n_10805);
  and g19790 (n10987, n_9417, n_9415);
  not g19791 (n_10806, n10987);
  and g19792 (n10988, n_9416, n_10806);
  and g19793 (n10989, n_9410, n_9408);
  not g19794 (n_10807, n10989);
  and g19795 (n10990, n_9409, n_10807);
  and g19796 (n10991, n9513, n_9402);
  not g19797 (n_10808, n10991);
  and g19798 (n10992, n_9403, n_10808);
  and g19799 (n10993, n_9315, n_9314);
  not g19800 (n_10809, n10993);
  and g19801 (n10994, n_9313, n_10809);
  and g19802 (n10995, n_9359, n_9358);
  not g19803 (n_10810, n10995);
  and g19804 (n10996, n_9357, n_10810);
  not g19805 (n_10811, n10994);
  and g19806 (n10997, n_10811, n10996);
  not g19807 (n_10812, n10996);
  and g19808 (n10998, n10994, n_10812);
  not g19809 (n_10813, n10997);
  not g19810 (n_10814, n10998);
  and g19811 (n10999, n_10813, n_10814);
  not g19812 (n_10815, n10992);
  not g19813 (n_10816, n10999);
  and g19814 (n11000, n_10815, n_10816);
  not g19818 (n_10817, n11000);
  not g19819 (n_10818, n11003);
  and g19820 (n11004, n_10817, n_10818);
  and g19821 (n11005, n9489, n_9381);
  not g19822 (n_10819, n11005);
  and g19823 (n11006, n_9382, n_10819);
  and g19824 (n11007, n_9223, n_9222);
  not g19825 (n_10820, n11007);
  and g19826 (n11008, n_9221, n_10820);
  and g19827 (n11009, n_9267, n_9266);
  not g19828 (n_10821, n11009);
  and g19829 (n11010, n_9265, n_10821);
  not g19830 (n_10822, n11008);
  and g19831 (n11011, n_10822, n11010);
  not g19832 (n_10823, n11010);
  and g19833 (n11012, n11008, n_10823);
  not g19834 (n_10824, n11011);
  not g19835 (n_10825, n11012);
  and g19836 (n11013, n_10824, n_10825);
  not g19837 (n_10826, n11006);
  not g19838 (n_10827, n11013);
  and g19839 (n11014, n_10826, n_10827);
  not g19843 (n_10828, n11014);
  not g19844 (n_10829, n11017);
  and g19845 (n11018, n_10828, n_10829);
  not g19846 (n_10830, n11004);
  and g19847 (n11019, n_10830, n11018);
  not g19848 (n_10831, n11018);
  and g19849 (n11020, n11004, n_10831);
  not g19850 (n_10832, n11019);
  not g19851 (n_10833, n11020);
  and g19852 (n11021, n_10832, n_10833);
  not g19853 (n_10834, n10990);
  not g19854 (n_10835, n11021);
  and g19855 (n11022, n_10834, n_10835);
  and g19856 (n11023, n10990, n11021);
  not g19857 (n_10836, n11022);
  not g19858 (n_10837, n11023);
  and g19859 (n11024, n_10836, n_10837);
  and g19860 (n11025, n_9174, n_9172);
  not g19861 (n_10838, n11025);
  and g19862 (n11026, n_9173, n_10838);
  and g19863 (n11027, n9162, n_9054);
  not g19864 (n_10839, n11027);
  and g19865 (n11028, n_9055, n_10839);
  and g19866 (n11029, n_9041, n_9044);
  not g19867 (n_10840, n11029);
  and g19868 (n11030, n_9040, n_10840);
  and g19869 (n11031, n_9000, n_8998);
  not g19870 (n_10841, n11031);
  and g19871 (n11032, n_8999, n_10841);
  not g19872 (n_10842, n11030);
  and g19873 (n11033, n_10842, n11032);
  not g19874 (n_10843, n11032);
  and g19875 (n11034, n11030, n_10843);
  not g19876 (n_10844, n11033);
  not g19877 (n_10845, n11034);
  and g19878 (n11035, n_10844, n_10845);
  not g19879 (n_10846, n11028);
  not g19880 (n_10847, n11035);
  and g19881 (n11036, n_10846, n_10847);
  not g19885 (n_10848, n11036);
  not g19886 (n_10849, n11039);
  and g19887 (n11040, n_10848, n_10849);
  and g19888 (n11041, n9251, n_9151);
  not g19889 (n_10850, n11041);
  and g19890 (n11042, n_9152, n_10850);
  and g19891 (n11043, n_9142, n_9145);
  not g19892 (n_10851, n11043);
  and g19893 (n11044, n_9141, n_10851);
  and g19894 (n11045, n_9101, n_9099);
  not g19895 (n_10852, n11045);
  and g19896 (n11046, n_9100, n_10852);
  not g19897 (n_10853, n11044);
  and g19898 (n11047, n_10853, n11046);
  not g19899 (n_10854, n11046);
  and g19900 (n11048, n11044, n_10854);
  not g19901 (n_10855, n11047);
  not g19902 (n_10856, n11048);
  and g19903 (n11049, n_10855, n_10856);
  not g19904 (n_10857, n11042);
  not g19905 (n_10858, n11049);
  and g19906 (n11050, n_10857, n_10858);
  not g19910 (n_10859, n11050);
  not g19911 (n_10860, n11053);
  and g19912 (n11054, n_10859, n_10860);
  not g19913 (n_10861, n11040);
  and g19914 (n11055, n_10861, n11054);
  not g19915 (n_10862, n11054);
  and g19916 (n11056, n11040, n_10862);
  not g19917 (n_10863, n11055);
  not g19918 (n_10864, n11056);
  and g19919 (n11057, n_10863, n_10864);
  not g19920 (n_10865, n11026);
  not g19921 (n_10866, n11057);
  and g19922 (n11058, n_10865, n_10866);
  and g19923 (n11059, n11026, n11057);
  not g19924 (n_10867, n11058);
  not g19925 (n_10868, n11059);
  and g19926 (n11060, n_10867, n_10868);
  not g19927 (n_10869, n11024);
  and g19928 (n11061, n_10869, n11060);
  not g19929 (n_10870, n11060);
  and g19930 (n11062, n11024, n_10870);
  not g19931 (n_10871, n11061);
  not g19932 (n_10872, n11062);
  and g19933 (n11063, n_10871, n_10872);
  not g19934 (n_10873, n10988);
  not g19935 (n_10874, n11063);
  and g19936 (n11064, n_10873, n_10874);
  and g19937 (n11065, n10988, n11063);
  not g19938 (n_10875, n11064);
  not g19939 (n_10876, n11065);
  and g19940 (n11066, n_10875, n_10876);
  and g19941 (n11067, n_9877, n_9875);
  not g19942 (n_10877, n11067);
  and g19943 (n11068, n_9876, n_10877);
  and g19944 (n11069, n_9640, n_9638);
  not g19945 (n_10878, n11069);
  and g19946 (n11070, n_9639, n_10878);
  and g19947 (n11071, n9720, n_9632);
  not g19948 (n_10879, n11071);
  and g19949 (n11072, n_9633, n_10879);
  and g19950 (n11073, n_9566, n_9565);
  not g19951 (n_10880, n11073);
  and g19952 (n11074, n_9564, n_10880);
  and g19953 (n11075, n_9610, n_9609);
  not g19954 (n_10881, n11075);
  and g19955 (n11076, n_9608, n_10881);
  not g19956 (n_10882, n11074);
  and g19957 (n11077, n_10882, n11076);
  not g19958 (n_10883, n11076);
  and g19959 (n11078, n11074, n_10883);
  not g19960 (n_10884, n11077);
  not g19961 (n_10885, n11078);
  and g19962 (n11079, n_10884, n_10885);
  not g19963 (n_10886, n11072);
  not g19964 (n_10887, n11079);
  and g19965 (n11080, n_10886, n_10887);
  not g19969 (n_10888, n11080);
  not g19970 (n_10889, n11083);
  and g19971 (n11084, n_10888, n_10889);
  and g19972 (n11085, n9580, n_9513);
  not g19973 (n_10890, n11085);
  and g19974 (n11086, n_9514, n_10890);
  and g19975 (n11087, n_9504, n_9507);
  not g19976 (n_10891, n11087);
  and g19977 (n11088, n_9503, n_10891);
  and g19978 (n11089, n_9463, n_9461);
  not g19979 (n_10892, n11089);
  and g19980 (n11090, n_9462, n_10892);
  not g19981 (n_10893, n11088);
  and g19982 (n11091, n_10893, n11090);
  not g19983 (n_10894, n11090);
  and g19984 (n11092, n11088, n_10894);
  not g19985 (n_10895, n11091);
  not g19986 (n_10896, n11092);
  and g19987 (n11093, n_10895, n_10896);
  not g19988 (n_10897, n11086);
  not g19989 (n_10898, n11093);
  and g19990 (n11094, n_10897, n_10898);
  not g19994 (n_10899, n11094);
  not g19995 (n_10900, n11097);
  and g19996 (n11098, n_10899, n_10900);
  not g19997 (n_10901, n11084);
  and g19998 (n11099, n_10901, n11098);
  not g19999 (n_10902, n11098);
  and g20000 (n11100, n11084, n_10902);
  not g20001 (n_10903, n11099);
  not g20002 (n_10904, n11100);
  and g20003 (n11101, n_10903, n_10904);
  not g20004 (n_10905, n11070);
  not g20005 (n_10906, n11101);
  and g20006 (n11102, n_10905, n_10906);
  and g20007 (n11103, n11070, n11101);
  not g20008 (n_10907, n11102);
  not g20009 (n_10908, n11103);
  and g20010 (n11104, n_10907, n_10908);
  and g20011 (n11105, n_9860, n_9858);
  not g20012 (n_10909, n11105);
  and g20013 (n11106, n_9859, n_10909);
  and g20014 (n11107, n9780, n_9740);
  not g20015 (n_10910, n11107);
  and g20016 (n11108, n_9741, n_10910);
  and g20017 (n11109, n_9727, n_9730);
  not g20018 (n_10911, n11109);
  and g20019 (n11110, n_9726, n_10911);
  and g20020 (n11111, n_9686, n_9684);
  not g20021 (n_10912, n11111);
  and g20022 (n11112, n_9685, n_10912);
  not g20023 (n_10913, n11110);
  and g20024 (n11113, n_10913, n11112);
  not g20025 (n_10914, n11112);
  and g20026 (n11114, n11110, n_10914);
  not g20027 (n_10915, n11113);
  not g20028 (n_10916, n11114);
  and g20029 (n11115, n_10915, n_10916);
  not g20030 (n_10917, n11108);
  not g20031 (n_10918, n11115);
  and g20032 (n11116, n_10917, n_10918);
  not g20036 (n_10919, n11116);
  not g20037 (n_10920, n11119);
  and g20038 (n11120, n_10919, n_10920);
  and g20039 (n11121, n9869, n_9837);
  not g20040 (n_10921, n11121);
  and g20041 (n11122, n_9838, n_10921);
  and g20042 (n11123, n_9828, n_9831);
  not g20043 (n_10922, n11123);
  and g20044 (n11124, n_9827, n_10922);
  and g20045 (n11125, n_9787, n_9785);
  not g20046 (n_10923, n11125);
  and g20047 (n11126, n_9786, n_10923);
  not g20048 (n_10924, n11124);
  and g20049 (n11127, n_10924, n11126);
  not g20050 (n_10925, n11126);
  and g20051 (n11128, n11124, n_10925);
  not g20052 (n_10926, n11127);
  not g20053 (n_10927, n11128);
  and g20054 (n11129, n_10926, n_10927);
  not g20055 (n_10928, n11122);
  not g20056 (n_10929, n11129);
  and g20057 (n11130, n_10928, n_10929);
  not g20061 (n_10930, n11130);
  not g20062 (n_10931, n11133);
  and g20063 (n11134, n_10930, n_10931);
  not g20064 (n_10932, n11120);
  and g20065 (n11135, n_10932, n11134);
  not g20066 (n_10933, n11134);
  and g20067 (n11136, n11120, n_10933);
  not g20068 (n_10934, n11135);
  not g20069 (n_10935, n11136);
  and g20070 (n11137, n_10934, n_10935);
  not g20071 (n_10936, n11106);
  not g20072 (n_10937, n11137);
  and g20073 (n11138, n_10936, n_10937);
  and g20074 (n11139, n11106, n11137);
  not g20075 (n_10938, n11138);
  not g20076 (n_10939, n11139);
  and g20077 (n11140, n_10938, n_10939);
  not g20078 (n_10940, n11104);
  and g20079 (n11141, n_10940, n11140);
  not g20080 (n_10941, n11140);
  and g20081 (n11142, n11104, n_10941);
  not g20082 (n_10942, n11141);
  not g20083 (n_10943, n11142);
  and g20084 (n11143, n_10942, n_10943);
  not g20085 (n_10944, n11068);
  not g20086 (n_10945, n11143);
  and g20087 (n11144, n_10944, n_10945);
  and g20088 (n11145, n11068, n11143);
  not g20089 (n_10946, n11144);
  not g20090 (n_10947, n11145);
  and g20091 (n11146, n_10946, n_10947);
  not g20092 (n_10948, n11066);
  and g20093 (n11147, n_10948, n11146);
  not g20094 (n_10949, n11146);
  and g20095 (n11148, n11066, n_10949);
  not g20096 (n_10950, n11147);
  not g20097 (n_10951, n11148);
  and g20098 (n11149, n_10950, n_10951);
  not g20099 (n_10952, n10986);
  not g20100 (n_10953, n11149);
  and g20101 (n11150, n_10952, n_10953);
  and g20102 (n11151, n10986, n11149);
  not g20103 (n_10954, n11150);
  not g20104 (n_10955, n11151);
  and g20105 (n11152, n_10954, n_10955);
  not g20106 (n_10956, n10984);
  and g20107 (n11153, n_10956, n11152);
  not g20108 (n_10957, n11152);
  and g20109 (n11154, n10984, n_10957);
  not g20110 (n_10958, n11153);
  not g20111 (n_10959, n11154);
  and g20112 (n11155, n_10958, n_10959);
  not g20113 (n_10960, n10816);
  not g20114 (n_10961, n11155);
  and g20115 (n11156, n_10960, n_10961);
  and g20116 (n11157, n10816, n11155);
  not g20117 (n_10962, n11156);
  not g20118 (n_10963, n11157);
  and g20119 (n11158, n_10962, n_10963);
  not g20120 (n_10964, n10814);
  and g20121 (n11159, n_10964, n11158);
  not g20122 (n_10965, n11158);
  and g20123 (n11160, n10814, n_10965);
  not g20124 (n_10966, n11159);
  not g20125 (n_10967, n11160);
  and g20126 (n11161, n_10966, n_10967);
  not g20127 (n_10968, n10470);
  not g20128 (n_10969, n11161);
  and g20129 (n11162, n_10968, n_10969);
  and g20130 (n11163, n10470, n11161);
  not g20131 (n_10970, n11162);
  not g20132 (n_10971, n11163);
  and g20133 (n11164, n_10970, n_10971);
  not g20134 (n_10972, n10468);
  and g20135 (n11165, n_10972, n11164);
  not g20136 (n_10973, n11164);
  and g20137 (n11166, n10468, n_10973);
  not g20138 (n_10974, n11165);
  not g20139 (n_10975, n11166);
  and g20140 (n11167, n_10974, n_10975);
  not g20141 (n_10976, n10049);
  not g20142 (n_10977, n11167);
  and g20143 (n11168, n_10976, n_10977);
  and g20144 (n11169, n10049, n11167);
  not g20145 (n_10978, n11168);
  not g20146 (n_10979, n11169);
  and g20147 (n11170, n_10978, n_10979);
  and g20148 (n11171, n_3820, n_3818);
  not g20149 (n_10980, n11171);
  and g20150 (n11172, n_3819, n_10980);
  and g20151 (n11173, n_3813, n_3811);
  not g20152 (n_10981, n11173);
  and g20153 (n11174, n_3812, n_10981);
  and g20154 (n11175, n_3806, n_3804);
  not g20155 (n_10982, n11175);
  and g20156 (n11176, n_3805, n_10982);
  and g20157 (n11177, n_3799, n_3797);
  not g20158 (n_10983, n11177);
  and g20159 (n11178, n_3798, n_10983);
  and g20160 (n11179, n_3792, n_3790);
  not g20161 (n_10984, n11179);
  and g20162 (n11180, n_3791, n_10984);
  and g20163 (n11181, n4420, n_3784);
  not g20164 (n_10985, n11181);
  and g20165 (n11182, n_3785, n_10985);
  and g20166 (n11183, n_1944, n_1943);
  not g20167 (n_10986, n11183);
  and g20168 (n11184, n_1942, n_10986);
  and g20169 (n11185, n_1988, n_1986);
  not g20170 (n_10987, n11185);
  and g20171 (n11186, n_1987, n_10987);
  not g20172 (n_10988, n11184);
  and g20173 (n11187, n_10988, n11186);
  not g20174 (n_10989, n11186);
  and g20175 (n11188, n11184, n_10989);
  not g20176 (n_10990, n11187);
  not g20177 (n_10991, n11188);
  and g20178 (n11189, n_10990, n_10991);
  not g20179 (n_10992, n11182);
  not g20180 (n_10993, n11189);
  and g20181 (n11190, n_10992, n_10993);
  not g20185 (n_10994, n11190);
  not g20186 (n_10995, n11193);
  and g20187 (n11194, n_10994, n_10995);
  and g20188 (n11195, n4396, n_3763);
  not g20189 (n_10996, n11195);
  and g20190 (n11196, n_3764, n_10996);
  and g20191 (n11197, n_2036, n_2035);
  not g20192 (n_10997, n11197);
  and g20193 (n11198, n_2034, n_10997);
  and g20194 (n11199, n_2080, n_2079);
  not g20195 (n_10998, n11199);
  and g20196 (n11200, n_2078, n_10998);
  not g20197 (n_10999, n11198);
  and g20198 (n11201, n_10999, n11200);
  not g20199 (n_11000, n11200);
  and g20200 (n11202, n11198, n_11000);
  not g20201 (n_11001, n11201);
  not g20202 (n_11002, n11202);
  and g20203 (n11203, n_11001, n_11002);
  not g20204 (n_11003, n11196);
  not g20205 (n_11004, n11203);
  and g20206 (n11204, n_11003, n_11004);
  not g20210 (n_11005, n11204);
  not g20211 (n_11006, n11207);
  and g20212 (n11208, n_11005, n_11006);
  not g20213 (n_11007, n11194);
  and g20214 (n11209, n_11007, n11208);
  not g20215 (n_11008, n11208);
  and g20216 (n11210, n11194, n_11008);
  not g20217 (n_11009, n11209);
  not g20218 (n_11010, n11210);
  and g20219 (n11211, n_11009, n_11010);
  not g20220 (n_11011, n11180);
  not g20221 (n_11012, n11211);
  and g20222 (n11212, n_11011, n_11012);
  and g20223 (n11213, n11180, n11211);
  not g20224 (n_11013, n11212);
  not g20225 (n_11014, n11213);
  and g20226 (n11214, n_11013, n_11014);
  and g20227 (n11215, n_3748, n_3746);
  not g20228 (n_11015, n11215);
  and g20229 (n11216, n_3747, n_11015);
  and g20230 (n11217, n4341, n_3726);
  not g20231 (n_11016, n11217);
  and g20232 (n11218, n_3727, n_11016);
  and g20233 (n11219, n_2224, n_2223);
  not g20234 (n_11017, n11219);
  and g20235 (n11220, n_2222, n_11017);
  and g20236 (n11221, n_2268, n_2267);
  not g20237 (n_11018, n11221);
  and g20238 (n11222, n_2266, n_11018);
  not g20239 (n_11019, n11220);
  and g20240 (n11223, n_11019, n11222);
  not g20241 (n_11020, n11222);
  and g20242 (n11224, n11220, n_11020);
  not g20243 (n_11021, n11223);
  not g20244 (n_11022, n11224);
  and g20245 (n11225, n_11021, n_11022);
  not g20246 (n_11023, n11218);
  not g20247 (n_11024, n11225);
  and g20248 (n11226, n_11023, n_11024);
  not g20252 (n_11025, n11226);
  not g20253 (n_11026, n11229);
  and g20254 (n11230, n_11025, n_11026);
  and g20255 (n11231, n4360, n_3735);
  not g20256 (n_11027, n11231);
  and g20257 (n11232, n_3736, n_11027);
  and g20258 (n11233, n_2132, n_2131);
  not g20259 (n_11028, n11233);
  and g20260 (n11234, n_2130, n_11028);
  and g20261 (n11235, n_2176, n_2175);
  not g20262 (n_11029, n11235);
  and g20263 (n11236, n_2174, n_11029);
  not g20264 (n_11030, n11234);
  and g20265 (n11237, n_11030, n11236);
  not g20266 (n_11031, n11236);
  and g20267 (n11238, n11234, n_11031);
  not g20268 (n_11032, n11237);
  not g20269 (n_11033, n11238);
  and g20270 (n11239, n_11032, n_11033);
  not g20271 (n_11034, n11232);
  not g20272 (n_11035, n11239);
  and g20273 (n11240, n_11034, n_11035);
  not g20277 (n_11036, n11240);
  not g20278 (n_11037, n11243);
  and g20279 (n11244, n_11036, n_11037);
  not g20280 (n_11038, n11230);
  and g20281 (n11245, n_11038, n11244);
  not g20282 (n_11039, n11244);
  and g20283 (n11246, n11230, n_11039);
  not g20284 (n_11040, n11245);
  not g20285 (n_11041, n11246);
  and g20286 (n11247, n_11040, n_11041);
  not g20287 (n_11042, n11216);
  not g20288 (n_11043, n11247);
  and g20289 (n11248, n_11042, n_11043);
  and g20290 (n11249, n11216, n11247);
  not g20291 (n_11044, n11248);
  not g20292 (n_11045, n11249);
  and g20293 (n11250, n_11044, n_11045);
  not g20294 (n_11046, n11214);
  and g20295 (n11251, n_11046, n11250);
  not g20296 (n_11047, n11250);
  and g20297 (n11252, n11214, n_11047);
  not g20298 (n_11048, n11251);
  not g20299 (n_11049, n11252);
  and g20300 (n11253, n_11048, n_11049);
  not g20301 (n_11050, n11178);
  not g20302 (n_11051, n11253);
  and g20303 (n11254, n_11050, n_11051);
  and g20304 (n11255, n11178, n11253);
  not g20305 (n_11052, n11254);
  not g20306 (n_11053, n11255);
  and g20307 (n11256, n_11052, n_11053);
  and g20308 (n11257, n_3707, n_3705);
  not g20309 (n_11054, n11257);
  and g20310 (n11258, n_3706, n_11054);
  and g20311 (n11259, n_3662, n_3660);
  not g20312 (n_11055, n11259);
  and g20313 (n11260, n_3661, n_11055);
  and g20314 (n11261, n4248, n_3654);
  not g20315 (n_11056, n11261);
  and g20316 (n11262, n_3655, n_11056);
  and g20317 (n11263, n_2604, n_2603);
  not g20318 (n_11057, n11263);
  and g20319 (n11264, n_2602, n_11057);
  and g20320 (n11265, n_2648, n_2647);
  not g20321 (n_11058, n11265);
  and g20322 (n11266, n_2646, n_11058);
  not g20323 (n_11059, n11264);
  and g20324 (n11267, n_11059, n11266);
  not g20325 (n_11060, n11266);
  and g20326 (n11268, n11264, n_11060);
  not g20327 (n_11061, n11267);
  not g20328 (n_11062, n11268);
  and g20329 (n11269, n_11061, n_11062);
  not g20330 (n_11063, n11262);
  not g20331 (n_11064, n11269);
  and g20332 (n11270, n_11063, n_11064);
  not g20336 (n_11065, n11270);
  not g20337 (n_11066, n11273);
  and g20338 (n11274, n_11065, n_11066);
  and g20339 (n11275, n4224, n_3633);
  not g20340 (n_11067, n11275);
  and g20341 (n11276, n_3634, n_11067);
  and g20342 (n11277, n_2512, n_2511);
  not g20343 (n_11068, n11277);
  and g20344 (n11278, n_2510, n_11068);
  and g20345 (n11279, n_2556, n_2555);
  not g20346 (n_11069, n11279);
  and g20347 (n11280, n_2554, n_11069);
  not g20348 (n_11070, n11278);
  and g20349 (n11281, n_11070, n11280);
  not g20350 (n_11071, n11280);
  and g20351 (n11282, n11278, n_11071);
  not g20352 (n_11072, n11281);
  not g20353 (n_11073, n11282);
  and g20354 (n11283, n_11072, n_11073);
  not g20355 (n_11074, n11276);
  not g20356 (n_11075, n11283);
  and g20357 (n11284, n_11074, n_11075);
  not g20361 (n_11076, n11284);
  not g20362 (n_11077, n11287);
  and g20363 (n11288, n_11076, n_11077);
  not g20364 (n_11078, n11274);
  and g20365 (n11289, n_11078, n11288);
  not g20366 (n_11079, n11288);
  and g20367 (n11290, n11274, n_11079);
  not g20368 (n_11080, n11289);
  not g20369 (n_11081, n11290);
  and g20370 (n11291, n_11080, n_11081);
  not g20371 (n_11082, n11260);
  not g20372 (n_11083, n11291);
  and g20373 (n11292, n_11082, n_11083);
  and g20374 (n11293, n11260, n11291);
  not g20375 (n_11084, n11292);
  not g20376 (n_11085, n11293);
  and g20377 (n11294, n_11084, n_11085);
  and g20378 (n11295, n_3696, n_3694);
  not g20379 (n_11086, n11295);
  and g20380 (n11296, n_3695, n_11086);
  and g20381 (n11297, n4274, n_3674);
  not g20382 (n_11087, n11297);
  and g20383 (n11298, n_3675, n_11087);
  and g20384 (n11299, n_2416, n_2415);
  not g20385 (n_11088, n11299);
  and g20386 (n11300, n_2414, n_11088);
  and g20387 (n11301, n_2460, n_2459);
  not g20388 (n_11089, n11301);
  and g20389 (n11302, n_2458, n_11089);
  not g20390 (n_11090, n11300);
  and g20391 (n11303, n_11090, n11302);
  not g20392 (n_11091, n11302);
  and g20393 (n11304, n11300, n_11091);
  not g20394 (n_11092, n11303);
  not g20395 (n_11093, n11304);
  and g20396 (n11305, n_11092, n_11093);
  not g20397 (n_11094, n11298);
  not g20398 (n_11095, n11305);
  and g20399 (n11306, n_11094, n_11095);
  not g20403 (n_11096, n11306);
  not g20404 (n_11097, n11309);
  and g20405 (n11310, n_11096, n_11097);
  and g20406 (n11311, n4293, n_3683);
  not g20407 (n_11098, n11311);
  and g20408 (n11312, n_3684, n_11098);
  and g20409 (n11313, n_2324, n_2323);
  not g20410 (n_11099, n11313);
  and g20411 (n11314, n_2322, n_11099);
  and g20412 (n11315, n_2368, n_2367);
  not g20413 (n_11100, n11315);
  and g20414 (n11316, n_2366, n_11100);
  not g20415 (n_11101, n11314);
  and g20416 (n11317, n_11101, n11316);
  not g20417 (n_11102, n11316);
  and g20418 (n11318, n11314, n_11102);
  not g20419 (n_11103, n11317);
  not g20420 (n_11104, n11318);
  and g20421 (n11319, n_11103, n_11104);
  not g20422 (n_11105, n11312);
  not g20423 (n_11106, n11319);
  and g20424 (n11320, n_11105, n_11106);
  not g20428 (n_11107, n11320);
  not g20429 (n_11108, n11323);
  and g20430 (n11324, n_11107, n_11108);
  not g20431 (n_11109, n11310);
  and g20432 (n11325, n_11109, n11324);
  not g20433 (n_11110, n11324);
  and g20434 (n11326, n11310, n_11110);
  not g20435 (n_11111, n11325);
  not g20436 (n_11112, n11326);
  and g20437 (n11327, n_11111, n_11112);
  not g20438 (n_11113, n11296);
  not g20439 (n_11114, n11327);
  and g20440 (n11328, n_11113, n_11114);
  and g20441 (n11329, n11296, n11327);
  not g20442 (n_11115, n11328);
  not g20443 (n_11116, n11329);
  and g20444 (n11330, n_11115, n_11116);
  not g20445 (n_11117, n11294);
  and g20446 (n11331, n_11117, n11330);
  not g20447 (n_11118, n11330);
  and g20448 (n11332, n11294, n_11118);
  not g20449 (n_11119, n11331);
  not g20450 (n_11120, n11332);
  and g20451 (n11333, n_11119, n_11120);
  not g20452 (n_11121, n11258);
  not g20453 (n_11122, n11333);
  and g20454 (n11334, n_11121, n_11122);
  and g20455 (n11335, n11258, n11333);
  not g20456 (n_11123, n11334);
  not g20457 (n_11124, n11335);
  and g20458 (n11336, n_11123, n_11124);
  not g20459 (n_11125, n11256);
  and g20460 (n11337, n_11125, n11336);
  not g20461 (n_11126, n11336);
  and g20462 (n11338, n11256, n_11126);
  not g20463 (n_11127, n11337);
  not g20464 (n_11128, n11338);
  and g20465 (n11339, n_11127, n_11128);
  not g20466 (n_11129, n11176);
  not g20467 (n_11130, n11339);
  and g20468 (n11340, n_11129, n_11130);
  and g20469 (n11341, n11176, n11339);
  not g20470 (n_11131, n11340);
  not g20471 (n_11132, n11341);
  and g20472 (n11342, n_11131, n_11132);
  and g20473 (n11343, n_3618, n_3616);
  not g20474 (n_11133, n11343);
  and g20475 (n11344, n_3617, n_11133);
  and g20476 (n11345, n_3525, n_3523);
  not g20477 (n_11134, n11345);
  and g20478 (n11346, n_3524, n_11134);
  and g20479 (n11347, n_3518, n_3516);
  not g20480 (n_11135, n11347);
  and g20481 (n11348, n_3517, n_11135);
  and g20482 (n11349, n4062, n_3510);
  not g20483 (n_11136, n11349);
  and g20484 (n11350, n_3511, n_11136);
  and g20485 (n11351, n_3368, n_3367);
  not g20486 (n_11137, n11351);
  and g20487 (n11352, n_3366, n_11137);
  and g20488 (n11353, n_3412, n_3411);
  not g20489 (n_11138, n11353);
  and g20490 (n11354, n_3410, n_11138);
  not g20491 (n_11139, n11352);
  and g20492 (n11355, n_11139, n11354);
  not g20493 (n_11140, n11354);
  and g20494 (n11356, n11352, n_11140);
  not g20495 (n_11141, n11355);
  not g20496 (n_11142, n11356);
  and g20497 (n11357, n_11141, n_11142);
  not g20498 (n_11143, n11350);
  not g20499 (n_11144, n11357);
  and g20500 (n11358, n_11143, n_11144);
  not g20504 (n_11145, n11358);
  not g20505 (n_11146, n11361);
  and g20506 (n11362, n_11145, n_11146);
  and g20507 (n11363, n4038, n_3489);
  not g20508 (n_11147, n11363);
  and g20509 (n11364, n_3490, n_11147);
  and g20510 (n11365, n_3276, n_3275);
  not g20511 (n_11148, n11365);
  and g20512 (n11366, n_3274, n_11148);
  and g20513 (n11367, n_3320, n_3319);
  not g20514 (n_11149, n11367);
  and g20515 (n11368, n_3318, n_11149);
  not g20516 (n_11150, n11366);
  and g20517 (n11369, n_11150, n11368);
  not g20518 (n_11151, n11368);
  and g20519 (n11370, n11366, n_11151);
  not g20520 (n_11152, n11369);
  not g20521 (n_11153, n11370);
  and g20522 (n11371, n_11152, n_11153);
  not g20523 (n_11154, n11364);
  not g20524 (n_11155, n11371);
  and g20525 (n11372, n_11154, n_11155);
  not g20529 (n_11156, n11372);
  not g20530 (n_11157, n11375);
  and g20531 (n11376, n_11156, n_11157);
  not g20532 (n_11158, n11362);
  and g20533 (n11377, n_11158, n11376);
  not g20534 (n_11159, n11376);
  and g20535 (n11378, n11362, n_11159);
  not g20536 (n_11160, n11377);
  not g20537 (n_11161, n11378);
  and g20538 (n11379, n_11160, n_11161);
  not g20539 (n_11162, n11348);
  not g20540 (n_11163, n11379);
  and g20541 (n11380, n_11162, n_11163);
  and g20542 (n11381, n11348, n11379);
  not g20543 (n_11164, n11380);
  not g20544 (n_11165, n11381);
  and g20545 (n11382, n_11164, n_11165);
  and g20546 (n11383, n_3474, n_3472);
  not g20547 (n_11166, n11383);
  and g20548 (n11384, n_3473, n_11166);
  and g20549 (n11385, n3983, n_3452);
  not g20550 (n_11167, n11385);
  and g20551 (n11386, n_3453, n_11167);
  and g20552 (n11387, n_3180, n_3179);
  not g20553 (n_11168, n11387);
  and g20554 (n11388, n_3178, n_11168);
  and g20555 (n11389, n_3224, n_3223);
  not g20556 (n_11169, n11389);
  and g20557 (n11390, n_3222, n_11169);
  not g20558 (n_11170, n11388);
  and g20559 (n11391, n_11170, n11390);
  not g20560 (n_11171, n11390);
  and g20561 (n11392, n11388, n_11171);
  not g20562 (n_11172, n11391);
  not g20563 (n_11173, n11392);
  and g20564 (n11393, n_11172, n_11173);
  not g20565 (n_11174, n11386);
  not g20566 (n_11175, n11393);
  and g20567 (n11394, n_11174, n_11175);
  not g20571 (n_11176, n11394);
  not g20572 (n_11177, n11397);
  and g20573 (n11398, n_11176, n_11177);
  and g20574 (n11399, n4002, n_3461);
  not g20575 (n_11178, n11399);
  and g20576 (n11400, n_3462, n_11178);
  and g20577 (n11401, n_3088, n_3087);
  not g20578 (n_11179, n11401);
  and g20579 (n11402, n_3086, n_11179);
  and g20580 (n11403, n_3132, n_3131);
  not g20581 (n_11180, n11403);
  and g20582 (n11404, n_3130, n_11180);
  not g20583 (n_11181, n11402);
  and g20584 (n11405, n_11181, n11404);
  not g20585 (n_11182, n11404);
  and g20586 (n11406, n11402, n_11182);
  not g20587 (n_11183, n11405);
  not g20588 (n_11184, n11406);
  and g20589 (n11407, n_11183, n_11184);
  not g20590 (n_11185, n11400);
  not g20591 (n_11186, n11407);
  and g20592 (n11408, n_11185, n_11186);
  not g20596 (n_11187, n11408);
  not g20597 (n_11188, n11411);
  and g20598 (n11412, n_11187, n_11188);
  not g20599 (n_11189, n11398);
  and g20600 (n11413, n_11189, n11412);
  not g20601 (n_11190, n11412);
  and g20602 (n11414, n11398, n_11190);
  not g20603 (n_11191, n11413);
  not g20604 (n_11192, n11414);
  and g20605 (n11415, n_11191, n_11192);
  not g20606 (n_11193, n11384);
  not g20607 (n_11194, n11415);
  and g20608 (n11416, n_11193, n_11194);
  and g20609 (n11417, n11384, n11415);
  not g20610 (n_11195, n11416);
  not g20611 (n_11196, n11417);
  and g20612 (n11418, n_11195, n_11196);
  not g20613 (n_11197, n11382);
  and g20614 (n11419, n_11197, n11418);
  not g20615 (n_11198, n11418);
  and g20616 (n11420, n11382, n_11198);
  not g20617 (n_11199, n11419);
  not g20618 (n_11200, n11420);
  and g20619 (n11421, n_11199, n_11200);
  not g20620 (n_11201, n11346);
  not g20621 (n_11202, n11421);
  and g20622 (n11422, n_11201, n_11202);
  and g20623 (n11423, n11346, n11421);
  not g20624 (n_11203, n11422);
  not g20625 (n_11204, n11423);
  and g20626 (n11424, n_11203, n_11204);
  and g20627 (n11425, n_3607, n_3605);
  not g20628 (n_11205, n11425);
  and g20629 (n11426, n_3606, n_11205);
  and g20630 (n11427, n_3562, n_3560);
  not g20631 (n_11206, n11427);
  and g20632 (n11428, n_3561, n_11206);
  and g20633 (n11429, n4119, n_3554);
  not g20634 (n_11207, n11429);
  and g20635 (n11430, n_3555, n_11207);
  and g20636 (n11431, n_2988, n_2987);
  not g20637 (n_11208, n11431);
  and g20638 (n11432, n_2986, n_11208);
  and g20639 (n11433, n_3032, n_3031);
  not g20640 (n_11209, n11433);
  and g20641 (n11434, n_3030, n_11209);
  not g20642 (n_11210, n11432);
  and g20643 (n11435, n_11210, n11434);
  not g20644 (n_11211, n11434);
  and g20645 (n11436, n11432, n_11211);
  not g20646 (n_11212, n11435);
  not g20647 (n_11213, n11436);
  and g20648 (n11437, n_11212, n_11213);
  not g20649 (n_11214, n11430);
  not g20650 (n_11215, n11437);
  and g20651 (n11438, n_11214, n_11215);
  not g20655 (n_11216, n11438);
  not g20656 (n_11217, n11441);
  and g20657 (n11442, n_11216, n_11217);
  and g20658 (n11443, n4095, n_3533);
  not g20659 (n_11218, n11443);
  and g20660 (n11444, n_3534, n_11218);
  and g20661 (n11445, n_2896, n_2895);
  not g20662 (n_11219, n11445);
  and g20663 (n11446, n_2894, n_11219);
  and g20664 (n11447, n_2940, n_2939);
  not g20665 (n_11220, n11447);
  and g20666 (n11448, n_2938, n_11220);
  not g20667 (n_11221, n11446);
  and g20668 (n11449, n_11221, n11448);
  not g20669 (n_11222, n11448);
  and g20670 (n11450, n11446, n_11222);
  not g20671 (n_11223, n11449);
  not g20672 (n_11224, n11450);
  and g20673 (n11451, n_11223, n_11224);
  not g20674 (n_11225, n11444);
  not g20675 (n_11226, n11451);
  and g20676 (n11452, n_11225, n_11226);
  not g20680 (n_11227, n11452);
  not g20681 (n_11228, n11455);
  and g20682 (n11456, n_11227, n_11228);
  not g20683 (n_11229, n11442);
  and g20684 (n11457, n_11229, n11456);
  not g20685 (n_11230, n11456);
  and g20686 (n11458, n11442, n_11230);
  not g20687 (n_11231, n11457);
  not g20688 (n_11232, n11458);
  and g20689 (n11459, n_11231, n_11232);
  not g20690 (n_11233, n11428);
  not g20691 (n_11234, n11459);
  and g20692 (n11460, n_11233, n_11234);
  and g20693 (n11461, n11428, n11459);
  not g20694 (n_11235, n11460);
  not g20695 (n_11236, n11461);
  and g20696 (n11462, n_11235, n_11236);
  and g20697 (n11463, n_3596, n_3594);
  not g20698 (n_11237, n11463);
  and g20699 (n11464, n_3595, n_11237);
  and g20700 (n11465, n4145, n_3574);
  not g20701 (n_11238, n11465);
  and g20702 (n11466, n_3575, n_11238);
  and g20703 (n11467, n_2800, n_2799);
  not g20704 (n_11239, n11467);
  and g20705 (n11468, n_2798, n_11239);
  and g20706 (n11469, n_2844, n_2843);
  not g20707 (n_11240, n11469);
  and g20708 (n11470, n_2842, n_11240);
  not g20709 (n_11241, n11468);
  and g20710 (n11471, n_11241, n11470);
  not g20711 (n_11242, n11470);
  and g20712 (n11472, n11468, n_11242);
  not g20713 (n_11243, n11471);
  not g20714 (n_11244, n11472);
  and g20715 (n11473, n_11243, n_11244);
  not g20716 (n_11245, n11466);
  not g20717 (n_11246, n11473);
  and g20718 (n11474, n_11245, n_11246);
  not g20722 (n_11247, n11474);
  not g20723 (n_11248, n11477);
  and g20724 (n11478, n_11247, n_11248);
  and g20725 (n11479, n4164, n_3583);
  not g20726 (n_11249, n11479);
  and g20727 (n11480, n_3584, n_11249);
  and g20728 (n11481, n_2708, n_2707);
  not g20729 (n_11250, n11481);
  and g20730 (n11482, n_2706, n_11250);
  and g20731 (n11483, n_2752, n_2751);
  not g20732 (n_11251, n11483);
  and g20733 (n11484, n_2750, n_11251);
  not g20734 (n_11252, n11482);
  and g20735 (n11485, n_11252, n11484);
  not g20736 (n_11253, n11484);
  and g20737 (n11486, n11482, n_11253);
  not g20738 (n_11254, n11485);
  not g20739 (n_11255, n11486);
  and g20740 (n11487, n_11254, n_11255);
  not g20741 (n_11256, n11480);
  not g20742 (n_11257, n11487);
  and g20743 (n11488, n_11256, n_11257);
  not g20747 (n_11258, n11488);
  not g20748 (n_11259, n11491);
  and g20749 (n11492, n_11258, n_11259);
  not g20750 (n_11260, n11478);
  and g20751 (n11493, n_11260, n11492);
  not g20752 (n_11261, n11492);
  and g20753 (n11494, n11478, n_11261);
  not g20754 (n_11262, n11493);
  not g20755 (n_11263, n11494);
  and g20756 (n11495, n_11262, n_11263);
  not g20757 (n_11264, n11464);
  not g20758 (n_11265, n11495);
  and g20759 (n11496, n_11264, n_11265);
  and g20760 (n11497, n11464, n11495);
  not g20761 (n_11266, n11496);
  not g20762 (n_11267, n11497);
  and g20763 (n11498, n_11266, n_11267);
  not g20764 (n_11268, n11462);
  and g20765 (n11499, n_11268, n11498);
  not g20766 (n_11269, n11498);
  and g20767 (n11500, n11462, n_11269);
  not g20768 (n_11270, n11499);
  not g20769 (n_11271, n11500);
  and g20770 (n11501, n_11270, n_11271);
  not g20771 (n_11272, n11426);
  not g20772 (n_11273, n11501);
  and g20773 (n11502, n_11272, n_11273);
  and g20774 (n11503, n11426, n11501);
  not g20775 (n_11274, n11502);
  not g20776 (n_11275, n11503);
  and g20777 (n11504, n_11274, n_11275);
  not g20778 (n_11276, n11424);
  and g20779 (n11505, n_11276, n11504);
  not g20780 (n_11277, n11504);
  and g20781 (n11506, n11424, n_11277);
  not g20782 (n_11278, n11505);
  not g20783 (n_11279, n11506);
  and g20784 (n11507, n_11278, n_11279);
  not g20785 (n_11280, n11344);
  not g20786 (n_11281, n11507);
  and g20787 (n11508, n_11280, n_11281);
  and g20788 (n11509, n11344, n11507);
  not g20789 (n_11282, n11508);
  not g20790 (n_11283, n11509);
  and g20791 (n11510, n_11282, n_11283);
  not g20792 (n_11284, n11342);
  and g20793 (n11511, n_11284, n11510);
  not g20794 (n_11285, n11510);
  and g20795 (n11512, n11342, n_11285);
  not g20796 (n_11286, n11511);
  not g20797 (n_11287, n11512);
  and g20798 (n11513, n_11286, n_11287);
  not g20799 (n_11288, n11174);
  not g20800 (n_11289, n11513);
  and g20801 (n11514, n_11288, n_11289);
  and g20802 (n11515, n11174, n11513);
  not g20803 (n_11290, n11514);
  not g20804 (n_11291, n11515);
  and g20805 (n11516, n_11290, n_11291);
  and g20806 (n11517, n_1897, n_1895);
  not g20807 (n_11292, n11517);
  and g20808 (n11518, n_1896, n_11292);
  and g20809 (n11519, n_940, n_938);
  not g20810 (n_11293, n11519);
  and g20811 (n11520, n_939, n_11293);
  and g20812 (n11521, n_933, n_931);
  not g20813 (n_11294, n11521);
  and g20814 (n11522, n_932, n_11294);
  and g20815 (n11523, n_926, n_924);
  not g20816 (n_11295, n11523);
  and g20817 (n11524, n_925, n_11295);
  and g20818 (n11525, n1818, n_918);
  not g20819 (n_11296, n11525);
  and g20820 (n11526, n_919, n_11296);
  and g20821 (n11527, n_786, n_785);
  not g20822 (n_11297, n11527);
  and g20823 (n11528, n_784, n_11297);
  and g20824 (n11529, n_830, n_829);
  not g20825 (n_11298, n11529);
  and g20826 (n11530, n_828, n_11298);
  not g20827 (n_11299, n11528);
  and g20828 (n11531, n_11299, n11530);
  not g20829 (n_11300, n11530);
  and g20830 (n11532, n11528, n_11300);
  not g20831 (n_11301, n11531);
  not g20832 (n_11302, n11532);
  and g20833 (n11533, n_11301, n_11302);
  not g20834 (n_11303, n11526);
  not g20835 (n_11304, n11533);
  and g20836 (n11534, n_11303, n_11304);
  not g20840 (n_11305, n11534);
  not g20841 (n_11306, n11537);
  and g20842 (n11538, n_11305, n_11306);
  and g20843 (n11539, n1794, n_897);
  not g20844 (n_11307, n11539);
  and g20845 (n11540, n_898, n_11307);
  and g20846 (n11541, n_694, n_693);
  not g20847 (n_11308, n11541);
  and g20848 (n11542, n_692, n_11308);
  and g20849 (n11543, n_738, n_737);
  not g20850 (n_11309, n11543);
  and g20851 (n11544, n_736, n_11309);
  not g20852 (n_11310, n11542);
  and g20853 (n11545, n_11310, n11544);
  not g20854 (n_11311, n11544);
  and g20855 (n11546, n11542, n_11311);
  not g20856 (n_11312, n11545);
  not g20857 (n_11313, n11546);
  and g20858 (n11547, n_11312, n_11313);
  not g20859 (n_11314, n11540);
  not g20860 (n_11315, n11547);
  and g20861 (n11548, n_11314, n_11315);
  not g20865 (n_11316, n11548);
  not g20866 (n_11317, n11551);
  and g20867 (n11552, n_11316, n_11317);
  not g20868 (n_11318, n11538);
  and g20869 (n11553, n_11318, n11552);
  not g20870 (n_11319, n11552);
  and g20871 (n11554, n11538, n_11319);
  not g20872 (n_11320, n11553);
  not g20873 (n_11321, n11554);
  and g20874 (n11555, n_11320, n_11321);
  not g20875 (n_11322, n11524);
  not g20876 (n_11323, n11555);
  and g20877 (n11556, n_11322, n_11323);
  and g20878 (n11557, n11524, n11555);
  not g20879 (n_11324, n11556);
  not g20880 (n_11325, n11557);
  and g20881 (n11558, n_11324, n_11325);
  and g20882 (n11559, n_882, n_880);
  not g20883 (n_11326, n11559);
  and g20884 (n11560, n_881, n_11326);
  and g20885 (n11561, n1739, n_860);
  not g20886 (n_11327, n11561);
  and g20887 (n11562, n_861, n_11327);
  and g20888 (n11563, n_598, n_597);
  not g20889 (n_11328, n11563);
  and g20890 (n11564, n_596, n_11328);
  and g20891 (n11565, n_642, n_641);
  not g20892 (n_11329, n11565);
  and g20893 (n11566, n_640, n_11329);
  not g20894 (n_11330, n11564);
  and g20895 (n11567, n_11330, n11566);
  not g20896 (n_11331, n11566);
  and g20897 (n11568, n11564, n_11331);
  not g20898 (n_11332, n11567);
  not g20899 (n_11333, n11568);
  and g20900 (n11569, n_11332, n_11333);
  not g20901 (n_11334, n11562);
  not g20902 (n_11335, n11569);
  and g20903 (n11570, n_11334, n_11335);
  not g20907 (n_11336, n11570);
  not g20908 (n_11337, n11573);
  and g20909 (n11574, n_11336, n_11337);
  and g20910 (n11575, n1758, n_869);
  not g20911 (n_11338, n11575);
  and g20912 (n11576, n_870, n_11338);
  and g20913 (n11577, n_506, n_505);
  not g20914 (n_11339, n11577);
  and g20915 (n11578, n_504, n_11339);
  and g20916 (n11579, n_550, n_549);
  not g20917 (n_11340, n11579);
  and g20918 (n11580, n_548, n_11340);
  not g20919 (n_11341, n11578);
  and g20920 (n11581, n_11341, n11580);
  not g20921 (n_11342, n11580);
  and g20922 (n11582, n11578, n_11342);
  not g20923 (n_11343, n11581);
  not g20924 (n_11344, n11582);
  and g20925 (n11583, n_11343, n_11344);
  not g20926 (n_11345, n11576);
  not g20927 (n_11346, n11583);
  and g20928 (n11584, n_11345, n_11346);
  not g20932 (n_11347, n11584);
  not g20933 (n_11348, n11587);
  and g20934 (n11588, n_11347, n_11348);
  not g20935 (n_11349, n11574);
  and g20936 (n11589, n_11349, n11588);
  not g20937 (n_11350, n11588);
  and g20938 (n11590, n11574, n_11350);
  not g20939 (n_11351, n11589);
  not g20940 (n_11352, n11590);
  and g20941 (n11591, n_11351, n_11352);
  not g20942 (n_11353, n11560);
  not g20943 (n_11354, n11591);
  and g20944 (n11592, n_11353, n_11354);
  and g20945 (n11593, n11560, n11591);
  not g20946 (n_11355, n11592);
  not g20947 (n_11356, n11593);
  and g20948 (n11594, n_11355, n_11356);
  not g20949 (n_11357, n11558);
  and g20950 (n11595, n_11357, n11594);
  not g20951 (n_11358, n11594);
  and g20952 (n11596, n11558, n_11358);
  not g20953 (n_11359, n11595);
  not g20954 (n_11360, n11596);
  and g20955 (n11597, n_11359, n_11360);
  not g20956 (n_11361, n11522);
  not g20957 (n_11362, n11597);
  and g20958 (n11598, n_11361, n_11362);
  and g20959 (n11599, n11522, n11597);
  not g20960 (n_11363, n11598);
  not g20961 (n_11364, n11599);
  and g20962 (n11600, n_11363, n_11364);
  and g20963 (n11601, n_457, n_455);
  not g20964 (n_11365, n11601);
  and g20965 (n11602, n_456, n_11365);
  and g20966 (n11603, n_220, n_218);
  not g20967 (n_11366, n11603);
  and g20968 (n11604, n_219, n_11366);
  and g20969 (n11605, n1178, n_212);
  not g20970 (n_11367, n11605);
  and g20971 (n11606, n_213, n_11367);
  and g20972 (n11607, n_146, n_145);
  not g20973 (n_11368, n11607);
  and g20974 (n11608, n_144, n_11368);
  and g20975 (n11609, n_190, n_189);
  not g20976 (n_11369, n11609);
  and g20977 (n11610, n_188, n_11369);
  not g20978 (n_11370, n11608);
  and g20979 (n11611, n_11370, n11610);
  not g20980 (n_11371, n11610);
  and g20981 (n11612, n11608, n_11371);
  not g20982 (n_11372, n11611);
  not g20983 (n_11373, n11612);
  and g20984 (n11613, n_11372, n_11373);
  not g20985 (n_11374, n11606);
  not g20986 (n_11375, n11613);
  and g20987 (n11614, n_11374, n_11375);
  not g20991 (n_11376, n11614);
  not g20992 (n_11377, n11617);
  and g20993 (n11618, n_11376, n_11377);
  and g20994 (n11619, n1038, n_93);
  not g20995 (n_11378, n11619);
  and g20996 (n11620, n_94, n_11378);
  and g20997 (n11621, n_84, n_87);
  not g20998 (n_11379, n11621);
  and g20999 (n11622, n_83, n_11379);
  and g21000 (n11623, n_43, n_41);
  not g21001 (n_11380, n11623);
  and g21002 (n11624, n_42, n_11380);
  not g21003 (n_11381, n11622);
  and g21004 (n11625, n_11381, n11624);
  not g21005 (n_11382, n11624);
  and g21006 (n11626, n11622, n_11382);
  not g21007 (n_11383, n11625);
  not g21008 (n_11384, n11626);
  and g21009 (n11627, n_11383, n_11384);
  not g21010 (n_11385, n11620);
  not g21011 (n_11386, n11627);
  and g21012 (n11628, n_11385, n_11386);
  not g21016 (n_11387, n11628);
  not g21017 (n_11388, n11631);
  and g21018 (n11632, n_11387, n_11388);
  not g21019 (n_11389, n11618);
  and g21020 (n11633, n_11389, n11632);
  not g21021 (n_11390, n11632);
  and g21022 (n11634, n11618, n_11390);
  not g21023 (n_11391, n11633);
  not g21024 (n_11392, n11634);
  and g21025 (n11635, n_11391, n_11392);
  not g21026 (n_11393, n11604);
  not g21027 (n_11394, n11635);
  and g21028 (n11636, n_11393, n_11394);
  and g21029 (n11637, n11604, n11635);
  not g21030 (n_11395, n11636);
  not g21031 (n_11396, n11637);
  and g21032 (n11638, n_11395, n_11396);
  and g21033 (n11639, n_440, n_438);
  not g21034 (n_11397, n11639);
  and g21035 (n11640, n_439, n_11397);
  and g21036 (n11641, n1238, n_320);
  not g21037 (n_11398, n11641);
  and g21038 (n11642, n_321, n_11398);
  and g21039 (n11643, n_307, n_310);
  not g21040 (n_11399, n11643);
  and g21041 (n11644, n_306, n_11399);
  and g21042 (n11645, n_266, n_264);
  not g21043 (n_11400, n11645);
  and g21044 (n11646, n_265, n_11400);
  not g21045 (n_11401, n11644);
  and g21046 (n11647, n_11401, n11646);
  not g21047 (n_11402, n11646);
  and g21048 (n11648, n11644, n_11402);
  not g21049 (n_11403, n11647);
  not g21050 (n_11404, n11648);
  and g21051 (n11649, n_11403, n_11404);
  not g21052 (n_11405, n11642);
  not g21053 (n_11406, n11649);
  and g21054 (n11650, n_11405, n_11406);
  not g21058 (n_11407, n11650);
  not g21059 (n_11408, n11653);
  and g21060 (n11654, n_11407, n_11408);
  and g21061 (n11655, n1327, n_417);
  not g21062 (n_11409, n11655);
  and g21063 (n11656, n_418, n_11409);
  and g21064 (n11657, n_408, n_411);
  not g21065 (n_11410, n11657);
  and g21066 (n11658, n_407, n_11410);
  and g21067 (n11659, n_367, n_365);
  not g21068 (n_11411, n11659);
  and g21069 (n11660, n_366, n_11411);
  not g21070 (n_11412, n11658);
  and g21071 (n11661, n_11412, n11660);
  not g21072 (n_11413, n11660);
  and g21073 (n11662, n11658, n_11413);
  not g21074 (n_11414, n11661);
  not g21075 (n_11415, n11662);
  and g21076 (n11663, n_11414, n_11415);
  not g21077 (n_11416, n11656);
  not g21078 (n_11417, n11663);
  and g21079 (n11664, n_11416, n_11417);
  not g21083 (n_11418, n11664);
  not g21084 (n_11419, n11667);
  and g21085 (n11668, n_11418, n_11419);
  not g21086 (n_11420, n11654);
  and g21087 (n11669, n_11420, n11668);
  not g21088 (n_11421, n11668);
  and g21089 (n11670, n11654, n_11421);
  not g21090 (n_11422, n11669);
  not g21091 (n_11423, n11670);
  and g21092 (n11671, n_11422, n_11423);
  not g21093 (n_11424, n11640);
  not g21094 (n_11425, n11671);
  and g21095 (n11672, n_11424, n_11425);
  and g21096 (n11673, n11640, n11671);
  not g21097 (n_11426, n11672);
  not g21098 (n_11427, n11673);
  and g21099 (n11674, n_11426, n_11427);
  not g21100 (n_11428, n11638);
  and g21101 (n11675, n_11428, n11674);
  not g21102 (n_11429, n11674);
  and g21103 (n11676, n11638, n_11429);
  not g21104 (n_11430, n11675);
  not g21105 (n_11431, n11676);
  and g21106 (n11677, n_11430, n_11431);
  not g21107 (n_11432, n11602);
  not g21108 (n_11433, n11677);
  and g21109 (n11678, n_11432, n_11433);
  and g21110 (n11679, n11602, n11677);
  not g21111 (n_11434, n11678);
  not g21112 (n_11435, n11679);
  and g21113 (n11680, n_11434, n_11435);
  not g21114 (n_11436, n11600);
  and g21115 (n11681, n_11436, n11680);
  not g21116 (n_11437, n11680);
  and g21117 (n11682, n11600, n_11437);
  not g21118 (n_11438, n11681);
  not g21119 (n_11439, n11682);
  and g21120 (n11683, n_11438, n_11439);
  not g21121 (n_11440, n11520);
  not g21122 (n_11441, n11683);
  and g21123 (n11684, n_11440, n_11441);
  and g21124 (n11685, n11520, n11683);
  not g21125 (n_11442, n11684);
  not g21126 (n_11443, n11685);
  and g21127 (n11686, n_11442, n_11443);
  and g21128 (n11687, n_1880, n_1878);
  not g21129 (n_11444, n11687);
  and g21130 (n11688, n_1879, n_11444);
  and g21131 (n11689, n_1403, n_1401);
  not g21132 (n_11445, n11689);
  and g21133 (n11690, n_1402, n_11445);
  and g21134 (n11691, n_1396, n_1394);
  not g21135 (n_11446, n11691);
  and g21136 (n11692, n_1395, n_11446);
  and g21137 (n11693, n2243, n_1388);
  not g21138 (n_11447, n11693);
  and g21139 (n11694, n_1389, n_11447);
  and g21140 (n11695, n_1301, n_1300);
  not g21141 (n_11448, n11695);
  and g21142 (n11696, n_1299, n_11448);
  and g21143 (n11697, n_1345, n_1344);
  not g21144 (n_11449, n11697);
  and g21145 (n11698, n_1343, n_11449);
  not g21146 (n_11450, n11696);
  and g21147 (n11699, n_11450, n11698);
  not g21148 (n_11451, n11698);
  and g21149 (n11700, n11696, n_11451);
  not g21150 (n_11452, n11699);
  not g21151 (n_11453, n11700);
  and g21152 (n11701, n_11452, n_11453);
  not g21153 (n_11454, n11694);
  not g21154 (n_11455, n11701);
  and g21155 (n11702, n_11454, n_11455);
  not g21159 (n_11456, n11702);
  not g21160 (n_11457, n11705);
  and g21161 (n11706, n_11456, n_11457);
  and g21162 (n11707, n2219, n_1367);
  not g21163 (n_11458, n11707);
  and g21164 (n11708, n_1368, n_11458);
  and g21165 (n11709, n_1209, n_1208);
  not g21166 (n_11459, n11709);
  and g21167 (n11710, n_1207, n_11459);
  and g21168 (n11711, n_1253, n_1252);
  not g21169 (n_11460, n11711);
  and g21170 (n11712, n_1251, n_11460);
  not g21171 (n_11461, n11710);
  and g21172 (n11713, n_11461, n11712);
  not g21173 (n_11462, n11712);
  and g21174 (n11714, n11710, n_11462);
  not g21175 (n_11463, n11713);
  not g21176 (n_11464, n11714);
  and g21177 (n11715, n_11463, n_11464);
  not g21178 (n_11465, n11708);
  not g21179 (n_11466, n11715);
  and g21180 (n11716, n_11465, n_11466);
  not g21184 (n_11467, n11716);
  not g21185 (n_11468, n11719);
  and g21186 (n11720, n_11467, n_11468);
  not g21187 (n_11469, n11706);
  and g21188 (n11721, n_11469, n11720);
  not g21189 (n_11470, n11720);
  and g21190 (n11722, n11706, n_11470);
  not g21191 (n_11471, n11721);
  not g21192 (n_11472, n11722);
  and g21193 (n11723, n_11471, n_11472);
  not g21194 (n_11473, n11692);
  not g21195 (n_11474, n11723);
  and g21196 (n11724, n_11473, n_11474);
  and g21197 (n11725, n11692, n11723);
  not g21198 (n_11475, n11724);
  not g21199 (n_11476, n11725);
  and g21200 (n11726, n_11475, n_11476);
  and g21201 (n11727, n_1160, n_1158);
  not g21202 (n_11477, n11727);
  and g21203 (n11728, n_1159, n_11477);
  and g21204 (n11729, n1892, n_1040);
  not g21205 (n_11478, n11729);
  and g21206 (n11730, n_1041, n_11478);
  and g21207 (n11731, n_1027, n_1030);
  not g21208 (n_11479, n11731);
  and g21209 (n11732, n_1026, n_11479);
  and g21210 (n11733, n_986, n_984);
  not g21211 (n_11480, n11733);
  and g21212 (n11734, n_985, n_11480);
  not g21213 (n_11481, n11732);
  and g21214 (n11735, n_11481, n11734);
  not g21215 (n_11482, n11734);
  and g21216 (n11736, n11732, n_11482);
  not g21217 (n_11483, n11735);
  not g21218 (n_11484, n11736);
  and g21219 (n11737, n_11483, n_11484);
  not g21220 (n_11485, n11730);
  not g21221 (n_11486, n11737);
  and g21222 (n11738, n_11485, n_11486);
  not g21226 (n_11487, n11738);
  not g21227 (n_11488, n11741);
  and g21228 (n11742, n_11487, n_11488);
  and g21229 (n11743, n1981, n_1137);
  not g21230 (n_11489, n11743);
  and g21231 (n11744, n_1138, n_11489);
  and g21232 (n11745, n_1128, n_1131);
  not g21233 (n_11490, n11745);
  and g21234 (n11746, n_1127, n_11490);
  and g21235 (n11747, n_1087, n_1085);
  not g21236 (n_11491, n11747);
  and g21237 (n11748, n_1086, n_11491);
  not g21238 (n_11492, n11746);
  and g21239 (n11749, n_11492, n11748);
  not g21240 (n_11493, n11748);
  and g21241 (n11750, n11746, n_11493);
  not g21242 (n_11494, n11749);
  not g21243 (n_11495, n11750);
  and g21244 (n11751, n_11494, n_11495);
  not g21245 (n_11496, n11744);
  not g21246 (n_11497, n11751);
  and g21247 (n11752, n_11496, n_11497);
  not g21251 (n_11498, n11752);
  not g21252 (n_11499, n11755);
  and g21253 (n11756, n_11498, n_11499);
  not g21254 (n_11500, n11742);
  and g21255 (n11757, n_11500, n11756);
  not g21256 (n_11501, n11756);
  and g21257 (n11758, n11742, n_11501);
  not g21258 (n_11502, n11757);
  not g21259 (n_11503, n11758);
  and g21260 (n11759, n_11502, n_11503);
  not g21261 (n_11504, n11728);
  not g21262 (n_11505, n11759);
  and g21263 (n11760, n_11504, n_11505);
  and g21264 (n11761, n11728, n11759);
  not g21265 (n_11506, n11760);
  not g21266 (n_11507, n11761);
  and g21267 (n11762, n_11506, n_11507);
  not g21268 (n_11508, n11726);
  and g21269 (n11763, n_11508, n11762);
  not g21270 (n_11509, n11762);
  and g21271 (n11764, n11726, n_11509);
  not g21272 (n_11510, n11763);
  not g21273 (n_11511, n11764);
  and g21274 (n11765, n_11510, n_11511);
  not g21275 (n_11512, n11690);
  not g21276 (n_11513, n11765);
  and g21277 (n11766, n_11512, n_11513);
  and g21278 (n11767, n11690, n11765);
  not g21279 (n_11514, n11766);
  not g21280 (n_11515, n11767);
  and g21281 (n11768, n_11514, n_11515);
  and g21282 (n11769, n_1863, n_1861);
  not g21283 (n_11516, n11769);
  and g21284 (n11770, n_1862, n_11516);
  and g21285 (n11771, n_1626, n_1624);
  not g21286 (n_11517, n11771);
  and g21287 (n11772, n_1625, n_11517);
  and g21288 (n11773, n2450, n_1618);
  not g21289 (n_11518, n11773);
  and g21290 (n11774, n_1619, n_11518);
  and g21291 (n11775, n_1552, n_1551);
  not g21292 (n_11519, n11775);
  and g21293 (n11776, n_1550, n_11519);
  and g21294 (n11777, n_1596, n_1595);
  not g21295 (n_11520, n11777);
  and g21296 (n11778, n_1594, n_11520);
  not g21297 (n_11521, n11776);
  and g21298 (n11779, n_11521, n11778);
  not g21299 (n_11522, n11778);
  and g21300 (n11780, n11776, n_11522);
  not g21301 (n_11523, n11779);
  not g21302 (n_11524, n11780);
  and g21303 (n11781, n_11523, n_11524);
  not g21304 (n_11525, n11774);
  not g21305 (n_11526, n11781);
  and g21306 (n11782, n_11525, n_11526);
  not g21310 (n_11527, n11782);
  not g21311 (n_11528, n11785);
  and g21312 (n11786, n_11527, n_11528);
  and g21313 (n11787, n2310, n_1499);
  not g21314 (n_11529, n11787);
  and g21315 (n11788, n_1500, n_11529);
  and g21316 (n11789, n_1490, n_1493);
  not g21317 (n_11530, n11789);
  and g21318 (n11790, n_1489, n_11530);
  and g21319 (n11791, n_1449, n_1447);
  not g21320 (n_11531, n11791);
  and g21321 (n11792, n_1448, n_11531);
  not g21322 (n_11532, n11790);
  and g21323 (n11793, n_11532, n11792);
  not g21324 (n_11533, n11792);
  and g21325 (n11794, n11790, n_11533);
  not g21326 (n_11534, n11793);
  not g21327 (n_11535, n11794);
  and g21328 (n11795, n_11534, n_11535);
  not g21329 (n_11536, n11788);
  not g21330 (n_11537, n11795);
  and g21331 (n11796, n_11536, n_11537);
  not g21335 (n_11538, n11796);
  not g21336 (n_11539, n11799);
  and g21337 (n11800, n_11538, n_11539);
  not g21338 (n_11540, n11786);
  and g21339 (n11801, n_11540, n11800);
  not g21340 (n_11541, n11800);
  and g21341 (n11802, n11786, n_11541);
  not g21342 (n_11542, n11801);
  not g21343 (n_11543, n11802);
  and g21344 (n11803, n_11542, n_11543);
  not g21345 (n_11544, n11772);
  not g21346 (n_11545, n11803);
  and g21347 (n11804, n_11544, n_11545);
  and g21348 (n11805, n11772, n11803);
  not g21349 (n_11546, n11804);
  not g21350 (n_11547, n11805);
  and g21351 (n11806, n_11546, n_11547);
  and g21352 (n11807, n_1846, n_1844);
  not g21353 (n_11548, n11807);
  and g21354 (n11808, n_1845, n_11548);
  and g21355 (n11809, n2510, n_1726);
  not g21356 (n_11549, n11809);
  and g21357 (n11810, n_1727, n_11549);
  and g21358 (n11811, n_1713, n_1716);
  not g21359 (n_11550, n11811);
  and g21360 (n11812, n_1712, n_11550);
  and g21361 (n11813, n_1672, n_1670);
  not g21362 (n_11551, n11813);
  and g21363 (n11814, n_1671, n_11551);
  not g21364 (n_11552, n11812);
  and g21365 (n11815, n_11552, n11814);
  not g21366 (n_11553, n11814);
  and g21367 (n11816, n11812, n_11553);
  not g21368 (n_11554, n11815);
  not g21369 (n_11555, n11816);
  and g21370 (n11817, n_11554, n_11555);
  not g21371 (n_11556, n11810);
  not g21372 (n_11557, n11817);
  and g21373 (n11818, n_11556, n_11557);
  not g21377 (n_11558, n11818);
  not g21378 (n_11559, n11821);
  and g21379 (n11822, n_11558, n_11559);
  and g21380 (n11823, n2599, n_1823);
  not g21381 (n_11560, n11823);
  and g21382 (n11824, n_1824, n_11560);
  and g21383 (n11825, n_1814, n_1817);
  not g21384 (n_11561, n11825);
  and g21385 (n11826, n_1813, n_11561);
  and g21386 (n11827, n_1773, n_1771);
  not g21387 (n_11562, n11827);
  and g21388 (n11828, n_1772, n_11562);
  not g21389 (n_11563, n11826);
  and g21390 (n11829, n_11563, n11828);
  not g21391 (n_11564, n11828);
  and g21392 (n11830, n11826, n_11564);
  not g21393 (n_11565, n11829);
  not g21394 (n_11566, n11830);
  and g21395 (n11831, n_11565, n_11566);
  not g21396 (n_11567, n11824);
  not g21397 (n_11568, n11831);
  and g21398 (n11832, n_11567, n_11568);
  not g21402 (n_11569, n11832);
  not g21403 (n_11570, n11835);
  and g21404 (n11836, n_11569, n_11570);
  not g21405 (n_11571, n11822);
  and g21406 (n11837, n_11571, n11836);
  not g21407 (n_11572, n11836);
  and g21408 (n11838, n11822, n_11572);
  not g21409 (n_11573, n11837);
  not g21410 (n_11574, n11838);
  and g21411 (n11839, n_11573, n_11574);
  not g21412 (n_11575, n11808);
  not g21413 (n_11576, n11839);
  and g21414 (n11840, n_11575, n_11576);
  and g21415 (n11841, n11808, n11839);
  not g21416 (n_11577, n11840);
  not g21417 (n_11578, n11841);
  and g21418 (n11842, n_11577, n_11578);
  not g21419 (n_11579, n11806);
  and g21420 (n11843, n_11579, n11842);
  not g21421 (n_11580, n11842);
  and g21422 (n11844, n11806, n_11580);
  not g21423 (n_11581, n11843);
  not g21424 (n_11582, n11844);
  and g21425 (n11845, n_11581, n_11582);
  not g21426 (n_11583, n11770);
  not g21427 (n_11584, n11845);
  and g21428 (n11846, n_11583, n_11584);
  and g21429 (n11847, n11770, n11845);
  not g21430 (n_11585, n11846);
  not g21431 (n_11586, n11847);
  and g21432 (n11848, n_11585, n_11586);
  not g21433 (n_11587, n11768);
  and g21434 (n11849, n_11587, n11848);
  not g21435 (n_11588, n11848);
  and g21436 (n11850, n11768, n_11588);
  not g21437 (n_11589, n11849);
  not g21438 (n_11590, n11850);
  and g21439 (n11851, n_11589, n_11590);
  not g21440 (n_11591, n11688);
  not g21441 (n_11592, n11851);
  and g21442 (n11852, n_11591, n_11592);
  and g21443 (n11853, n11688, n11851);
  not g21444 (n_11593, n11852);
  not g21445 (n_11594, n11853);
  and g21446 (n11854, n_11593, n_11594);
  not g21447 (n_11595, n11686);
  and g21448 (n11855, n_11595, n11854);
  not g21449 (n_11596, n11854);
  and g21450 (n11856, n11686, n_11596);
  not g21451 (n_11597, n11855);
  not g21452 (n_11598, n11856);
  and g21453 (n11857, n_11597, n_11598);
  not g21454 (n_11599, n11518);
  not g21455 (n_11600, n11857);
  and g21456 (n11858, n_11599, n_11600);
  and g21457 (n11859, n11518, n11857);
  not g21458 (n_11601, n11858);
  not g21459 (n_11602, n11859);
  and g21460 (n11860, n_11601, n_11602);
  not g21461 (n_11603, n11516);
  and g21462 (n11861, n_11603, n11860);
  not g21463 (n_11604, n11860);
  and g21464 (n11862, n11516, n_11604);
  not g21465 (n_11605, n11861);
  not g21466 (n_11606, n11862);
  and g21467 (n11863, n_11605, n_11606);
  not g21468 (n_11607, n11172);
  not g21469 (n_11608, n11863);
  and g21470 (n11864, n_11607, n_11608);
  and g21471 (n11865, n11172, n11863);
  not g21472 (n_11609, n11864);
  not g21473 (n_11610, n11865);
  and g21474 (n11866, n_11609, n_11610);
  not g21475 (n_11611, n11170);
  not g21476 (n_11612, n11866);
  and g21477 (n11867, n_11611, n_11612);
  not g21478 (n_11613, n10047);
  not g21479 (n_11614, n11867);
  and g21480 (n11868, n_11613, n_11614);
  and g21481 (n11869, n_10978, n11866);
  and g21482 (n11870, n_10979, n11869);
  not g21483 (n_11615, n11868);
  not g21484 (n_11616, n11870);
  and g21485 (n11871, n_11615, n_11616);
  and g21486 (n11872, n_10972, n_10973);
  not g21487 (n_11617, n11872);
  and g21488 (n11873, n_10976, n_11617);
  and g21489 (n11874, n10468, n11164);
  not g21490 (n_11618, n11873);
  not g21491 (n_11619, n11874);
  and g21492 (n11875, n_11618, n_11619);
  and g21493 (n11876, n_10964, n_10965);
  not g21494 (n_11620, n11876);
  and g21495 (n11877, n_10968, n_11620);
  and g21496 (n11878, n10814, n11158);
  not g21497 (n_11621, n11877);
  not g21498 (n_11622, n11878);
  and g21499 (n11879, n_11621, n_11622);
  and g21500 (n11880, n_10956, n_10957);
  not g21501 (n_11623, n11880);
  and g21502 (n11881, n_10960, n_11623);
  and g21503 (n11882, n10984, n11152);
  not g21504 (n_11624, n11881);
  not g21505 (n_11625, n11882);
  and g21506 (n11883, n_11624, n_11625);
  and g21507 (n11884, n_10948, n_10949);
  not g21508 (n_11626, n11884);
  and g21509 (n11885, n_10952, n_11626);
  and g21510 (n11886, n11066, n11146);
  not g21511 (n_11627, n11885);
  not g21512 (n_11628, n11886);
  and g21513 (n11887, n_11627, n_11628);
  and g21514 (n11888, n_10940, n_10941);
  not g21515 (n_11629, n11888);
  and g21516 (n11889, n_10944, n_11629);
  and g21517 (n11890, n11104, n11140);
  not g21518 (n_11630, n11889);
  not g21519 (n_11631, n11890);
  and g21520 (n11891, n_11630, n_11631);
  and g21521 (n11892, n_10932, n_10933);
  not g21522 (n_11632, n11892);
  and g21523 (n11893, n_10936, n_11632);
  not g21527 (n_11633, n11893);
  not g21528 (n_11634, n11896);
  and g21529 (n11897, n_11633, n_11634);
  and g21530 (n11898, n_9838, n_10924);
  and g21531 (n11899, n_10921, n11898);
  not g21532 (n_11635, n11899);
  and g21533 (n11900, n11126, n_11635);
  and g21534 (n11901, n_10928, n11124);
  not g21535 (n_11636, n11900);
  not g21536 (n_11637, n11901);
  and g21537 (n11902, n_11636, n_11637);
  and g21538 (n11903, n_9741, n_10913);
  and g21539 (n11904, n_10910, n11903);
  not g21540 (n_11638, n11904);
  and g21541 (n11905, n11112, n_11638);
  and g21542 (n11906, n_10917, n11110);
  not g21543 (n_11639, n11905);
  not g21544 (n_11640, n11906);
  and g21545 (n11907, n_11639, n_11640);
  not g21546 (n_11641, n11902);
  and g21547 (n11908, n_11641, n11907);
  not g21548 (n_11642, n11907);
  and g21549 (n11909, n11902, n_11642);
  not g21550 (n_11643, n11908);
  not g21551 (n_11644, n11909);
  and g21552 (n11910, n_11643, n_11644);
  not g21553 (n_11645, n11897);
  not g21554 (n_11646, n11910);
  and g21555 (n11911, n_11645, n_11646);
  not g21559 (n_11647, n11911);
  not g21560 (n_11648, n11914);
  and g21561 (n11915, n_11647, n_11648);
  and g21562 (n11916, n_10901, n_10902);
  not g21563 (n_11649, n11916);
  and g21564 (n11917, n_10905, n_11649);
  not g21568 (n_11650, n11917);
  not g21569 (n_11651, n11920);
  and g21570 (n11921, n_11650, n_11651);
  and g21571 (n11922, n_9514, n_10893);
  and g21572 (n11923, n_10890, n11922);
  not g21573 (n_11652, n11923);
  and g21574 (n11924, n11090, n_11652);
  and g21575 (n11925, n_10897, n11088);
  not g21576 (n_11653, n11924);
  not g21577 (n_11654, n11925);
  and g21578 (n11926, n_11653, n_11654);
  and g21579 (n11927, n_9633, n_10882);
  and g21580 (n11928, n_10879, n11927);
  not g21581 (n_11655, n11928);
  and g21582 (n11929, n11076, n_11655);
  and g21583 (n11930, n_10886, n11074);
  not g21584 (n_11656, n11929);
  not g21585 (n_11657, n11930);
  and g21586 (n11931, n_11656, n_11657);
  not g21587 (n_11658, n11926);
  and g21588 (n11932, n_11658, n11931);
  not g21589 (n_11659, n11931);
  and g21590 (n11933, n11926, n_11659);
  not g21591 (n_11660, n11932);
  not g21592 (n_11661, n11933);
  and g21593 (n11934, n_11660, n_11661);
  not g21594 (n_11662, n11921);
  not g21595 (n_11663, n11934);
  and g21596 (n11935, n_11662, n_11663);
  not g21600 (n_11664, n11935);
  not g21601 (n_11665, n11938);
  and g21602 (n11939, n_11664, n_11665);
  not g21603 (n_11666, n11915);
  and g21604 (n11940, n_11666, n11939);
  not g21605 (n_11667, n11939);
  and g21606 (n11941, n11915, n_11667);
  not g21607 (n_11668, n11940);
  not g21608 (n_11669, n11941);
  and g21609 (n11942, n_11668, n_11669);
  not g21610 (n_11670, n11891);
  not g21611 (n_11671, n11942);
  and g21612 (n11943, n_11670, n_11671);
  and g21613 (n11944, n11891, n11942);
  not g21614 (n_11672, n11943);
  not g21615 (n_11673, n11944);
  and g21616 (n11945, n_11672, n_11673);
  and g21617 (n11946, n_10869, n_10870);
  not g21618 (n_11674, n11946);
  and g21619 (n11947, n_10873, n_11674);
  and g21620 (n11948, n11024, n11060);
  not g21621 (n_11675, n11947);
  not g21622 (n_11676, n11948);
  and g21623 (n11949, n_11675, n_11676);
  and g21624 (n11950, n_10861, n_10862);
  not g21625 (n_11677, n11950);
  and g21626 (n11951, n_10865, n_11677);
  not g21630 (n_11678, n11951);
  not g21631 (n_11679, n11954);
  and g21632 (n11955, n_11678, n_11679);
  and g21633 (n11956, n_9152, n_10853);
  and g21634 (n11957, n_10850, n11956);
  not g21635 (n_11680, n11957);
  and g21636 (n11958, n11046, n_11680);
  and g21637 (n11959, n_10857, n11044);
  not g21638 (n_11681, n11958);
  not g21639 (n_11682, n11959);
  and g21640 (n11960, n_11681, n_11682);
  and g21641 (n11961, n_9055, n_10842);
  and g21642 (n11962, n_10839, n11961);
  not g21643 (n_11683, n11962);
  and g21644 (n11963, n11032, n_11683);
  and g21645 (n11964, n_10846, n11030);
  not g21646 (n_11684, n11963);
  not g21647 (n_11685, n11964);
  and g21648 (n11965, n_11684, n_11685);
  not g21649 (n_11686, n11960);
  and g21650 (n11966, n_11686, n11965);
  not g21651 (n_11687, n11965);
  and g21652 (n11967, n11960, n_11687);
  not g21653 (n_11688, n11966);
  not g21654 (n_11689, n11967);
  and g21655 (n11968, n_11688, n_11689);
  not g21656 (n_11690, n11955);
  not g21657 (n_11691, n11968);
  and g21658 (n11969, n_11690, n_11691);
  not g21662 (n_11692, n11969);
  not g21663 (n_11693, n11972);
  and g21664 (n11973, n_11692, n_11693);
  and g21665 (n11974, n_10830, n_10831);
  not g21666 (n_11694, n11974);
  and g21667 (n11975, n_10834, n_11694);
  not g21671 (n_11695, n11975);
  not g21672 (n_11696, n11978);
  and g21673 (n11979, n_11695, n_11696);
  and g21674 (n11980, n_9382, n_10822);
  and g21675 (n11981, n_10819, n11980);
  not g21676 (n_11697, n11981);
  and g21677 (n11982, n11010, n_11697);
  and g21678 (n11983, n_10826, n11008);
  not g21679 (n_11698, n11982);
  not g21680 (n_11699, n11983);
  and g21681 (n11984, n_11698, n_11699);
  and g21682 (n11985, n_9403, n_10811);
  and g21683 (n11986, n_10808, n11985);
  not g21684 (n_11700, n11986);
  and g21685 (n11987, n10996, n_11700);
  and g21686 (n11988, n_10815, n10994);
  not g21687 (n_11701, n11987);
  not g21688 (n_11702, n11988);
  and g21689 (n11989, n_11701, n_11702);
  not g21690 (n_11703, n11984);
  and g21691 (n11990, n_11703, n11989);
  not g21692 (n_11704, n11989);
  and g21693 (n11991, n11984, n_11704);
  not g21694 (n_11705, n11990);
  not g21695 (n_11706, n11991);
  and g21696 (n11992, n_11705, n_11706);
  not g21697 (n_11707, n11979);
  not g21698 (n_11708, n11992);
  and g21699 (n11993, n_11707, n_11708);
  not g21703 (n_11709, n11993);
  not g21704 (n_11710, n11996);
  and g21705 (n11997, n_11709, n_11710);
  not g21706 (n_11711, n11973);
  and g21707 (n11998, n_11711, n11997);
  not g21708 (n_11712, n11997);
  and g21709 (n11999, n11973, n_11712);
  not g21710 (n_11713, n11998);
  not g21711 (n_11714, n11999);
  and g21712 (n12000, n_11713, n_11714);
  not g21713 (n_11715, n11949);
  not g21714 (n_11716, n12000);
  and g21715 (n12001, n_11715, n_11716);
  and g21716 (n12002, n11949, n12000);
  not g21717 (n_11717, n12001);
  not g21718 (n_11718, n12002);
  and g21719 (n12003, n_11717, n_11718);
  not g21720 (n_11719, n11945);
  and g21721 (n12004, n_11719, n12003);
  not g21722 (n_11720, n12003);
  and g21723 (n12005, n11945, n_11720);
  not g21724 (n_11721, n12004);
  not g21725 (n_11722, n12005);
  and g21726 (n12006, n_11721, n_11722);
  not g21727 (n_11723, n11887);
  not g21728 (n_11724, n12006);
  and g21729 (n12007, n_11723, n_11724);
  and g21730 (n12008, n11887, n12006);
  not g21731 (n_11725, n12007);
  not g21732 (n_11726, n12008);
  and g21733 (n12009, n_11725, n_11726);
  and g21734 (n12010, n_10797, n_10798);
  not g21735 (n_11727, n12010);
  and g21736 (n12011, n_10801, n_11727);
  and g21737 (n12012, n10898, n10978);
  not g21738 (n_11728, n12011);
  not g21739 (n_11729, n12012);
  and g21740 (n12013, n_11728, n_11729);
  and g21741 (n12014, n_10789, n_10790);
  not g21742 (n_11730, n12014);
  and g21743 (n12015, n_10793, n_11730);
  and g21744 (n12016, n10936, n10972);
  not g21745 (n_11731, n12015);
  not g21746 (n_11732, n12016);
  and g21747 (n12017, n_11731, n_11732);
  and g21748 (n12018, n_10781, n_10782);
  not g21749 (n_11733, n12018);
  and g21750 (n12019, n_10785, n_11733);
  not g21754 (n_11734, n12019);
  not g21755 (n_11735, n12022);
  and g21756 (n12023, n_11734, n_11735);
  and g21757 (n12024, n_8432, n_10773);
  and g21758 (n12025, n_10770, n12024);
  not g21759 (n_11736, n12025);
  and g21760 (n12026, n10958, n_11736);
  and g21761 (n12027, n_10777, n10956);
  not g21762 (n_11737, n12026);
  not g21763 (n_11738, n12027);
  and g21764 (n12028, n_11737, n_11738);
  and g21765 (n12029, n_8335, n_10762);
  and g21766 (n12030, n_10759, n12029);
  not g21767 (n_11739, n12030);
  and g21768 (n12031, n10944, n_11739);
  and g21769 (n12032, n_10766, n10942);
  not g21770 (n_11740, n12031);
  not g21771 (n_11741, n12032);
  and g21772 (n12033, n_11740, n_11741);
  not g21773 (n_11742, n12028);
  and g21774 (n12034, n_11742, n12033);
  not g21775 (n_11743, n12033);
  and g21776 (n12035, n12028, n_11743);
  not g21777 (n_11744, n12034);
  not g21778 (n_11745, n12035);
  and g21779 (n12036, n_11744, n_11745);
  not g21780 (n_11746, n12023);
  not g21781 (n_11747, n12036);
  and g21782 (n12037, n_11746, n_11747);
  not g21786 (n_11748, n12037);
  not g21787 (n_11749, n12040);
  and g21788 (n12041, n_11748, n_11749);
  and g21789 (n12042, n_10750, n_10751);
  not g21790 (n_11750, n12042);
  and g21791 (n12043, n_10754, n_11750);
  not g21795 (n_11751, n12043);
  not g21796 (n_11752, n12046);
  and g21797 (n12047, n_11751, n_11752);
  and g21798 (n12048, n_8108, n_10742);
  and g21799 (n12049, n_10739, n12048);
  not g21800 (n_11753, n12049);
  and g21801 (n12050, n10922, n_11753);
  and g21802 (n12051, n_10746, n10920);
  not g21803 (n_11754, n12050);
  not g21804 (n_11755, n12051);
  and g21805 (n12052, n_11754, n_11755);
  and g21806 (n12053, n_8227, n_10731);
  and g21807 (n12054, n_10728, n12053);
  not g21808 (n_11756, n12054);
  and g21809 (n12055, n10908, n_11756);
  and g21810 (n12056, n_10735, n10906);
  not g21811 (n_11757, n12055);
  not g21812 (n_11758, n12056);
  and g21813 (n12057, n_11757, n_11758);
  not g21814 (n_11759, n12052);
  and g21815 (n12058, n_11759, n12057);
  not g21816 (n_11760, n12057);
  and g21817 (n12059, n12052, n_11760);
  not g21818 (n_11761, n12058);
  not g21819 (n_11762, n12059);
  and g21820 (n12060, n_11761, n_11762);
  not g21821 (n_11763, n12047);
  not g21822 (n_11764, n12060);
  and g21823 (n12061, n_11763, n_11764);
  not g21827 (n_11765, n12061);
  not g21828 (n_11766, n12064);
  and g21829 (n12065, n_11765, n_11766);
  not g21830 (n_11767, n12041);
  and g21831 (n12066, n_11767, n12065);
  not g21832 (n_11768, n12065);
  and g21833 (n12067, n12041, n_11768);
  not g21834 (n_11769, n12066);
  not g21835 (n_11770, n12067);
  and g21836 (n12068, n_11769, n_11770);
  not g21837 (n_11771, n12017);
  not g21838 (n_11772, n12068);
  and g21839 (n12069, n_11771, n_11772);
  and g21840 (n12070, n12017, n12068);
  not g21841 (n_11773, n12069);
  not g21842 (n_11774, n12070);
  and g21843 (n12071, n_11773, n_11774);
  and g21844 (n12072, n_10718, n_10719);
  not g21845 (n_11775, n12072);
  and g21846 (n12073, n_10722, n_11775);
  and g21847 (n12074, n10856, n10892);
  not g21848 (n_11776, n12073);
  not g21849 (n_11777, n12074);
  and g21850 (n12075, n_11776, n_11777);
  and g21851 (n12076, n_10710, n_10711);
  not g21852 (n_11778, n12076);
  and g21853 (n12077, n_10714, n_11778);
  not g21857 (n_11779, n12077);
  not g21858 (n_11780, n12080);
  and g21859 (n12081, n_11779, n_11780);
  and g21860 (n12082, n_8884, n_10702);
  and g21861 (n12083, n_10699, n12082);
  not g21862 (n_11781, n12083);
  and g21863 (n12084, n10878, n_11781);
  and g21864 (n12085, n_10706, n10876);
  not g21865 (n_11782, n12084);
  not g21866 (n_11783, n12085);
  and g21867 (n12086, n_11782, n_11783);
  and g21868 (n12087, n_8875, n_10691);
  and g21869 (n12088, n_10688, n12087);
  not g21870 (n_11784, n12088);
  and g21871 (n12089, n10864, n_11784);
  and g21872 (n12090, n_10695, n10862);
  not g21873 (n_11785, n12089);
  not g21874 (n_11786, n12090);
  and g21875 (n12091, n_11785, n_11786);
  not g21876 (n_11787, n12086);
  and g21877 (n12092, n_11787, n12091);
  not g21878 (n_11788, n12091);
  and g21879 (n12093, n12086, n_11788);
  not g21880 (n_11789, n12092);
  not g21881 (n_11790, n12093);
  and g21882 (n12094, n_11789, n_11790);
  not g21883 (n_11791, n12081);
  not g21884 (n_11792, n12094);
  and g21885 (n12095, n_11791, n_11792);
  not g21889 (n_11793, n12095);
  not g21890 (n_11794, n12098);
  and g21891 (n12099, n_11793, n_11794);
  and g21892 (n12100, n_10679, n_10680);
  not g21893 (n_11795, n12100);
  and g21894 (n12101, n_10683, n_11795);
  not g21898 (n_11796, n12101);
  not g21899 (n_11797, n12104);
  and g21900 (n12105, n_11796, n_11797);
  and g21901 (n12106, n_8912, n_10671);
  and g21902 (n12107, n_10668, n12106);
  not g21903 (n_11798, n12107);
  and g21904 (n12108, n10842, n_11798);
  and g21905 (n12109, n_10675, n10840);
  not g21906 (n_11799, n12108);
  not g21907 (n_11800, n12109);
  and g21908 (n12110, n_11799, n_11800);
  and g21909 (n12111, n_8933, n_10660);
  and g21910 (n12112, n_10657, n12111);
  not g21911 (n_11801, n12112);
  and g21912 (n12113, n10828, n_11801);
  and g21913 (n12114, n_10664, n10826);
  not g21914 (n_11802, n12113);
  not g21915 (n_11803, n12114);
  and g21916 (n12115, n_11802, n_11803);
  not g21917 (n_11804, n12110);
  and g21918 (n12116, n_11804, n12115);
  not g21919 (n_11805, n12115);
  and g21920 (n12117, n12110, n_11805);
  not g21921 (n_11806, n12116);
  not g21922 (n_11807, n12117);
  and g21923 (n12118, n_11806, n_11807);
  not g21924 (n_11808, n12105);
  not g21925 (n_11809, n12118);
  and g21926 (n12119, n_11808, n_11809);
  not g21930 (n_11810, n12119);
  not g21931 (n_11811, n12122);
  and g21932 (n12123, n_11810, n_11811);
  not g21933 (n_11812, n12099);
  and g21934 (n12124, n_11812, n12123);
  not g21935 (n_11813, n12123);
  and g21936 (n12125, n12099, n_11813);
  not g21937 (n_11814, n12124);
  not g21938 (n_11815, n12125);
  and g21939 (n12126, n_11814, n_11815);
  not g21940 (n_11816, n12075);
  not g21941 (n_11817, n12126);
  and g21942 (n12127, n_11816, n_11817);
  and g21943 (n12128, n12075, n12126);
  not g21944 (n_11818, n12127);
  not g21945 (n_11819, n12128);
  and g21946 (n12129, n_11818, n_11819);
  not g21947 (n_11820, n12071);
  and g21948 (n12130, n_11820, n12129);
  not g21949 (n_11821, n12129);
  and g21950 (n12131, n12071, n_11821);
  not g21951 (n_11822, n12130);
  not g21952 (n_11823, n12131);
  and g21953 (n12132, n_11822, n_11823);
  not g21954 (n_11824, n12013);
  not g21955 (n_11825, n12132);
  and g21956 (n12133, n_11824, n_11825);
  and g21957 (n12134, n12013, n12132);
  not g21958 (n_11826, n12133);
  not g21959 (n_11827, n12134);
  and g21960 (n12135, n_11826, n_11827);
  not g21961 (n_11828, n12009);
  and g21962 (n12136, n_11828, n12135);
  not g21963 (n_11829, n12135);
  and g21964 (n12137, n12009, n_11829);
  not g21965 (n_11830, n12136);
  not g21966 (n_11831, n12137);
  and g21967 (n12138, n_11830, n_11831);
  not g21968 (n_11832, n11883);
  not g21969 (n_11833, n12138);
  and g21970 (n12139, n_11832, n_11833);
  and g21971 (n12140, n11883, n12138);
  not g21972 (n_11834, n12139);
  not g21973 (n_11835, n12140);
  and g21974 (n12141, n_11834, n_11835);
  and g21975 (n12142, n_10645, n_10646);
  not g21976 (n_11836, n12142);
  and g21977 (n12143, n_10649, n_11836);
  and g21978 (n12144, n10640, n10808);
  not g21979 (n_11837, n12143);
  not g21980 (n_11838, n12144);
  and g21981 (n12145, n_11837, n_11838);
  and g21982 (n12146, n_10637, n_10638);
  not g21983 (n_11839, n12146);
  and g21984 (n12147, n_10641, n_11839);
  and g21985 (n12148, n10722, n10802);
  not g21986 (n_11840, n12147);
  not g21987 (n_11841, n12148);
  and g21988 (n12149, n_11840, n_11841);
  and g21989 (n12150, n_10629, n_10630);
  not g21990 (n_11842, n12150);
  and g21991 (n12151, n_10633, n_11842);
  and g21992 (n12152, n10760, n10796);
  not g21993 (n_11843, n12151);
  not g21994 (n_11844, n12152);
  and g21995 (n12153, n_11843, n_11844);
  and g21996 (n12154, n_10621, n_10622);
  not g21997 (n_11845, n12154);
  and g21998 (n12155, n_10625, n_11845);
  not g22002 (n_11846, n12155);
  not g22003 (n_11847, n12158);
  and g22004 (n12159, n_11846, n_11847);
  and g22005 (n12160, n_6992, n_10613);
  and g22006 (n12161, n_10610, n12160);
  not g22007 (n_11848, n12161);
  and g22008 (n12162, n10782, n_11848);
  and g22009 (n12163, n_10617, n10780);
  not g22010 (n_11849, n12162);
  not g22011 (n_11850, n12163);
  and g22012 (n12164, n_11849, n_11850);
  and g22013 (n12165, n_6895, n_10602);
  and g22014 (n12166, n_10599, n12165);
  not g22015 (n_11851, n12166);
  and g22016 (n12167, n10768, n_11851);
  and g22017 (n12168, n_10606, n10766);
  not g22018 (n_11852, n12167);
  not g22019 (n_11853, n12168);
  and g22020 (n12169, n_11852, n_11853);
  not g22021 (n_11854, n12164);
  and g22022 (n12170, n_11854, n12169);
  not g22023 (n_11855, n12169);
  and g22024 (n12171, n12164, n_11855);
  not g22025 (n_11856, n12170);
  not g22026 (n_11857, n12171);
  and g22027 (n12172, n_11856, n_11857);
  not g22028 (n_11858, n12159);
  not g22029 (n_11859, n12172);
  and g22030 (n12173, n_11858, n_11859);
  not g22034 (n_11860, n12173);
  not g22035 (n_11861, n12176);
  and g22036 (n12177, n_11860, n_11861);
  and g22037 (n12178, n_10590, n_10591);
  not g22038 (n_11862, n12178);
  and g22039 (n12179, n_10594, n_11862);
  not g22043 (n_11863, n12179);
  not g22044 (n_11864, n12182);
  and g22045 (n12183, n_11863, n_11864);
  and g22046 (n12184, n_6668, n_10582);
  and g22047 (n12185, n_10579, n12184);
  not g22048 (n_11865, n12185);
  and g22049 (n12186, n10746, n_11865);
  and g22050 (n12187, n_10586, n10744);
  not g22051 (n_11866, n12186);
  not g22052 (n_11867, n12187);
  and g22053 (n12188, n_11866, n_11867);
  and g22054 (n12189, n_6787, n_10571);
  and g22055 (n12190, n_10568, n12189);
  not g22056 (n_11868, n12190);
  and g22057 (n12191, n10732, n_11868);
  and g22058 (n12192, n_10575, n10730);
  not g22059 (n_11869, n12191);
  not g22060 (n_11870, n12192);
  and g22061 (n12193, n_11869, n_11870);
  not g22062 (n_11871, n12188);
  and g22063 (n12194, n_11871, n12193);
  not g22064 (n_11872, n12193);
  and g22065 (n12195, n12188, n_11872);
  not g22066 (n_11873, n12194);
  not g22067 (n_11874, n12195);
  and g22068 (n12196, n_11873, n_11874);
  not g22069 (n_11875, n12183);
  not g22070 (n_11876, n12196);
  and g22071 (n12197, n_11875, n_11876);
  not g22075 (n_11877, n12197);
  not g22076 (n_11878, n12200);
  and g22077 (n12201, n_11877, n_11878);
  not g22078 (n_11879, n12177);
  and g22079 (n12202, n_11879, n12201);
  not g22080 (n_11880, n12201);
  and g22081 (n12203, n12177, n_11880);
  not g22082 (n_11881, n12202);
  not g22083 (n_11882, n12203);
  and g22084 (n12204, n_11881, n_11882);
  not g22085 (n_11883, n12153);
  not g22086 (n_11884, n12204);
  and g22087 (n12205, n_11883, n_11884);
  and g22088 (n12206, n12153, n12204);
  not g22089 (n_11885, n12205);
  not g22090 (n_11886, n12206);
  and g22091 (n12207, n_11885, n_11886);
  and g22092 (n12208, n_10558, n_10559);
  not g22093 (n_11887, n12208);
  and g22094 (n12209, n_10562, n_11887);
  and g22095 (n12210, n10680, n10716);
  not g22096 (n_11888, n12209);
  not g22097 (n_11889, n12210);
  and g22098 (n12211, n_11888, n_11889);
  and g22099 (n12212, n_10550, n_10551);
  not g22100 (n_11890, n12212);
  and g22101 (n12213, n_10554, n_11890);
  not g22105 (n_11891, n12213);
  not g22106 (n_11892, n12216);
  and g22107 (n12217, n_11891, n_11892);
  and g22108 (n12218, n_6306, n_10542);
  and g22109 (n12219, n_10539, n12218);
  not g22110 (n_11893, n12219);
  and g22111 (n12220, n10702, n_11893);
  and g22112 (n12221, n_10546, n10700);
  not g22113 (n_11894, n12220);
  not g22114 (n_11895, n12221);
  and g22115 (n12222, n_11894, n_11895);
  and g22116 (n12223, n_6209, n_10531);
  and g22117 (n12224, n_10528, n12223);
  not g22118 (n_11896, n12224);
  and g22119 (n12225, n10688, n_11896);
  and g22120 (n12226, n_10535, n10686);
  not g22121 (n_11897, n12225);
  not g22122 (n_11898, n12226);
  and g22123 (n12227, n_11897, n_11898);
  not g22124 (n_11899, n12222);
  and g22125 (n12228, n_11899, n12227);
  not g22126 (n_11900, n12227);
  and g22127 (n12229, n12222, n_11900);
  not g22128 (n_11901, n12228);
  not g22129 (n_11902, n12229);
  and g22130 (n12230, n_11901, n_11902);
  not g22131 (n_11903, n12217);
  not g22132 (n_11904, n12230);
  and g22133 (n12231, n_11903, n_11904);
  not g22137 (n_11905, n12231);
  not g22138 (n_11906, n12234);
  and g22139 (n12235, n_11905, n_11906);
  and g22140 (n12236, n_10519, n_10520);
  not g22141 (n_11907, n12236);
  and g22142 (n12237, n_10523, n_11907);
  not g22146 (n_11908, n12237);
  not g22147 (n_11909, n12240);
  and g22148 (n12241, n_11908, n_11909);
  and g22149 (n12242, n_6536, n_10511);
  and g22150 (n12243, n_10508, n12242);
  not g22151 (n_11910, n12243);
  and g22152 (n12244, n10666, n_11910);
  and g22153 (n12245, n_10515, n10664);
  not g22154 (n_11911, n12244);
  not g22155 (n_11912, n12245);
  and g22156 (n12246, n_11911, n_11912);
  and g22157 (n12247, n_6557, n_10500);
  and g22158 (n12248, n_10497, n12247);
  not g22159 (n_11913, n12248);
  and g22160 (n12249, n10652, n_11913);
  and g22161 (n12250, n_10504, n10650);
  not g22162 (n_11914, n12249);
  not g22163 (n_11915, n12250);
  and g22164 (n12251, n_11914, n_11915);
  not g22165 (n_11916, n12246);
  and g22166 (n12252, n_11916, n12251);
  not g22167 (n_11917, n12251);
  and g22168 (n12253, n12246, n_11917);
  not g22169 (n_11918, n12252);
  not g22170 (n_11919, n12253);
  and g22171 (n12254, n_11918, n_11919);
  not g22172 (n_11920, n12241);
  not g22173 (n_11921, n12254);
  and g22174 (n12255, n_11920, n_11921);
  not g22178 (n_11922, n12255);
  not g22179 (n_11923, n12258);
  and g22180 (n12259, n_11922, n_11923);
  not g22181 (n_11924, n12235);
  and g22182 (n12260, n_11924, n12259);
  not g22183 (n_11925, n12259);
  and g22184 (n12261, n12235, n_11925);
  not g22185 (n_11926, n12260);
  not g22186 (n_11927, n12261);
  and g22187 (n12262, n_11926, n_11927);
  not g22188 (n_11928, n12211);
  not g22189 (n_11929, n12262);
  and g22190 (n12263, n_11928, n_11929);
  and g22191 (n12264, n12211, n12262);
  not g22192 (n_11930, n12263);
  not g22193 (n_11931, n12264);
  and g22194 (n12265, n_11930, n_11931);
  not g22195 (n_11932, n12207);
  and g22196 (n12266, n_11932, n12265);
  not g22197 (n_11933, n12265);
  and g22198 (n12267, n12207, n_11933);
  not g22199 (n_11934, n12266);
  not g22200 (n_11935, n12267);
  and g22201 (n12268, n_11934, n_11935);
  not g22202 (n_11936, n12149);
  not g22203 (n_11937, n12268);
  and g22204 (n12269, n_11936, n_11937);
  and g22205 (n12270, n12149, n12268);
  not g22206 (n_11938, n12269);
  not g22207 (n_11939, n12270);
  and g22208 (n12271, n_11938, n_11939);
  and g22209 (n12272, n_10486, n_10487);
  not g22210 (n_11940, n12272);
  and g22211 (n12273, n_10490, n_11940);
  and g22212 (n12274, n10554, n10634);
  not g22213 (n_11941, n12273);
  not g22214 (n_11942, n12274);
  and g22215 (n12275, n_11941, n_11942);
  and g22216 (n12276, n_10478, n_10479);
  not g22217 (n_11943, n12276);
  and g22218 (n12277, n_10482, n_11943);
  and g22219 (n12278, n10592, n10628);
  not g22220 (n_11944, n12277);
  not g22221 (n_11945, n12278);
  and g22222 (n12279, n_11944, n_11945);
  and g22223 (n12280, n_10470, n_10471);
  not g22224 (n_11946, n12280);
  and g22225 (n12281, n_10474, n_11946);
  not g22229 (n_11947, n12281);
  not g22230 (n_11948, n12284);
  and g22231 (n12285, n_11947, n_11948);
  and g22232 (n12286, n_7882, n_10462);
  and g22233 (n12287, n_10459, n12286);
  not g22234 (n_11949, n12287);
  and g22235 (n12288, n10614, n_11949);
  and g22236 (n12289, n_10466, n10612);
  not g22237 (n_11950, n12288);
  not g22238 (n_11951, n12289);
  and g22239 (n12290, n_11950, n_11951);
  and g22240 (n12291, n_7873, n_10451);
  and g22241 (n12292, n_10448, n12291);
  not g22242 (n_11952, n12292);
  and g22243 (n12293, n10600, n_11952);
  and g22244 (n12294, n_10455, n10598);
  not g22245 (n_11953, n12293);
  not g22246 (n_11954, n12294);
  and g22247 (n12295, n_11953, n_11954);
  not g22248 (n_11955, n12290);
  and g22249 (n12296, n_11955, n12295);
  not g22250 (n_11956, n12295);
  and g22251 (n12297, n12290, n_11956);
  not g22252 (n_11957, n12296);
  not g22253 (n_11958, n12297);
  and g22254 (n12298, n_11957, n_11958);
  not g22255 (n_11959, n12285);
  not g22256 (n_11960, n12298);
  and g22257 (n12299, n_11959, n_11960);
  not g22261 (n_11961, n12299);
  not g22262 (n_11962, n12302);
  and g22263 (n12303, n_11961, n_11962);
  and g22264 (n12304, n_10439, n_10440);
  not g22265 (n_11963, n12304);
  and g22266 (n12305, n_10443, n_11963);
  not g22270 (n_11964, n12305);
  not g22271 (n_11965, n12308);
  and g22272 (n12309, n_11964, n_11965);
  and g22273 (n12310, n_7832, n_10431);
  and g22274 (n12311, n_10428, n12310);
  not g22275 (n_11966, n12311);
  and g22276 (n12312, n10578, n_11966);
  and g22277 (n12313, n_10435, n10576);
  not g22278 (n_11967, n12312);
  not g22279 (n_11968, n12313);
  and g22280 (n12314, n_11967, n_11968);
  and g22281 (n12315, n_7853, n_10420);
  and g22282 (n12316, n_10417, n12315);
  not g22283 (n_11969, n12316);
  and g22284 (n12317, n10564, n_11969);
  and g22285 (n12318, n_10424, n10562);
  not g22286 (n_11970, n12317);
  not g22287 (n_11971, n12318);
  and g22288 (n12319, n_11970, n_11971);
  not g22289 (n_11972, n12314);
  and g22290 (n12320, n_11972, n12319);
  not g22291 (n_11973, n12319);
  and g22292 (n12321, n12314, n_11973);
  not g22293 (n_11974, n12320);
  not g22294 (n_11975, n12321);
  and g22295 (n12322, n_11974, n_11975);
  not g22296 (n_11976, n12309);
  not g22297 (n_11977, n12322);
  and g22298 (n12323, n_11976, n_11977);
  not g22302 (n_11978, n12323);
  not g22303 (n_11979, n12326);
  and g22304 (n12327, n_11978, n_11979);
  not g22305 (n_11980, n12303);
  and g22306 (n12328, n_11980, n12327);
  not g22307 (n_11981, n12327);
  and g22308 (n12329, n12303, n_11981);
  not g22309 (n_11982, n12328);
  not g22310 (n_11983, n12329);
  and g22311 (n12330, n_11982, n_11983);
  not g22312 (n_11984, n12279);
  not g22313 (n_11985, n12330);
  and g22314 (n12331, n_11984, n_11985);
  and g22315 (n12332, n12279, n12330);
  not g22316 (n_11986, n12331);
  not g22317 (n_11987, n12332);
  and g22318 (n12333, n_11986, n_11987);
  and g22319 (n12334, n_10407, n_10408);
  not g22320 (n_11988, n12334);
  and g22321 (n12335, n_10411, n_11988);
  and g22322 (n12336, n10512, n10548);
  not g22323 (n_11989, n12335);
  not g22324 (n_11990, n12336);
  and g22325 (n12337, n_11989, n_11990);
  and g22326 (n12338, n_10399, n_10400);
  not g22327 (n_11991, n12338);
  and g22328 (n12339, n_10403, n_11991);
  not g22332 (n_11992, n12339);
  not g22333 (n_11993, n12342);
  and g22334 (n12343, n_11992, n_11993);
  and g22335 (n12344, n_7934, n_10391);
  and g22336 (n12345, n_10388, n12344);
  not g22337 (n_11994, n12345);
  and g22338 (n12346, n10534, n_11994);
  and g22339 (n12347, n_10395, n10532);
  not g22340 (n_11995, n12346);
  not g22341 (n_11996, n12347);
  and g22342 (n12348, n_11995, n_11996);
  and g22343 (n12349, n_7925, n_10380);
  and g22344 (n12350, n_10377, n12349);
  not g22345 (n_11997, n12350);
  and g22346 (n12351, n10520, n_11997);
  and g22347 (n12352, n_10384, n10518);
  not g22348 (n_11998, n12351);
  not g22349 (n_11999, n12352);
  and g22350 (n12353, n_11998, n_11999);
  not g22351 (n_12000, n12348);
  and g22352 (n12354, n_12000, n12353);
  not g22353 (n_12001, n12353);
  and g22354 (n12355, n12348, n_12001);
  not g22355 (n_12002, n12354);
  not g22356 (n_12003, n12355);
  and g22357 (n12356, n_12002, n_12003);
  not g22358 (n_12004, n12343);
  not g22359 (n_12005, n12356);
  and g22360 (n12357, n_12004, n_12005);
  not g22364 (n_12006, n12357);
  not g22365 (n_12007, n12360);
  and g22366 (n12361, n_12006, n_12007);
  and g22367 (n12362, n_10368, n_10369);
  not g22368 (n_12008, n12362);
  and g22369 (n12363, n_10372, n_12008);
  not g22373 (n_12009, n12363);
  not g22374 (n_12010, n12366);
  and g22375 (n12367, n_12009, n_12010);
  and g22376 (n12368, n_7962, n_10360);
  and g22377 (n12369, n_10357, n12368);
  not g22378 (n_12011, n12369);
  and g22379 (n12370, n10498, n_12011);
  and g22380 (n12371, n_10364, n10496);
  not g22381 (n_12012, n12370);
  not g22382 (n_12013, n12371);
  and g22383 (n12372, n_12012, n_12013);
  and g22384 (n12373, n_7983, n_10349);
  and g22385 (n12374, n_10346, n12373);
  not g22386 (n_12014, n12374);
  and g22387 (n12375, n10484, n_12014);
  and g22388 (n12376, n_10353, n10482);
  not g22389 (n_12015, n12375);
  not g22390 (n_12016, n12376);
  and g22391 (n12377, n_12015, n_12016);
  not g22392 (n_12017, n12372);
  and g22393 (n12378, n_12017, n12377);
  not g22394 (n_12018, n12377);
  and g22395 (n12379, n12372, n_12018);
  not g22396 (n_12019, n12378);
  not g22397 (n_12020, n12379);
  and g22398 (n12380, n_12019, n_12020);
  not g22399 (n_12021, n12367);
  not g22400 (n_12022, n12380);
  and g22401 (n12381, n_12021, n_12022);
  not g22405 (n_12023, n12381);
  not g22406 (n_12024, n12384);
  and g22407 (n12385, n_12023, n_12024);
  not g22408 (n_12025, n12361);
  and g22409 (n12386, n_12025, n12385);
  not g22410 (n_12026, n12385);
  and g22411 (n12387, n12361, n_12026);
  not g22412 (n_12027, n12386);
  not g22413 (n_12028, n12387);
  and g22414 (n12388, n_12027, n_12028);
  not g22415 (n_12029, n12337);
  not g22416 (n_12030, n12388);
  and g22417 (n12389, n_12029, n_12030);
  and g22418 (n12390, n12337, n12388);
  not g22419 (n_12031, n12389);
  not g22420 (n_12032, n12390);
  and g22421 (n12391, n_12031, n_12032);
  not g22422 (n_12033, n12333);
  and g22423 (n12392, n_12033, n12391);
  not g22424 (n_12034, n12391);
  and g22425 (n12393, n12333, n_12034);
  not g22426 (n_12035, n12392);
  not g22427 (n_12036, n12393);
  and g22428 (n12394, n_12035, n_12036);
  not g22429 (n_12037, n12275);
  not g22430 (n_12038, n12394);
  and g22431 (n12395, n_12037, n_12038);
  and g22432 (n12396, n12275, n12394);
  not g22433 (n_12039, n12395);
  not g22434 (n_12040, n12396);
  and g22435 (n12397, n_12039, n_12040);
  not g22436 (n_12041, n12271);
  and g22437 (n12398, n_12041, n12397);
  not g22438 (n_12042, n12397);
  and g22439 (n12399, n12271, n_12042);
  not g22440 (n_12043, n12398);
  not g22441 (n_12044, n12399);
  and g22442 (n12400, n_12043, n_12044);
  not g22443 (n_12045, n12145);
  not g22444 (n_12046, n12400);
  and g22445 (n12401, n_12045, n_12046);
  and g22446 (n12402, n12145, n12400);
  not g22447 (n_12047, n12401);
  not g22448 (n_12048, n12402);
  and g22449 (n12403, n_12047, n_12048);
  not g22450 (n_12049, n12141);
  and g22451 (n12404, n_12049, n12403);
  not g22452 (n_12050, n12403);
  and g22453 (n12405, n12141, n_12050);
  not g22454 (n_12051, n12404);
  not g22455 (n_12052, n12405);
  and g22456 (n12406, n_12051, n_12052);
  not g22457 (n_12053, n11879);
  not g22458 (n_12054, n12406);
  and g22459 (n12407, n_12053, n_12054);
  and g22460 (n12408, n11879, n12406);
  not g22461 (n_12055, n12407);
  not g22462 (n_12056, n12408);
  and g22463 (n12409, n_12055, n_12056);
  and g22464 (n12410, n_10332, n_10334);
  not g22465 (n_12057, n12410);
  and g22466 (n12411, n_10337, n_12057);
  and g22467 (n12412, n_10331, n10460);
  and g22468 (n12413, n_10333, n12412);
  not g22469 (n_12058, n12411);
  not g22470 (n_12059, n12413);
  and g22471 (n12414, n_12058, n_12059);
  and g22472 (n12415, n_10173, n_10175);
  not g22473 (n_12060, n12415);
  and g22474 (n12416, n_10178, n_12060);
  and g22475 (n12417, n_10172, n10285);
  and g22476 (n12418, n_10174, n12417);
  not g22477 (n_12061, n12416);
  not g22478 (n_12062, n12418);
  and g22479 (n12419, n_12061, n_12062);
  and g22480 (n12420, n_10095, n_10096);
  not g22481 (n_12063, n12420);
  and g22482 (n12421, n_10099, n_12063);
  and g22483 (n12422, n10120, n10200);
  not g22484 (n_12064, n12421);
  not g22485 (n_12065, n12422);
  and g22486 (n12423, n_12064, n_12065);
  and g22487 (n12424, n_10087, n_10088);
  not g22488 (n_12066, n12424);
  and g22489 (n12425, n_10091, n_12066);
  and g22490 (n12426, n10158, n10194);
  not g22491 (n_12067, n12425);
  not g22492 (n_12068, n12426);
  and g22493 (n12427, n_12067, n_12068);
  and g22494 (n12428, n_10079, n_10080);
  not g22495 (n_12069, n12428);
  and g22496 (n12429, n_10083, n_12069);
  not g22500 (n_12070, n12429);
  not g22501 (n_12071, n12432);
  and g22502 (n12433, n_12070, n_12071);
  and g22503 (n12434, n_5072, n_10071);
  and g22504 (n12435, n_10068, n12434);
  not g22505 (n_12072, n12435);
  and g22506 (n12436, n10180, n_12072);
  and g22507 (n12437, n_10075, n10178);
  not g22508 (n_12073, n12436);
  not g22509 (n_12074, n12437);
  and g22510 (n12438, n_12073, n_12074);
  and g22511 (n12439, n_4975, n_10060);
  and g22512 (n12440, n_10057, n12439);
  not g22513 (n_12075, n12440);
  and g22514 (n12441, n10166, n_12075);
  and g22515 (n12442, n_10064, n10164);
  not g22516 (n_12076, n12441);
  not g22517 (n_12077, n12442);
  and g22518 (n12443, n_12076, n_12077);
  not g22519 (n_12078, n12438);
  and g22520 (n12444, n_12078, n12443);
  not g22521 (n_12079, n12443);
  and g22522 (n12445, n12438, n_12079);
  not g22523 (n_12080, n12444);
  not g22524 (n_12081, n12445);
  and g22525 (n12446, n_12080, n_12081);
  not g22526 (n_12082, n12433);
  not g22527 (n_12083, n12446);
  and g22528 (n12447, n_12082, n_12083);
  not g22532 (n_12084, n12447);
  not g22533 (n_12085, n12450);
  and g22534 (n12451, n_12084, n_12085);
  and g22535 (n12452, n_10048, n_10049);
  not g22536 (n_12086, n12452);
  and g22537 (n12453, n_10052, n_12086);
  not g22541 (n_12087, n12453);
  not g22542 (n_12088, n12456);
  and g22543 (n12457, n_12087, n_12088);
  and g22544 (n12458, n_4748, n_10040);
  and g22545 (n12459, n_10037, n12458);
  not g22546 (n_12089, n12459);
  and g22547 (n12460, n10144, n_12089);
  and g22548 (n12461, n_10044, n10142);
  not g22549 (n_12090, n12460);
  not g22550 (n_12091, n12461);
  and g22551 (n12462, n_12090, n_12091);
  and g22552 (n12463, n_4867, n_10029);
  and g22553 (n12464, n_10026, n12463);
  not g22554 (n_12092, n12464);
  and g22555 (n12465, n10130, n_12092);
  and g22556 (n12466, n_10033, n10128);
  not g22557 (n_12093, n12465);
  not g22558 (n_12094, n12466);
  and g22559 (n12467, n_12093, n_12094);
  not g22560 (n_12095, n12462);
  and g22561 (n12468, n_12095, n12467);
  not g22562 (n_12096, n12467);
  and g22563 (n12469, n12462, n_12096);
  not g22564 (n_12097, n12468);
  not g22565 (n_12098, n12469);
  and g22566 (n12470, n_12097, n_12098);
  not g22567 (n_12099, n12457);
  not g22568 (n_12100, n12470);
  and g22569 (n12471, n_12099, n_12100);
  not g22573 (n_12101, n12471);
  not g22574 (n_12102, n12474);
  and g22575 (n12475, n_12101, n_12102);
  not g22576 (n_12103, n12451);
  and g22577 (n12476, n_12103, n12475);
  not g22578 (n_12104, n12475);
  and g22579 (n12477, n12451, n_12104);
  not g22580 (n_12105, n12476);
  not g22581 (n_12106, n12477);
  and g22582 (n12478, n_12105, n_12106);
  not g22583 (n_12107, n12427);
  not g22584 (n_12108, n12478);
  and g22585 (n12479, n_12107, n_12108);
  and g22586 (n12480, n12427, n12478);
  not g22587 (n_12109, n12479);
  not g22588 (n_12110, n12480);
  and g22589 (n12481, n_12109, n_12110);
  and g22590 (n12482, n_10016, n_10017);
  not g22591 (n_12111, n12482);
  and g22592 (n12483, n_10020, n_12111);
  and g22593 (n12484, n10078, n_10014);
  and g22594 (n12485, n_10015, n12484);
  not g22595 (n_12112, n12483);
  not g22596 (n_12113, n12485);
  and g22597 (n12486, n_12112, n_12113);
  and g22598 (n12487, n_4644, n10071);
  and g22599 (n12488, n_9969, n12487);
  not g22600 (n_12114, n12488);
  and g22601 (n12489, n10068, n_12114);
  and g22602 (n12490, n_9981, n_9978);
  not g22603 (n_12115, n12489);
  not g22604 (n_12116, n12490);
  and g22605 (n12491, n_12115, n_12116);
  and g22606 (n12492, n_9972, n_9973);
  not g22607 (n_12117, n12491);
  and g22608 (n12493, n_12117, n12492);
  not g22609 (n_12118, n12492);
  and g22610 (n12494, n_12115, n_12118);
  and g22611 (n12495, n_12116, n12494);
  not g22612 (n_12119, n12493);
  not g22613 (n_12120, n12495);
  and g22614 (n12496, n_12119, n_12120);
  and g22615 (n12497, n_10008, n_10009);
  not g22616 (n_12121, n12497);
  and g22617 (n12498, n_10012, n_12121);
  not g22621 (n_12122, n12498);
  not g22622 (n_12123, n12501);
  and g22623 (n12502, n_12122, n_12123);
  and g22624 (n12503, n_4481, n_10000);
  and g22625 (n12504, n_9997, n12503);
  not g22626 (n_12124, n12504);
  and g22627 (n12505, n10100, n_12124);
  and g22628 (n12506, n_10004, n10098);
  not g22629 (n_12125, n12505);
  not g22630 (n_12126, n12506);
  and g22631 (n12507, n_12125, n_12126);
  and g22632 (n12508, n_4384, n_9989);
  and g22633 (n12509, n_9986, n12508);
  not g22634 (n_12127, n12509);
  and g22635 (n12510, n10086, n_12127);
  and g22636 (n12511, n_9993, n10084);
  not g22637 (n_12128, n12510);
  not g22638 (n_12129, n12511);
  and g22639 (n12512, n_12128, n_12129);
  not g22640 (n_12130, n12507);
  and g22641 (n12513, n_12130, n12512);
  not g22642 (n_12131, n12512);
  and g22643 (n12514, n12507, n_12131);
  not g22644 (n_12132, n12513);
  not g22645 (n_12133, n12514);
  and g22646 (n12515, n_12132, n_12133);
  not g22647 (n_12134, n12502);
  not g22648 (n_12135, n12515);
  and g22649 (n12516, n_12134, n_12135);
  not g22653 (n_12136, n12516);
  not g22654 (n_12137, n12519);
  and g22655 (n12520, n_12136, n_12137);
  not g22656 (n_12138, n12496);
  not g22657 (n_12139, n12520);
  and g22658 (n12521, n_12138, n_12139);
  and g22659 (n12522, n12496, n12520);
  not g22660 (n_12140, n12521);
  not g22661 (n_12141, n12522);
  and g22662 (n12523, n_12140, n_12141);
  not g22663 (n_12142, n12486);
  and g22664 (n12524, n_12142, n12523);
  not g22665 (n_12143, n12523);
  and g22666 (n12525, n12486, n_12143);
  not g22667 (n_12144, n12524);
  not g22668 (n_12145, n12525);
  and g22669 (n12526, n_12144, n_12145);
  not g22670 (n_12146, n12481);
  and g22671 (n12527, n_12146, n12526);
  not g22672 (n_12147, n12526);
  and g22673 (n12528, n12481, n_12147);
  not g22674 (n_12148, n12527);
  not g22675 (n_12149, n12528);
  and g22676 (n12529, n_12148, n_12149);
  not g22677 (n_12150, n12423);
  not g22678 (n_12151, n12529);
  and g22679 (n12530, n_12150, n_12151);
  and g22680 (n12531, n12423, n12529);
  not g22681 (n_12152, n12530);
  not g22682 (n_12153, n12531);
  and g22683 (n12532, n_12152, n_12153);
  and g22684 (n12533, n_10164, n_10165);
  not g22685 (n_12154, n12533);
  and g22686 (n12534, n_10168, n_12154);
  and g22687 (n12535, n10243, n10279);
  not g22688 (n_12155, n12534);
  not g22689 (n_12156, n12535);
  and g22690 (n12536, n_12155, n_12156);
  and g22691 (n12537, n_10156, n_10157);
  not g22692 (n_12157, n12537);
  and g22693 (n12538, n_10160, n_12157);
  not g22697 (n_12158, n12538);
  not g22698 (n_12159, n12541);
  and g22699 (n12542, n_12158, n_12159);
  and g22700 (n12543, n_4018, n_10148);
  and g22701 (n12544, n_10145, n12543);
  not g22702 (n_12160, n12544);
  and g22703 (n12545, n10265, n_12160);
  and g22704 (n12546, n_10152, n10263);
  not g22705 (n_12161, n12545);
  not g22706 (n_12162, n12546);
  and g22707 (n12547, n_12161, n_12162);
  and g22708 (n12548, n_3921, n_10137);
  and g22709 (n12549, n_10134, n12548);
  not g22710 (n_12163, n12549);
  and g22711 (n12550, n10251, n_12163);
  and g22712 (n12551, n_10141, n10249);
  not g22713 (n_12164, n12550);
  not g22714 (n_12165, n12551);
  and g22715 (n12552, n_12164, n_12165);
  not g22716 (n_12166, n12547);
  and g22717 (n12553, n_12166, n12552);
  not g22718 (n_12167, n12552);
  and g22719 (n12554, n12547, n_12167);
  not g22720 (n_12168, n12553);
  not g22721 (n_12169, n12554);
  and g22722 (n12555, n_12168, n_12169);
  not g22723 (n_12170, n12542);
  not g22724 (n_12171, n12555);
  and g22725 (n12556, n_12170, n_12171);
  not g22729 (n_12172, n12556);
  not g22730 (n_12173, n12559);
  and g22731 (n12560, n_12172, n_12173);
  and g22732 (n12561, n_10125, n_10126);
  not g22733 (n_12174, n12561);
  and g22734 (n12562, n_10129, n_12174);
  not g22738 (n_12175, n12562);
  not g22739 (n_12176, n12565);
  and g22740 (n12566, n_12175, n_12176);
  and g22741 (n12567, n_4248, n_10117);
  and g22742 (n12568, n_10114, n12567);
  not g22743 (n_12177, n12568);
  and g22744 (n12569, n10229, n_12177);
  and g22745 (n12570, n_10121, n10227);
  not g22746 (n_12178, n12569);
  not g22747 (n_12179, n12570);
  and g22748 (n12571, n_12178, n_12179);
  and g22749 (n12572, n_4269, n_10106);
  and g22750 (n12573, n_10103, n12572);
  not g22751 (n_12180, n12573);
  and g22752 (n12574, n10215, n_12180);
  and g22753 (n12575, n_10110, n10213);
  not g22754 (n_12181, n12574);
  not g22755 (n_12182, n12575);
  and g22756 (n12576, n_12181, n_12182);
  not g22757 (n_12183, n12571);
  and g22758 (n12577, n_12183, n12576);
  not g22759 (n_12184, n12576);
  and g22760 (n12578, n12571, n_12184);
  not g22761 (n_12185, n12577);
  not g22762 (n_12186, n12578);
  and g22763 (n12579, n_12185, n_12186);
  not g22764 (n_12187, n12566);
  not g22765 (n_12188, n12579);
  and g22766 (n12580, n_12187, n_12188);
  not g22770 (n_12189, n12580);
  not g22771 (n_12190, n12583);
  and g22772 (n12584, n_12189, n_12190);
  not g22773 (n_12191, n12560);
  and g22774 (n12585, n_12191, n12584);
  not g22775 (n_12192, n12584);
  and g22776 (n12586, n12560, n_12192);
  not g22777 (n_12193, n12585);
  not g22778 (n_12194, n12586);
  and g22779 (n12587, n_12193, n_12194);
  not g22780 (n_12195, n12536);
  not g22781 (n_12196, n12587);
  and g22782 (n12588, n_12195, n_12196);
  and g22783 (n12589, n12536, n12587);
  not g22784 (n_12197, n12588);
  not g22785 (n_12198, n12589);
  and g22786 (n12590, n_12197, n_12198);
  not g22787 (n_12199, n12532);
  and g22788 (n12591, n_12199, n12590);
  not g22789 (n_12200, n12590);
  and g22790 (n12592, n_12152, n_12200);
  and g22791 (n12593, n_12153, n12592);
  not g22792 (n_12201, n12591);
  not g22793 (n_12202, n12593);
  and g22794 (n12594, n_12201, n_12202);
  not g22795 (n_12203, n12419);
  not g22796 (n_12204, n12594);
  and g22797 (n12595, n_12203, n_12204);
  and g22798 (n12596, n12419, n12594);
  not g22799 (n_12205, n12595);
  not g22800 (n_12206, n12596);
  and g22801 (n12597, n_12205, n_12206);
  and g22802 (n12598, n_10323, n_10324);
  not g22803 (n_12207, n12598);
  and g22804 (n12599, n_10327, n_12207);
  and g22805 (n12600, n10374, n10454);
  not g22806 (n_12208, n12599);
  not g22807 (n_12209, n12600);
  and g22808 (n12601, n_12208, n_12209);
  and g22809 (n12602, n_10315, n_10316);
  not g22810 (n_12210, n12602);
  and g22811 (n12603, n_10319, n_12210);
  and g22812 (n12604, n10412, n10448);
  not g22813 (n_12211, n12603);
  not g22814 (n_12212, n12604);
  and g22815 (n12605, n_12211, n_12212);
  and g22816 (n12606, n_10307, n_10308);
  not g22817 (n_12213, n12606);
  and g22818 (n12607, n_10311, n_12213);
  not g22822 (n_12214, n12607);
  not g22823 (n_12215, n12610);
  and g22824 (n12611, n_12214, n_12215);
  and g22825 (n12612, n_5979, n_10299);
  and g22826 (n12613, n_10296, n12612);
  not g22827 (n_12216, n12613);
  and g22828 (n12614, n10434, n_12216);
  and g22829 (n12615, n_10303, n10432);
  not g22830 (n_12217, n12614);
  not g22831 (n_12218, n12615);
  and g22832 (n12616, n_12217, n_12218);
  and g22833 (n12617, n_5970, n_10288);
  and g22834 (n12618, n_10285, n12617);
  not g22835 (n_12219, n12618);
  and g22836 (n12619, n10420, n_12219);
  and g22837 (n12620, n_10292, n10418);
  not g22838 (n_12220, n12619);
  not g22839 (n_12221, n12620);
  and g22840 (n12621, n_12220, n_12221);
  not g22841 (n_12222, n12616);
  and g22842 (n12622, n_12222, n12621);
  not g22843 (n_12223, n12621);
  and g22844 (n12623, n12616, n_12223);
  not g22845 (n_12224, n12622);
  not g22846 (n_12225, n12623);
  and g22847 (n12624, n_12224, n_12225);
  not g22848 (n_12226, n12611);
  not g22849 (n_12227, n12624);
  and g22850 (n12625, n_12226, n_12227);
  not g22854 (n_12228, n12625);
  not g22855 (n_12229, n12628);
  and g22856 (n12629, n_12228, n_12229);
  and g22857 (n12630, n_10276, n_10277);
  not g22858 (n_12230, n12630);
  and g22859 (n12631, n_10280, n_12230);
  not g22863 (n_12231, n12631);
  not g22864 (n_12232, n12634);
  and g22865 (n12635, n_12231, n_12232);
  and g22866 (n12636, n_5929, n_10268);
  and g22867 (n12637, n_10265, n12636);
  not g22868 (n_12233, n12637);
  and g22869 (n12638, n10398, n_12233);
  and g22870 (n12639, n_10272, n10396);
  not g22871 (n_12234, n12638);
  not g22872 (n_12235, n12639);
  and g22873 (n12640, n_12234, n_12235);
  and g22874 (n12641, n_5950, n_10257);
  and g22875 (n12642, n_10254, n12641);
  not g22876 (n_12236, n12642);
  and g22877 (n12643, n10384, n_12236);
  and g22878 (n12644, n_10261, n10382);
  not g22879 (n_12237, n12643);
  not g22880 (n_12238, n12644);
  and g22881 (n12645, n_12237, n_12238);
  not g22882 (n_12239, n12640);
  and g22883 (n12646, n_12239, n12645);
  not g22884 (n_12240, n12645);
  and g22885 (n12647, n12640, n_12240);
  not g22886 (n_12241, n12646);
  not g22887 (n_12242, n12647);
  and g22888 (n12648, n_12241, n_12242);
  not g22889 (n_12243, n12635);
  not g22890 (n_12244, n12648);
  and g22891 (n12649, n_12243, n_12244);
  not g22895 (n_12245, n12649);
  not g22896 (n_12246, n12652);
  and g22897 (n12653, n_12245, n_12246);
  not g22898 (n_12247, n12629);
  and g22899 (n12654, n_12247, n12653);
  not g22900 (n_12248, n12653);
  and g22901 (n12655, n12629, n_12248);
  not g22902 (n_12249, n12654);
  not g22903 (n_12250, n12655);
  and g22904 (n12656, n_12249, n_12250);
  not g22905 (n_12251, n12605);
  not g22906 (n_12252, n12656);
  and g22907 (n12657, n_12251, n_12252);
  and g22908 (n12658, n12605, n12656);
  not g22909 (n_12253, n12657);
  not g22910 (n_12254, n12658);
  and g22911 (n12659, n_12253, n_12254);
  and g22912 (n12660, n_10244, n_10245);
  not g22913 (n_12255, n12660);
  and g22914 (n12661, n_10248, n_12255);
  and g22915 (n12662, n10332, n10368);
  not g22916 (n_12256, n12661);
  not g22917 (n_12257, n12662);
  and g22918 (n12663, n_12256, n_12257);
  and g22919 (n12664, n_10236, n_10237);
  not g22920 (n_12258, n12664);
  and g22921 (n12665, n_10240, n_12258);
  not g22925 (n_12259, n12665);
  not g22926 (n_12260, n12668);
  and g22927 (n12669, n_12259, n_12260);
  and g22928 (n12670, n_6031, n_10228);
  and g22929 (n12671, n_10225, n12670);
  not g22930 (n_12261, n12671);
  and g22931 (n12672, n10354, n_12261);
  and g22932 (n12673, n_10232, n10352);
  not g22933 (n_12262, n12672);
  not g22934 (n_12263, n12673);
  and g22935 (n12674, n_12262, n_12263);
  and g22936 (n12675, n_6022, n_10217);
  and g22937 (n12676, n_10214, n12675);
  not g22938 (n_12264, n12676);
  and g22939 (n12677, n10340, n_12264);
  and g22940 (n12678, n_10221, n10338);
  not g22941 (n_12265, n12677);
  not g22942 (n_12266, n12678);
  and g22943 (n12679, n_12265, n_12266);
  not g22944 (n_12267, n12674);
  and g22945 (n12680, n_12267, n12679);
  not g22946 (n_12268, n12679);
  and g22947 (n12681, n12674, n_12268);
  not g22948 (n_12269, n12680);
  not g22949 (n_12270, n12681);
  and g22950 (n12682, n_12269, n_12270);
  not g22951 (n_12271, n12669);
  not g22952 (n_12272, n12682);
  and g22953 (n12683, n_12271, n_12272);
  not g22957 (n_12273, n12683);
  not g22958 (n_12274, n12686);
  and g22959 (n12687, n_12273, n_12274);
  and g22960 (n12688, n_10205, n_10206);
  not g22961 (n_12275, n12688);
  and g22962 (n12689, n_10209, n_12275);
  not g22966 (n_12276, n12689);
  not g22967 (n_12277, n12692);
  and g22968 (n12693, n_12276, n_12277);
  and g22969 (n12694, n_6059, n_10197);
  and g22970 (n12695, n_10194, n12694);
  not g22971 (n_12278, n12695);
  and g22972 (n12696, n10318, n_12278);
  and g22973 (n12697, n_10201, n10316);
  not g22974 (n_12279, n12696);
  not g22975 (n_12280, n12697);
  and g22976 (n12698, n_12279, n_12280);
  and g22977 (n12699, n_6080, n_10186);
  and g22978 (n12700, n_10183, n12699);
  not g22979 (n_12281, n12700);
  and g22980 (n12701, n10304, n_12281);
  and g22981 (n12702, n_10190, n10302);
  not g22982 (n_12282, n12701);
  not g22983 (n_12283, n12702);
  and g22984 (n12703, n_12282, n_12283);
  not g22985 (n_12284, n12698);
  and g22986 (n12704, n_12284, n12703);
  not g22987 (n_12285, n12703);
  and g22988 (n12705, n12698, n_12285);
  not g22989 (n_12286, n12704);
  not g22990 (n_12287, n12705);
  and g22991 (n12706, n_12286, n_12287);
  not g22992 (n_12288, n12693);
  not g22993 (n_12289, n12706);
  and g22994 (n12707, n_12288, n_12289);
  not g22998 (n_12290, n12707);
  not g22999 (n_12291, n12710);
  and g23000 (n12711, n_12290, n_12291);
  not g23001 (n_12292, n12687);
  and g23002 (n12712, n_12292, n12711);
  not g23003 (n_12293, n12711);
  and g23004 (n12713, n12687, n_12293);
  not g23005 (n_12294, n12712);
  not g23006 (n_12295, n12713);
  and g23007 (n12714, n_12294, n_12295);
  not g23008 (n_12296, n12663);
  not g23009 (n_12297, n12714);
  and g23010 (n12715, n_12296, n_12297);
  and g23011 (n12716, n12663, n12714);
  not g23012 (n_12298, n12715);
  not g23013 (n_12299, n12716);
  and g23014 (n12717, n_12298, n_12299);
  not g23015 (n_12300, n12659);
  and g23016 (n12718, n_12300, n12717);
  not g23017 (n_12301, n12717);
  and g23018 (n12719, n12659, n_12301);
  not g23019 (n_12302, n12718);
  not g23020 (n_12303, n12719);
  and g23021 (n12720, n_12302, n_12303);
  not g23022 (n_12304, n12601);
  not g23023 (n_12305, n12720);
  and g23024 (n12721, n_12304, n_12305);
  and g23025 (n12722, n12601, n12720);
  not g23026 (n_12306, n12721);
  not g23027 (n_12307, n12722);
  and g23028 (n12723, n_12306, n_12307);
  not g23029 (n_12308, n12597);
  and g23030 (n12724, n_12308, n12723);
  not g23031 (n_12309, n12723);
  and g23032 (n12725, n_12205, n_12309);
  and g23033 (n12726, n_12206, n12725);
  not g23034 (n_12310, n12724);
  not g23035 (n_12311, n12726);
  and g23036 (n12727, n_12310, n_12311);
  not g23037 (n_12312, n12414);
  not g23038 (n_12313, n12727);
  and g23039 (n12728, n_12312, n_12313);
  and g23040 (n12729, n12414, n12727);
  not g23041 (n_12314, n12728);
  not g23042 (n_12315, n12729);
  and g23043 (n12730, n_12314, n_12315);
  not g23044 (n_12316, n12409);
  and g23045 (n12731, n_12316, n12730);
  not g23046 (n_12317, n12730);
  and g23047 (n12732, n12409, n_12317);
  not g23048 (n_12318, n12731);
  not g23049 (n_12319, n12732);
  and g23050 (n12733, n_12318, n_12319);
  not g23051 (n_12320, n11875);
  not g23052 (n_12321, n12733);
  and g23053 (n12734, n_12320, n_12321);
  and g23054 (n12735, n11875, n12733);
  not g23055 (n_12322, n12734);
  not g23056 (n_12323, n12735);
  and g23057 (n12736, n_12322, n_12323);
  and g23058 (n12737, n_11603, n_11604);
  not g23059 (n_12324, n12737);
  and g23060 (n12738, n_11607, n_12324);
  and g23061 (n12739, n11516, n11860);
  not g23062 (n_12325, n12738);
  not g23063 (n_12326, n12739);
  and g23064 (n12740, n_12325, n_12326);
  and g23065 (n12741, n_11595, n_11596);
  not g23066 (n_12327, n12741);
  and g23067 (n12742, n_11599, n_12327);
  and g23068 (n12743, n11686, n11854);
  not g23069 (n_12328, n12742);
  not g23070 (n_12329, n12743);
  and g23071 (n12744, n_12328, n_12329);
  and g23072 (n12745, n_11587, n_11588);
  not g23073 (n_12330, n12745);
  and g23074 (n12746, n_11591, n_12330);
  and g23075 (n12747, n11768, n11848);
  not g23076 (n_12331, n12746);
  not g23077 (n_12332, n12747);
  and g23078 (n12748, n_12331, n_12332);
  and g23079 (n12749, n_11579, n_11580);
  not g23080 (n_12333, n12749);
  and g23081 (n12750, n_11583, n_12333);
  and g23082 (n12751, n11806, n11842);
  not g23083 (n_12334, n12750);
  not g23084 (n_12335, n12751);
  and g23085 (n12752, n_12334, n_12335);
  and g23086 (n12753, n_11571, n_11572);
  not g23087 (n_12336, n12753);
  and g23088 (n12754, n_11575, n_12336);
  not g23092 (n_12337, n12754);
  not g23093 (n_12338, n12757);
  and g23094 (n12758, n_12337, n_12338);
  and g23095 (n12759, n_1824, n_11563);
  and g23096 (n12760, n_11560, n12759);
  not g23097 (n_12339, n12760);
  and g23098 (n12761, n11828, n_12339);
  and g23099 (n12762, n_11567, n11826);
  not g23100 (n_12340, n12761);
  not g23101 (n_12341, n12762);
  and g23102 (n12763, n_12340, n_12341);
  and g23103 (n12764, n_1727, n_11552);
  and g23104 (n12765, n_11549, n12764);
  not g23105 (n_12342, n12765);
  and g23106 (n12766, n11814, n_12342);
  and g23107 (n12767, n_11556, n11812);
  not g23108 (n_12343, n12766);
  not g23109 (n_12344, n12767);
  and g23110 (n12768, n_12343, n_12344);
  not g23111 (n_12345, n12763);
  and g23112 (n12769, n_12345, n12768);
  not g23113 (n_12346, n12768);
  and g23114 (n12770, n12763, n_12346);
  not g23115 (n_12347, n12769);
  not g23116 (n_12348, n12770);
  and g23117 (n12771, n_12347, n_12348);
  not g23118 (n_12349, n12758);
  not g23119 (n_12350, n12771);
  and g23120 (n12772, n_12349, n_12350);
  not g23124 (n_12351, n12772);
  not g23125 (n_12352, n12775);
  and g23126 (n12776, n_12351, n_12352);
  and g23127 (n12777, n_11540, n_11541);
  not g23128 (n_12353, n12777);
  and g23129 (n12778, n_11544, n_12353);
  not g23133 (n_12354, n12778);
  not g23134 (n_12355, n12781);
  and g23135 (n12782, n_12354, n_12355);
  and g23136 (n12783, n_1500, n_11532);
  and g23137 (n12784, n_11529, n12783);
  not g23138 (n_12356, n12784);
  and g23139 (n12785, n11792, n_12356);
  and g23140 (n12786, n_11536, n11790);
  not g23141 (n_12357, n12785);
  not g23142 (n_12358, n12786);
  and g23143 (n12787, n_12357, n_12358);
  and g23144 (n12788, n_1619, n_11521);
  and g23145 (n12789, n_11518, n12788);
  not g23146 (n_12359, n12789);
  and g23147 (n12790, n11778, n_12359);
  and g23148 (n12791, n_11525, n11776);
  not g23149 (n_12360, n12790);
  not g23150 (n_12361, n12791);
  and g23151 (n12792, n_12360, n_12361);
  not g23152 (n_12362, n12787);
  and g23153 (n12793, n_12362, n12792);
  not g23154 (n_12363, n12792);
  and g23155 (n12794, n12787, n_12363);
  not g23156 (n_12364, n12793);
  not g23157 (n_12365, n12794);
  and g23158 (n12795, n_12364, n_12365);
  not g23159 (n_12366, n12782);
  not g23160 (n_12367, n12795);
  and g23161 (n12796, n_12366, n_12367);
  not g23165 (n_12368, n12796);
  not g23166 (n_12369, n12799);
  and g23167 (n12800, n_12368, n_12369);
  not g23168 (n_12370, n12776);
  and g23169 (n12801, n_12370, n12800);
  not g23170 (n_12371, n12800);
  and g23171 (n12802, n12776, n_12371);
  not g23172 (n_12372, n12801);
  not g23173 (n_12373, n12802);
  and g23174 (n12803, n_12372, n_12373);
  not g23175 (n_12374, n12752);
  not g23176 (n_12375, n12803);
  and g23177 (n12804, n_12374, n_12375);
  and g23178 (n12805, n12752, n12803);
  not g23179 (n_12376, n12804);
  not g23180 (n_12377, n12805);
  and g23181 (n12806, n_12376, n_12377);
  and g23182 (n12807, n_11508, n_11509);
  not g23183 (n_12378, n12807);
  and g23184 (n12808, n_11512, n_12378);
  and g23185 (n12809, n11726, n11762);
  not g23186 (n_12379, n12808);
  not g23187 (n_12380, n12809);
  and g23188 (n12810, n_12379, n_12380);
  and g23189 (n12811, n_11500, n_11501);
  not g23190 (n_12381, n12811);
  and g23191 (n12812, n_11504, n_12381);
  not g23195 (n_12382, n12812);
  not g23196 (n_12383, n12815);
  and g23197 (n12816, n_12382, n_12383);
  and g23198 (n12817, n_1138, n_11492);
  and g23199 (n12818, n_11489, n12817);
  not g23200 (n_12384, n12818);
  and g23201 (n12819, n11748, n_12384);
  and g23202 (n12820, n_11496, n11746);
  not g23203 (n_12385, n12819);
  not g23204 (n_12386, n12820);
  and g23205 (n12821, n_12385, n_12386);
  and g23206 (n12822, n_1041, n_11481);
  and g23207 (n12823, n_11478, n12822);
  not g23208 (n_12387, n12823);
  and g23209 (n12824, n11734, n_12387);
  and g23210 (n12825, n_11485, n11732);
  not g23211 (n_12388, n12824);
  not g23212 (n_12389, n12825);
  and g23213 (n12826, n_12388, n_12389);
  not g23214 (n_12390, n12821);
  and g23215 (n12827, n_12390, n12826);
  not g23216 (n_12391, n12826);
  and g23217 (n12828, n12821, n_12391);
  not g23218 (n_12392, n12827);
  not g23219 (n_12393, n12828);
  and g23220 (n12829, n_12392, n_12393);
  not g23221 (n_12394, n12816);
  not g23222 (n_12395, n12829);
  and g23223 (n12830, n_12394, n_12395);
  not g23227 (n_12396, n12830);
  not g23228 (n_12397, n12833);
  and g23229 (n12834, n_12396, n_12397);
  and g23230 (n12835, n_11469, n_11470);
  not g23231 (n_12398, n12835);
  and g23232 (n12836, n_11473, n_12398);
  not g23236 (n_12399, n12836);
  not g23237 (n_12400, n12839);
  and g23238 (n12840, n_12399, n_12400);
  and g23239 (n12841, n_1368, n_11461);
  and g23240 (n12842, n_11458, n12841);
  not g23241 (n_12401, n12842);
  and g23242 (n12843, n11712, n_12401);
  and g23243 (n12844, n_11465, n11710);
  not g23244 (n_12402, n12843);
  not g23245 (n_12403, n12844);
  and g23246 (n12845, n_12402, n_12403);
  and g23247 (n12846, n_1389, n_11450);
  and g23248 (n12847, n_11447, n12846);
  not g23249 (n_12404, n12847);
  and g23250 (n12848, n11698, n_12404);
  and g23251 (n12849, n_11454, n11696);
  not g23252 (n_12405, n12848);
  not g23253 (n_12406, n12849);
  and g23254 (n12850, n_12405, n_12406);
  not g23255 (n_12407, n12845);
  and g23256 (n12851, n_12407, n12850);
  not g23257 (n_12408, n12850);
  and g23258 (n12852, n12845, n_12408);
  not g23259 (n_12409, n12851);
  not g23260 (n_12410, n12852);
  and g23261 (n12853, n_12409, n_12410);
  not g23262 (n_12411, n12840);
  not g23263 (n_12412, n12853);
  and g23264 (n12854, n_12411, n_12412);
  not g23268 (n_12413, n12854);
  not g23269 (n_12414, n12857);
  and g23270 (n12858, n_12413, n_12414);
  not g23271 (n_12415, n12834);
  and g23272 (n12859, n_12415, n12858);
  not g23273 (n_12416, n12858);
  and g23274 (n12860, n12834, n_12416);
  not g23275 (n_12417, n12859);
  not g23276 (n_12418, n12860);
  and g23277 (n12861, n_12417, n_12418);
  not g23278 (n_12419, n12810);
  not g23279 (n_12420, n12861);
  and g23280 (n12862, n_12419, n_12420);
  and g23281 (n12863, n12810, n12861);
  not g23282 (n_12421, n12862);
  not g23283 (n_12422, n12863);
  and g23284 (n12864, n_12421, n_12422);
  not g23285 (n_12423, n12806);
  and g23286 (n12865, n_12423, n12864);
  not g23287 (n_12424, n12864);
  and g23288 (n12866, n12806, n_12424);
  not g23289 (n_12425, n12865);
  not g23290 (n_12426, n12866);
  and g23291 (n12867, n_12425, n_12426);
  not g23292 (n_12427, n12748);
  not g23293 (n_12428, n12867);
  and g23294 (n12868, n_12427, n_12428);
  and g23295 (n12869, n12748, n12867);
  not g23296 (n_12429, n12868);
  not g23297 (n_12430, n12869);
  and g23298 (n12870, n_12429, n_12430);
  and g23299 (n12871, n_11436, n_11437);
  not g23300 (n_12431, n12871);
  and g23301 (n12872, n_11440, n_12431);
  and g23302 (n12873, n11600, n11680);
  not g23303 (n_12432, n12872);
  not g23304 (n_12433, n12873);
  and g23305 (n12874, n_12432, n_12433);
  and g23306 (n12875, n_11428, n_11429);
  not g23307 (n_12434, n12875);
  and g23308 (n12876, n_11432, n_12434);
  and g23309 (n12877, n11638, n11674);
  not g23310 (n_12435, n12876);
  not g23311 (n_12436, n12877);
  and g23312 (n12878, n_12435, n_12436);
  and g23313 (n12879, n_11420, n_11421);
  not g23314 (n_12437, n12879);
  and g23315 (n12880, n_11424, n_12437);
  not g23319 (n_12438, n12880);
  not g23320 (n_12439, n12883);
  and g23321 (n12884, n_12438, n_12439);
  and g23322 (n12885, n_418, n_11412);
  and g23323 (n12886, n_11409, n12885);
  not g23324 (n_12440, n12886);
  and g23325 (n12887, n11660, n_12440);
  and g23326 (n12888, n_11416, n11658);
  not g23327 (n_12441, n12887);
  not g23328 (n_12442, n12888);
  and g23329 (n12889, n_12441, n_12442);
  and g23330 (n12890, n_321, n_11401);
  and g23331 (n12891, n_11398, n12890);
  not g23332 (n_12443, n12891);
  and g23333 (n12892, n11646, n_12443);
  and g23334 (n12893, n_11405, n11644);
  not g23335 (n_12444, n12892);
  not g23336 (n_12445, n12893);
  and g23337 (n12894, n_12444, n_12445);
  not g23338 (n_12446, n12889);
  and g23339 (n12895, n_12446, n12894);
  not g23340 (n_12447, n12894);
  and g23341 (n12896, n12889, n_12447);
  not g23342 (n_12448, n12895);
  not g23343 (n_12449, n12896);
  and g23344 (n12897, n_12448, n_12449);
  not g23345 (n_12450, n12884);
  not g23346 (n_12451, n12897);
  and g23347 (n12898, n_12450, n_12451);
  not g23351 (n_12452, n12898);
  not g23352 (n_12453, n12901);
  and g23353 (n12902, n_12452, n_12453);
  and g23354 (n12903, n_11389, n_11390);
  not g23355 (n_12454, n12903);
  and g23356 (n12904, n_11393, n_12454);
  not g23360 (n_12455, n12904);
  not g23361 (n_12456, n12907);
  and g23362 (n12908, n_12455, n_12456);
  and g23363 (n12909, n_94, n_11381);
  and g23364 (n12910, n_11378, n12909);
  not g23365 (n_12457, n12910);
  and g23366 (n12911, n11624, n_12457);
  and g23367 (n12912, n_11385, n11622);
  not g23368 (n_12458, n12911);
  not g23369 (n_12459, n12912);
  and g23370 (n12913, n_12458, n_12459);
  and g23371 (n12914, n_213, n_11370);
  and g23372 (n12915, n_11367, n12914);
  not g23373 (n_12460, n12915);
  and g23374 (n12916, n11610, n_12460);
  and g23375 (n12917, n_11374, n11608);
  not g23376 (n_12461, n12916);
  not g23377 (n_12462, n12917);
  and g23378 (n12918, n_12461, n_12462);
  not g23379 (n_12463, n12913);
  and g23380 (n12919, n_12463, n12918);
  not g23381 (n_12464, n12918);
  and g23382 (n12920, n12913, n_12464);
  not g23383 (n_12465, n12919);
  not g23384 (n_12466, n12920);
  and g23385 (n12921, n_12465, n_12466);
  not g23386 (n_12467, n12908);
  not g23387 (n_12468, n12921);
  and g23388 (n12922, n_12467, n_12468);
  not g23392 (n_12469, n12922);
  not g23393 (n_12470, n12925);
  and g23394 (n12926, n_12469, n_12470);
  not g23395 (n_12471, n12902);
  and g23396 (n12927, n_12471, n12926);
  not g23397 (n_12472, n12926);
  and g23398 (n12928, n12902, n_12472);
  not g23399 (n_12473, n12927);
  not g23400 (n_12474, n12928);
  and g23401 (n12929, n_12473, n_12474);
  not g23402 (n_12475, n12878);
  not g23403 (n_12476, n12929);
  and g23404 (n12930, n_12475, n_12476);
  and g23405 (n12931, n12878, n12929);
  not g23406 (n_12477, n12930);
  not g23407 (n_12478, n12931);
  and g23408 (n12932, n_12477, n_12478);
  and g23409 (n12933, n_11357, n_11358);
  not g23410 (n_12479, n12933);
  and g23411 (n12934, n_11361, n_12479);
  and g23412 (n12935, n11558, n11594);
  not g23413 (n_12480, n12934);
  not g23414 (n_12481, n12935);
  and g23415 (n12936, n_12480, n_12481);
  and g23416 (n12937, n_11349, n_11350);
  not g23417 (n_12482, n12937);
  and g23418 (n12938, n_11353, n_12482);
  not g23422 (n_12483, n12938);
  not g23423 (n_12484, n12941);
  and g23424 (n12942, n_12483, n_12484);
  and g23425 (n12943, n_870, n_11341);
  and g23426 (n12944, n_11338, n12943);
  not g23427 (n_12485, n12944);
  and g23428 (n12945, n11580, n_12485);
  and g23429 (n12946, n_11345, n11578);
  not g23430 (n_12486, n12945);
  not g23431 (n_12487, n12946);
  and g23432 (n12947, n_12486, n_12487);
  and g23433 (n12948, n_861, n_11330);
  and g23434 (n12949, n_11327, n12948);
  not g23435 (n_12488, n12949);
  and g23436 (n12950, n11566, n_12488);
  and g23437 (n12951, n_11334, n11564);
  not g23438 (n_12489, n12950);
  not g23439 (n_12490, n12951);
  and g23440 (n12952, n_12489, n_12490);
  not g23441 (n_12491, n12947);
  and g23442 (n12953, n_12491, n12952);
  not g23443 (n_12492, n12952);
  and g23444 (n12954, n12947, n_12492);
  not g23445 (n_12493, n12953);
  not g23446 (n_12494, n12954);
  and g23447 (n12955, n_12493, n_12494);
  not g23448 (n_12495, n12942);
  not g23449 (n_12496, n12955);
  and g23450 (n12956, n_12495, n_12496);
  not g23454 (n_12497, n12956);
  not g23455 (n_12498, n12959);
  and g23456 (n12960, n_12497, n_12498);
  and g23457 (n12961, n_11318, n_11319);
  not g23458 (n_12499, n12961);
  and g23459 (n12962, n_11322, n_12499);
  not g23463 (n_12500, n12962);
  not g23464 (n_12501, n12965);
  and g23465 (n12966, n_12500, n_12501);
  and g23466 (n12967, n_898, n_11310);
  and g23467 (n12968, n_11307, n12967);
  not g23468 (n_12502, n12968);
  and g23469 (n12969, n11544, n_12502);
  and g23470 (n12970, n_11314, n11542);
  not g23471 (n_12503, n12969);
  not g23472 (n_12504, n12970);
  and g23473 (n12971, n_12503, n_12504);
  and g23474 (n12972, n_919, n_11299);
  and g23475 (n12973, n_11296, n12972);
  not g23476 (n_12505, n12973);
  and g23477 (n12974, n11530, n_12505);
  and g23478 (n12975, n_11303, n11528);
  not g23479 (n_12506, n12974);
  not g23480 (n_12507, n12975);
  and g23481 (n12976, n_12506, n_12507);
  not g23482 (n_12508, n12971);
  and g23483 (n12977, n_12508, n12976);
  not g23484 (n_12509, n12976);
  and g23485 (n12978, n12971, n_12509);
  not g23486 (n_12510, n12977);
  not g23487 (n_12511, n12978);
  and g23488 (n12979, n_12510, n_12511);
  not g23489 (n_12512, n12966);
  not g23490 (n_12513, n12979);
  and g23491 (n12980, n_12512, n_12513);
  not g23495 (n_12514, n12980);
  not g23496 (n_12515, n12983);
  and g23497 (n12984, n_12514, n_12515);
  not g23498 (n_12516, n12960);
  and g23499 (n12985, n_12516, n12984);
  not g23500 (n_12517, n12984);
  and g23501 (n12986, n12960, n_12517);
  not g23502 (n_12518, n12985);
  not g23503 (n_12519, n12986);
  and g23504 (n12987, n_12518, n_12519);
  not g23505 (n_12520, n12936);
  not g23506 (n_12521, n12987);
  and g23507 (n12988, n_12520, n_12521);
  and g23508 (n12989, n12936, n12987);
  not g23509 (n_12522, n12988);
  not g23510 (n_12523, n12989);
  and g23511 (n12990, n_12522, n_12523);
  not g23512 (n_12524, n12932);
  and g23513 (n12991, n_12524, n12990);
  not g23514 (n_12525, n12990);
  and g23515 (n12992, n12932, n_12525);
  not g23516 (n_12526, n12991);
  not g23517 (n_12527, n12992);
  and g23518 (n12993, n_12526, n_12527);
  not g23519 (n_12528, n12874);
  not g23520 (n_12529, n12993);
  and g23521 (n12994, n_12528, n_12529);
  and g23522 (n12995, n12874, n12993);
  not g23523 (n_12530, n12994);
  not g23524 (n_12531, n12995);
  and g23525 (n12996, n_12530, n_12531);
  not g23526 (n_12532, n12870);
  and g23527 (n12997, n_12532, n12996);
  not g23528 (n_12533, n12996);
  and g23529 (n12998, n12870, n_12533);
  not g23530 (n_12534, n12997);
  not g23531 (n_12535, n12998);
  and g23532 (n12999, n_12534, n_12535);
  not g23533 (n_12536, n12744);
  not g23534 (n_12537, n12999);
  and g23535 (n13000, n_12536, n_12537);
  and g23536 (n13001, n12744, n12999);
  not g23537 (n_12538, n13000);
  not g23538 (n_12539, n13001);
  and g23539 (n13002, n_12538, n_12539);
  and g23540 (n13003, n_11284, n_11285);
  not g23541 (n_12540, n13003);
  and g23542 (n13004, n_11288, n_12540);
  and g23543 (n13005, n11342, n11510);
  not g23544 (n_12541, n13004);
  not g23545 (n_12542, n13005);
  and g23546 (n13006, n_12541, n_12542);
  and g23547 (n13007, n_11276, n_11277);
  not g23548 (n_12543, n13007);
  and g23549 (n13008, n_11280, n_12543);
  and g23550 (n13009, n11424, n11504);
  not g23551 (n_12544, n13008);
  not g23552 (n_12545, n13009);
  and g23553 (n13010, n_12544, n_12545);
  and g23554 (n13011, n_11268, n_11269);
  not g23555 (n_12546, n13011);
  and g23556 (n13012, n_11272, n_12546);
  and g23557 (n13013, n11462, n11498);
  not g23558 (n_12547, n13012);
  not g23559 (n_12548, n13013);
  and g23560 (n13014, n_12547, n_12548);
  and g23561 (n13015, n_11260, n_11261);
  not g23562 (n_12549, n13015);
  and g23563 (n13016, n_11264, n_12549);
  not g23567 (n_12550, n13016);
  not g23568 (n_12551, n13019);
  and g23569 (n13020, n_12550, n_12551);
  and g23570 (n13021, n_3584, n_11252);
  and g23571 (n13022, n_11249, n13021);
  not g23572 (n_12552, n13022);
  and g23573 (n13023, n11484, n_12552);
  and g23574 (n13024, n_11256, n11482);
  not g23575 (n_12553, n13023);
  not g23576 (n_12554, n13024);
  and g23577 (n13025, n_12553, n_12554);
  and g23578 (n13026, n_3575, n_11241);
  and g23579 (n13027, n_11238, n13026);
  not g23580 (n_12555, n13027);
  and g23581 (n13028, n11470, n_12555);
  and g23582 (n13029, n_11245, n11468);
  not g23583 (n_12556, n13028);
  not g23584 (n_12557, n13029);
  and g23585 (n13030, n_12556, n_12557);
  not g23586 (n_12558, n13025);
  and g23587 (n13031, n_12558, n13030);
  not g23588 (n_12559, n13030);
  and g23589 (n13032, n13025, n_12559);
  not g23590 (n_12560, n13031);
  not g23591 (n_12561, n13032);
  and g23592 (n13033, n_12560, n_12561);
  not g23593 (n_12562, n13020);
  not g23594 (n_12563, n13033);
  and g23595 (n13034, n_12562, n_12563);
  not g23599 (n_12564, n13034);
  not g23600 (n_12565, n13037);
  and g23601 (n13038, n_12564, n_12565);
  and g23602 (n13039, n_11229, n_11230);
  not g23603 (n_12566, n13039);
  and g23604 (n13040, n_11233, n_12566);
  not g23608 (n_12567, n13040);
  not g23609 (n_12568, n13043);
  and g23610 (n13044, n_12567, n_12568);
  and g23611 (n13045, n_3534, n_11221);
  and g23612 (n13046, n_11218, n13045);
  not g23613 (n_12569, n13046);
  and g23614 (n13047, n11448, n_12569);
  and g23615 (n13048, n_11225, n11446);
  not g23616 (n_12570, n13047);
  not g23617 (n_12571, n13048);
  and g23618 (n13049, n_12570, n_12571);
  and g23619 (n13050, n_3555, n_11210);
  and g23620 (n13051, n_11207, n13050);
  not g23621 (n_12572, n13051);
  and g23622 (n13052, n11434, n_12572);
  and g23623 (n13053, n_11214, n11432);
  not g23624 (n_12573, n13052);
  not g23625 (n_12574, n13053);
  and g23626 (n13054, n_12573, n_12574);
  not g23627 (n_12575, n13049);
  and g23628 (n13055, n_12575, n13054);
  not g23629 (n_12576, n13054);
  and g23630 (n13056, n13049, n_12576);
  not g23631 (n_12577, n13055);
  not g23632 (n_12578, n13056);
  and g23633 (n13057, n_12577, n_12578);
  not g23634 (n_12579, n13044);
  not g23635 (n_12580, n13057);
  and g23636 (n13058, n_12579, n_12580);
  not g23640 (n_12581, n13058);
  not g23641 (n_12582, n13061);
  and g23642 (n13062, n_12581, n_12582);
  not g23643 (n_12583, n13038);
  and g23644 (n13063, n_12583, n13062);
  not g23645 (n_12584, n13062);
  and g23646 (n13064, n13038, n_12584);
  not g23647 (n_12585, n13063);
  not g23648 (n_12586, n13064);
  and g23649 (n13065, n_12585, n_12586);
  not g23650 (n_12587, n13014);
  not g23651 (n_12588, n13065);
  and g23652 (n13066, n_12587, n_12588);
  and g23653 (n13067, n13014, n13065);
  not g23654 (n_12589, n13066);
  not g23655 (n_12590, n13067);
  and g23656 (n13068, n_12589, n_12590);
  and g23657 (n13069, n_11197, n_11198);
  not g23658 (n_12591, n13069);
  and g23659 (n13070, n_11201, n_12591);
  and g23660 (n13071, n11382, n11418);
  not g23661 (n_12592, n13070);
  not g23662 (n_12593, n13071);
  and g23663 (n13072, n_12592, n_12593);
  and g23664 (n13073, n_11189, n_11190);
  not g23665 (n_12594, n13073);
  and g23666 (n13074, n_11193, n_12594);
  not g23670 (n_12595, n13074);
  not g23671 (n_12596, n13077);
  and g23672 (n13078, n_12595, n_12596);
  and g23673 (n13079, n_3462, n_11181);
  and g23674 (n13080, n_11178, n13079);
  not g23675 (n_12597, n13080);
  and g23676 (n13081, n11404, n_12597);
  and g23677 (n13082, n_11185, n11402);
  not g23678 (n_12598, n13081);
  not g23679 (n_12599, n13082);
  and g23680 (n13083, n_12598, n_12599);
  and g23681 (n13084, n_3453, n_11170);
  and g23682 (n13085, n_11167, n13084);
  not g23683 (n_12600, n13085);
  and g23684 (n13086, n11390, n_12600);
  and g23685 (n13087, n_11174, n11388);
  not g23686 (n_12601, n13086);
  not g23687 (n_12602, n13087);
  and g23688 (n13088, n_12601, n_12602);
  not g23689 (n_12603, n13083);
  and g23690 (n13089, n_12603, n13088);
  not g23691 (n_12604, n13088);
  and g23692 (n13090, n13083, n_12604);
  not g23693 (n_12605, n13089);
  not g23694 (n_12606, n13090);
  and g23695 (n13091, n_12605, n_12606);
  not g23696 (n_12607, n13078);
  not g23697 (n_12608, n13091);
  and g23698 (n13092, n_12607, n_12608);
  not g23702 (n_12609, n13092);
  not g23703 (n_12610, n13095);
  and g23704 (n13096, n_12609, n_12610);
  and g23705 (n13097, n_11158, n_11159);
  not g23706 (n_12611, n13097);
  and g23707 (n13098, n_11162, n_12611);
  not g23711 (n_12612, n13098);
  not g23712 (n_12613, n13101);
  and g23713 (n13102, n_12612, n_12613);
  and g23714 (n13103, n_3490, n_11150);
  and g23715 (n13104, n_11147, n13103);
  not g23716 (n_12614, n13104);
  and g23717 (n13105, n11368, n_12614);
  and g23718 (n13106, n_11154, n11366);
  not g23719 (n_12615, n13105);
  not g23720 (n_12616, n13106);
  and g23721 (n13107, n_12615, n_12616);
  and g23722 (n13108, n_3511, n_11139);
  and g23723 (n13109, n_11136, n13108);
  not g23724 (n_12617, n13109);
  and g23725 (n13110, n11354, n_12617);
  and g23726 (n13111, n_11143, n11352);
  not g23727 (n_12618, n13110);
  not g23728 (n_12619, n13111);
  and g23729 (n13112, n_12618, n_12619);
  not g23730 (n_12620, n13107);
  and g23731 (n13113, n_12620, n13112);
  not g23732 (n_12621, n13112);
  and g23733 (n13114, n13107, n_12621);
  not g23734 (n_12622, n13113);
  not g23735 (n_12623, n13114);
  and g23736 (n13115, n_12622, n_12623);
  not g23737 (n_12624, n13102);
  not g23738 (n_12625, n13115);
  and g23739 (n13116, n_12624, n_12625);
  not g23743 (n_12626, n13116);
  not g23744 (n_12627, n13119);
  and g23745 (n13120, n_12626, n_12627);
  not g23746 (n_12628, n13096);
  and g23747 (n13121, n_12628, n13120);
  not g23748 (n_12629, n13120);
  and g23749 (n13122, n13096, n_12629);
  not g23750 (n_12630, n13121);
  not g23751 (n_12631, n13122);
  and g23752 (n13123, n_12630, n_12631);
  not g23753 (n_12632, n13072);
  not g23754 (n_12633, n13123);
  and g23755 (n13124, n_12632, n_12633);
  and g23756 (n13125, n13072, n13123);
  not g23757 (n_12634, n13124);
  not g23758 (n_12635, n13125);
  and g23759 (n13126, n_12634, n_12635);
  not g23760 (n_12636, n13068);
  and g23761 (n13127, n_12636, n13126);
  not g23762 (n_12637, n13126);
  and g23763 (n13128, n13068, n_12637);
  not g23764 (n_12638, n13127);
  not g23765 (n_12639, n13128);
  and g23766 (n13129, n_12638, n_12639);
  not g23767 (n_12640, n13010);
  not g23768 (n_12641, n13129);
  and g23769 (n13130, n_12640, n_12641);
  and g23770 (n13131, n13010, n13129);
  not g23771 (n_12642, n13130);
  not g23772 (n_12643, n13131);
  and g23773 (n13132, n_12642, n_12643);
  and g23774 (n13133, n_11125, n_11126);
  not g23775 (n_12644, n13133);
  and g23776 (n13134, n_11129, n_12644);
  and g23777 (n13135, n11256, n11336);
  not g23778 (n_12645, n13134);
  not g23779 (n_12646, n13135);
  and g23780 (n13136, n_12645, n_12646);
  and g23781 (n13137, n_11117, n_11118);
  not g23782 (n_12647, n13137);
  and g23783 (n13138, n_11121, n_12647);
  and g23784 (n13139, n11294, n11330);
  not g23785 (n_12648, n13138);
  not g23786 (n_12649, n13139);
  and g23787 (n13140, n_12648, n_12649);
  and g23788 (n13141, n_11109, n_11110);
  not g23789 (n_12650, n13141);
  and g23790 (n13142, n_11113, n_12650);
  not g23794 (n_12651, n13142);
  not g23795 (n_12652, n13145);
  and g23796 (n13146, n_12651, n_12652);
  and g23797 (n13147, n_3684, n_11101);
  and g23798 (n13148, n_11098, n13147);
  not g23799 (n_12653, n13148);
  and g23800 (n13149, n11316, n_12653);
  and g23801 (n13150, n_11105, n11314);
  not g23802 (n_12654, n13149);
  not g23803 (n_12655, n13150);
  and g23804 (n13151, n_12654, n_12655);
  and g23805 (n13152, n_3675, n_11090);
  and g23806 (n13153, n_11087, n13152);
  not g23807 (n_12656, n13153);
  and g23808 (n13154, n11302, n_12656);
  and g23809 (n13155, n_11094, n11300);
  not g23810 (n_12657, n13154);
  not g23811 (n_12658, n13155);
  and g23812 (n13156, n_12657, n_12658);
  not g23813 (n_12659, n13151);
  and g23814 (n13157, n_12659, n13156);
  not g23815 (n_12660, n13156);
  and g23816 (n13158, n13151, n_12660);
  not g23817 (n_12661, n13157);
  not g23818 (n_12662, n13158);
  and g23819 (n13159, n_12661, n_12662);
  not g23820 (n_12663, n13146);
  not g23821 (n_12664, n13159);
  and g23822 (n13160, n_12663, n_12664);
  not g23826 (n_12665, n13160);
  not g23827 (n_12666, n13163);
  and g23828 (n13164, n_12665, n_12666);
  and g23829 (n13165, n_11078, n_11079);
  not g23830 (n_12667, n13165);
  and g23831 (n13166, n_11082, n_12667);
  not g23835 (n_12668, n13166);
  not g23836 (n_12669, n13169);
  and g23837 (n13170, n_12668, n_12669);
  and g23838 (n13171, n_3634, n_11070);
  and g23839 (n13172, n_11067, n13171);
  not g23840 (n_12670, n13172);
  and g23841 (n13173, n11280, n_12670);
  and g23842 (n13174, n_11074, n11278);
  not g23843 (n_12671, n13173);
  not g23844 (n_12672, n13174);
  and g23845 (n13175, n_12671, n_12672);
  and g23846 (n13176, n_3655, n_11059);
  and g23847 (n13177, n_11056, n13176);
  not g23848 (n_12673, n13177);
  and g23849 (n13178, n11266, n_12673);
  and g23850 (n13179, n_11063, n11264);
  not g23851 (n_12674, n13178);
  not g23852 (n_12675, n13179);
  and g23853 (n13180, n_12674, n_12675);
  not g23854 (n_12676, n13175);
  and g23855 (n13181, n_12676, n13180);
  not g23856 (n_12677, n13180);
  and g23857 (n13182, n13175, n_12677);
  not g23858 (n_12678, n13181);
  not g23859 (n_12679, n13182);
  and g23860 (n13183, n_12678, n_12679);
  not g23861 (n_12680, n13170);
  not g23862 (n_12681, n13183);
  and g23863 (n13184, n_12680, n_12681);
  not g23867 (n_12682, n13184);
  not g23868 (n_12683, n13187);
  and g23869 (n13188, n_12682, n_12683);
  not g23870 (n_12684, n13164);
  and g23871 (n13189, n_12684, n13188);
  not g23872 (n_12685, n13188);
  and g23873 (n13190, n13164, n_12685);
  not g23874 (n_12686, n13189);
  not g23875 (n_12687, n13190);
  and g23876 (n13191, n_12686, n_12687);
  not g23877 (n_12688, n13140);
  not g23878 (n_12689, n13191);
  and g23879 (n13192, n_12688, n_12689);
  and g23880 (n13193, n13140, n13191);
  not g23881 (n_12690, n13192);
  not g23882 (n_12691, n13193);
  and g23883 (n13194, n_12690, n_12691);
  and g23884 (n13195, n_11046, n_11047);
  not g23885 (n_12692, n13195);
  and g23886 (n13196, n_11050, n_12692);
  and g23887 (n13197, n11214, n11250);
  not g23888 (n_12693, n13196);
  not g23889 (n_12694, n13197);
  and g23890 (n13198, n_12693, n_12694);
  and g23891 (n13199, n_11038, n_11039);
  not g23892 (n_12695, n13199);
  and g23893 (n13200, n_11042, n_12695);
  not g23897 (n_12696, n13200);
  not g23898 (n_12697, n13203);
  and g23899 (n13204, n_12696, n_12697);
  and g23900 (n13205, n_3736, n_11030);
  and g23901 (n13206, n_11027, n13205);
  not g23902 (n_12698, n13206);
  and g23903 (n13207, n11236, n_12698);
  and g23904 (n13208, n_11034, n11234);
  not g23905 (n_12699, n13207);
  not g23906 (n_12700, n13208);
  and g23907 (n13209, n_12699, n_12700);
  and g23908 (n13210, n_3727, n_11019);
  and g23909 (n13211, n_11016, n13210);
  not g23910 (n_12701, n13211);
  and g23911 (n13212, n11222, n_12701);
  and g23912 (n13213, n_11023, n11220);
  not g23913 (n_12702, n13212);
  not g23914 (n_12703, n13213);
  and g23915 (n13214, n_12702, n_12703);
  not g23916 (n_12704, n13209);
  and g23917 (n13215, n_12704, n13214);
  not g23918 (n_12705, n13214);
  and g23919 (n13216, n13209, n_12705);
  not g23920 (n_12706, n13215);
  not g23921 (n_12707, n13216);
  and g23922 (n13217, n_12706, n_12707);
  not g23923 (n_12708, n13204);
  not g23924 (n_12709, n13217);
  and g23925 (n13218, n_12708, n_12709);
  not g23929 (n_12710, n13218);
  not g23930 (n_12711, n13221);
  and g23931 (n13222, n_12710, n_12711);
  and g23932 (n13223, n_11007, n_11008);
  not g23933 (n_12712, n13223);
  and g23934 (n13224, n_11011, n_12712);
  not g23938 (n_12713, n13224);
  not g23939 (n_12714, n13227);
  and g23940 (n13228, n_12713, n_12714);
  and g23941 (n13229, n_3764, n_10999);
  and g23942 (n13230, n_10996, n13229);
  not g23943 (n_12715, n13230);
  and g23944 (n13231, n11200, n_12715);
  and g23945 (n13232, n_11003, n11198);
  not g23946 (n_12716, n13231);
  not g23947 (n_12717, n13232);
  and g23948 (n13233, n_12716, n_12717);
  and g23949 (n13234, n_3785, n_10988);
  and g23950 (n13235, n_10985, n13234);
  not g23951 (n_12718, n13235);
  and g23952 (n13236, n11186, n_12718);
  and g23953 (n13237, n_10992, n11184);
  not g23954 (n_12719, n13236);
  not g23955 (n_12720, n13237);
  and g23956 (n13238, n_12719, n_12720);
  not g23957 (n_12721, n13233);
  and g23958 (n13239, n_12721, n13238);
  not g23959 (n_12722, n13238);
  and g23960 (n13240, n13233, n_12722);
  not g23961 (n_12723, n13239);
  not g23962 (n_12724, n13240);
  and g23963 (n13241, n_12723, n_12724);
  not g23964 (n_12725, n13228);
  not g23965 (n_12726, n13241);
  and g23966 (n13242, n_12725, n_12726);
  not g23970 (n_12727, n13242);
  not g23971 (n_12728, n13245);
  and g23972 (n13246, n_12727, n_12728);
  not g23973 (n_12729, n13222);
  and g23974 (n13247, n_12729, n13246);
  not g23975 (n_12730, n13246);
  and g23976 (n13248, n13222, n_12730);
  not g23977 (n_12731, n13247);
  not g23978 (n_12732, n13248);
  and g23979 (n13249, n_12731, n_12732);
  not g23980 (n_12733, n13198);
  not g23981 (n_12734, n13249);
  and g23982 (n13250, n_12733, n_12734);
  and g23983 (n13251, n13198, n13249);
  not g23984 (n_12735, n13250);
  not g23985 (n_12736, n13251);
  and g23986 (n13252, n_12735, n_12736);
  not g23987 (n_12737, n13194);
  and g23988 (n13253, n_12737, n13252);
  not g23989 (n_12738, n13252);
  and g23990 (n13254, n13194, n_12738);
  not g23991 (n_12739, n13253);
  not g23992 (n_12740, n13254);
  and g23993 (n13255, n_12739, n_12740);
  not g23994 (n_12741, n13136);
  not g23995 (n_12742, n13255);
  and g23996 (n13256, n_12741, n_12742);
  and g23997 (n13257, n13136, n13255);
  not g23998 (n_12743, n13256);
  not g23999 (n_12744, n13257);
  and g24000 (n13258, n_12743, n_12744);
  not g24001 (n_12745, n13132);
  and g24002 (n13259, n_12745, n13258);
  not g24003 (n_12746, n13258);
  and g24004 (n13260, n13132, n_12746);
  not g24005 (n_12747, n13259);
  not g24006 (n_12748, n13260);
  and g24007 (n13261, n_12747, n_12748);
  not g24008 (n_12749, n13006);
  not g24009 (n_12750, n13261);
  and g24010 (n13262, n_12749, n_12750);
  and g24011 (n13263, n13006, n13261);
  not g24012 (n_12751, n13262);
  not g24013 (n_12752, n13263);
  and g24014 (n13264, n_12751, n_12752);
  not g24015 (n_12753, n13002);
  and g24016 (n13265, n_12753, n13264);
  not g24017 (n_12754, n13264);
  and g24018 (n13266, n13002, n_12754);
  not g24019 (n_12755, n13265);
  not g24020 (n_12756, n13266);
  and g24021 (n13267, n_12755, n_12756);
  not g24022 (n_12757, n12740);
  not g24023 (n_12758, n13267);
  and g24024 (n13268, n_12757, n_12758);
  and g24025 (n13269, n12740, n13267);
  not g24026 (n_12759, n13268);
  not g24027 (n_12760, n13269);
  and g24028 (n13270, n_12759, n_12760);
  not g24029 (n_12761, n12736);
  not g24030 (n_12762, n13270);
  and g24031 (n13271, n_12761, n_12762);
  not g24032 (n_12763, n11871);
  not g24033 (n_12764, n13271);
  and g24034 (n13272, n_12763, n_12764);
  and g24035 (n13273, n_12322, n13270);
  and g24036 (n13274, n_12323, n13273);
  not g24037 (n_12765, n13272);
  not g24038 (n_12766, n13274);
  and g24039 (n13275, n_12765, n_12766);
  and g24040 (n13276, n_12316, n_12317);
  not g24041 (n_12767, n13276);
  and g24042 (n13277, n_12320, n_12767);
  and g24043 (n13278, n12409, n12730);
  not g24044 (n_12768, n13277);
  not g24045 (n_12769, n13278);
  and g24046 (n13279, n_12768, n_12769);
  and g24047 (n13280, n_12308, n_12309);
  not g24048 (n_12770, n13280);
  and g24049 (n13281, n_12312, n_12770);
  and g24050 (n13282, n_12205, n12723);
  and g24051 (n13283, n_12206, n13282);
  not g24052 (n_12771, n13281);
  not g24053 (n_12772, n13283);
  and g24054 (n13284, n_12771, n_12772);
  and g24055 (n13285, n_12199, n_12200);
  not g24056 (n_12773, n13285);
  and g24057 (n13286, n_12203, n_12773);
  and g24058 (n13287, n_12152, n12590);
  and g24059 (n13288, n_12153, n13287);
  not g24060 (n_12774, n13286);
  not g24061 (n_12775, n13288);
  and g24062 (n13289, n_12774, n_12775);
  and g24063 (n13290, n_12146, n_12147);
  not g24064 (n_12776, n13290);
  and g24065 (n13291, n_12150, n_12776);
  and g24066 (n13292, n12481, n12526);
  not g24067 (n_12777, n13291);
  not g24068 (n_12778, n13292);
  and g24069 (n13293, n_12777, n_12778);
  and g24070 (n13294, n_12142, n_12140);
  not g24071 (n_12779, n13294);
  and g24072 (n13295, n_12141, n_12779);
  and g24073 (n13296, n12507, n12512);
  not g24074 (n_12780, n13296);
  and g24075 (n13297, n_12134, n_12780);
  and g24076 (n13298, n_12130, n_12131);
  not g24077 (n_12781, n13298);
  and g24078 (n13299, n_12119, n_12781);
  not g24079 (n_12782, n13297);
  and g24080 (n13300, n_12782, n13299);
  and g24081 (n13301, n_12782, n_12781);
  not g24082 (n_12783, n13301);
  and g24083 (n13302, n12493, n_12783);
  not g24084 (n_12784, n13300);
  not g24085 (n_12785, n13302);
  and g24086 (n13303, n_12784, n_12785);
  not g24087 (n_12786, n13295);
  and g24088 (n13304, n_12786, n13303);
  not g24089 (n_12787, n13303);
  and g24090 (n13305, n_12141, n_12787);
  and g24091 (n13306, n_12779, n13305);
  not g24092 (n_12788, n13304);
  not g24093 (n_12789, n13306);
  and g24094 (n13307, n_12788, n_12789);
  and g24095 (n13308, n_12103, n_12104);
  not g24096 (n_12790, n13308);
  and g24097 (n13309, n_12107, n_12790);
  not g24101 (n_12791, n13309);
  not g24102 (n_12792, n13312);
  and g24103 (n13313, n_12791, n_12792);
  and g24104 (n13314, n12438, n12443);
  not g24105 (n_12793, n13314);
  and g24106 (n13315, n_12082, n_12793);
  and g24107 (n13316, n_12078, n_12079);
  not g24108 (n_12794, n13315);
  not g24109 (n_12795, n13316);
  and g24110 (n13317, n_12794, n_12795);
  and g24111 (n13318, n12462, n12467);
  not g24112 (n_12796, n13318);
  and g24113 (n13319, n_12099, n_12796);
  and g24114 (n13320, n_12095, n_12096);
  not g24115 (n_12797, n13319);
  not g24116 (n_12798, n13320);
  and g24117 (n13321, n_12797, n_12798);
  not g24118 (n_12799, n13317);
  and g24119 (n13322, n_12799, n13321);
  not g24120 (n_12800, n13321);
  and g24121 (n13323, n13317, n_12800);
  not g24122 (n_12801, n13322);
  not g24123 (n_12802, n13323);
  and g24124 (n13324, n_12801, n_12802);
  not g24125 (n_12803, n13313);
  not g24126 (n_12804, n13324);
  and g24127 (n13325, n_12803, n_12804);
  not g24131 (n_12805, n13325);
  not g24132 (n_12806, n13328);
  and g24133 (n13329, n_12805, n_12806);
  not g24134 (n_12807, n13307);
  and g24135 (n13330, n_12807, n13329);
  not g24136 (n_12808, n13329);
  and g24137 (n13331, n13307, n_12808);
  not g24138 (n_12809, n13330);
  not g24139 (n_12810, n13331);
  and g24140 (n13332, n_12809, n_12810);
  and g24141 (n13333, n13293, n13332);
  not g24142 (n_12811, n13293);
  not g24143 (n_12812, n13332);
  and g24144 (n13334, n_12811, n_12812);
  and g24145 (n13335, n_12191, n_12192);
  not g24146 (n_12813, n13335);
  and g24147 (n13336, n_12195, n_12813);
  not g24151 (n_12814, n13336);
  not g24152 (n_12815, n13339);
  and g24153 (n13340, n_12814, n_12815);
  and g24154 (n13341, n12547, n12552);
  not g24155 (n_12816, n13341);
  and g24156 (n13342, n_12170, n_12816);
  and g24157 (n13343, n_12166, n_12167);
  not g24158 (n_12817, n13342);
  not g24159 (n_12818, n13343);
  and g24160 (n13344, n_12817, n_12818);
  and g24161 (n13345, n12571, n12576);
  not g24162 (n_12819, n13345);
  and g24163 (n13346, n_12187, n_12819);
  and g24164 (n13347, n_12183, n_12184);
  not g24165 (n_12820, n13346);
  not g24166 (n_12821, n13347);
  and g24167 (n13348, n_12820, n_12821);
  not g24168 (n_12822, n13344);
  and g24169 (n13349, n_12822, n13348);
  not g24170 (n_12823, n13348);
  and g24171 (n13350, n13344, n_12823);
  not g24172 (n_12824, n13349);
  not g24173 (n_12825, n13350);
  and g24174 (n13351, n_12824, n_12825);
  not g24175 (n_12826, n13340);
  not g24176 (n_12827, n13351);
  and g24177 (n13352, n_12826, n_12827);
  not g24181 (n_12828, n13352);
  not g24182 (n_12829, n13355);
  and g24183 (n13356, n_12828, n_12829);
  not g24184 (n_12830, n13334);
  not g24185 (n_12831, n13356);
  and g24186 (n13357, n_12830, n_12831);
  not g24187 (n_12832, n13333);
  and g24188 (n13358, n_12832, n13357);
  and g24189 (n13359, n_12832, n_12830);
  not g24190 (n_12833, n13359);
  and g24191 (n13360, n13356, n_12833);
  not g24192 (n_12834, n13358);
  not g24193 (n_12835, n13360);
  and g24194 (n13361, n_12834, n_12835);
  and g24195 (n13362, n13289, n13361);
  not g24196 (n_12836, n13289);
  not g24197 (n_12837, n13361);
  and g24198 (n13363, n_12836, n_12837);
  and g24199 (n13364, n_12300, n_12301);
  not g24200 (n_12838, n13364);
  and g24201 (n13365, n_12304, n_12838);
  and g24202 (n13366, n12659, n12717);
  not g24203 (n_12839, n13365);
  not g24204 (n_12840, n13366);
  and g24205 (n13367, n_12839, n_12840);
  and g24206 (n13368, n_12292, n_12293);
  not g24207 (n_12841, n13368);
  and g24208 (n13369, n_12296, n_12841);
  not g24212 (n_12842, n13369);
  not g24213 (n_12843, n13372);
  and g24214 (n13373, n_12842, n_12843);
  and g24215 (n13374, n12674, n12679);
  not g24216 (n_12844, n13374);
  and g24217 (n13375, n_12271, n_12844);
  and g24218 (n13376, n_12267, n_12268);
  not g24219 (n_12845, n13375);
  not g24220 (n_12846, n13376);
  and g24221 (n13377, n_12845, n_12846);
  and g24222 (n13378, n12698, n12703);
  not g24223 (n_12847, n13378);
  and g24224 (n13379, n_12288, n_12847);
  and g24225 (n13380, n_12284, n_12285);
  not g24226 (n_12848, n13379);
  not g24227 (n_12849, n13380);
  and g24228 (n13381, n_12848, n_12849);
  not g24229 (n_12850, n13377);
  and g24230 (n13382, n_12850, n13381);
  not g24231 (n_12851, n13381);
  and g24232 (n13383, n13377, n_12851);
  not g24233 (n_12852, n13382);
  not g24234 (n_12853, n13383);
  and g24235 (n13384, n_12852, n_12853);
  not g24236 (n_12854, n13373);
  not g24237 (n_12855, n13384);
  and g24238 (n13385, n_12854, n_12855);
  not g24242 (n_12856, n13385);
  not g24243 (n_12857, n13388);
  and g24244 (n13389, n_12856, n_12857);
  and g24245 (n13390, n_12247, n_12248);
  not g24246 (n_12858, n13390);
  and g24247 (n13391, n_12251, n_12858);
  not g24251 (n_12859, n13391);
  not g24252 (n_12860, n13394);
  and g24253 (n13395, n_12859, n_12860);
  and g24254 (n13396, n12616, n12621);
  not g24255 (n_12861, n13396);
  and g24256 (n13397, n_12226, n_12861);
  and g24257 (n13398, n_12222, n_12223);
  not g24258 (n_12862, n13397);
  not g24259 (n_12863, n13398);
  and g24260 (n13399, n_12862, n_12863);
  and g24261 (n13400, n12640, n12645);
  not g24262 (n_12864, n13400);
  and g24263 (n13401, n_12243, n_12864);
  and g24264 (n13402, n_12239, n_12240);
  not g24265 (n_12865, n13401);
  not g24266 (n_12866, n13402);
  and g24267 (n13403, n_12865, n_12866);
  not g24268 (n_12867, n13399);
  and g24269 (n13404, n_12867, n13403);
  not g24270 (n_12868, n13403);
  and g24271 (n13405, n13399, n_12868);
  not g24272 (n_12869, n13404);
  not g24273 (n_12870, n13405);
  and g24274 (n13406, n_12869, n_12870);
  not g24275 (n_12871, n13395);
  not g24276 (n_12872, n13406);
  and g24277 (n13407, n_12871, n_12872);
  not g24281 (n_12873, n13407);
  not g24282 (n_12874, n13410);
  and g24283 (n13411, n_12873, n_12874);
  not g24284 (n_12875, n13389);
  and g24285 (n13412, n_12875, n13411);
  not g24286 (n_12876, n13411);
  and g24287 (n13413, n13389, n_12876);
  not g24288 (n_12877, n13412);
  not g24289 (n_12878, n13413);
  and g24290 (n13414, n_12877, n_12878);
  not g24291 (n_12879, n13367);
  not g24292 (n_12880, n13414);
  and g24293 (n13415, n_12879, n_12880);
  and g24294 (n13416, n13367, n13414);
  not g24295 (n_12881, n13415);
  not g24296 (n_12882, n13416);
  and g24297 (n13417, n_12881, n_12882);
  not g24298 (n_12883, n13363);
  not g24299 (n_12884, n13417);
  and g24300 (n13418, n_12883, n_12884);
  not g24301 (n_12885, n13362);
  and g24302 (n13419, n_12885, n13418);
  and g24303 (n13420, n_12885, n_12883);
  not g24304 (n_12886, n13420);
  and g24305 (n13421, n13417, n_12886);
  not g24306 (n_12887, n13419);
  not g24307 (n_12888, n13421);
  and g24308 (n13422, n_12887, n_12888);
  not g24309 (n_12889, n13284);
  not g24310 (n_12890, n13422);
  and g24311 (n13423, n_12889, n_12890);
  and g24312 (n13424, n13284, n13422);
  not g24313 (n_12891, n13423);
  not g24314 (n_12892, n13424);
  and g24315 (n13425, n_12891, n_12892);
  and g24316 (n13426, n_12049, n_12050);
  not g24317 (n_12893, n13426);
  and g24318 (n13427, n_12053, n_12893);
  and g24319 (n13428, n12141, n12403);
  not g24320 (n_12894, n13427);
  not g24321 (n_12895, n13428);
  and g24322 (n13429, n_12894, n_12895);
  and g24323 (n13430, n_12041, n_12042);
  not g24324 (n_12896, n13430);
  and g24325 (n13431, n_12045, n_12896);
  and g24326 (n13432, n12271, n12397);
  not g24327 (n_12897, n13431);
  not g24328 (n_12898, n13432);
  and g24329 (n13433, n_12897, n_12898);
  and g24330 (n13434, n_12033, n_12034);
  not g24331 (n_12899, n13434);
  and g24332 (n13435, n_12037, n_12899);
  and g24333 (n13436, n12333, n12391);
  not g24334 (n_12900, n13435);
  not g24335 (n_12901, n13436);
  and g24336 (n13437, n_12900, n_12901);
  and g24337 (n13438, n_12025, n_12026);
  not g24338 (n_12902, n13438);
  and g24339 (n13439, n_12029, n_12902);
  not g24343 (n_12903, n13439);
  not g24344 (n_12904, n13442);
  and g24345 (n13443, n_12903, n_12904);
  and g24346 (n13444, n12348, n12353);
  not g24347 (n_12905, n13444);
  and g24348 (n13445, n_12004, n_12905);
  and g24349 (n13446, n_12000, n_12001);
  not g24350 (n_12906, n13445);
  not g24351 (n_12907, n13446);
  and g24352 (n13447, n_12906, n_12907);
  and g24353 (n13448, n12372, n12377);
  not g24354 (n_12908, n13448);
  and g24355 (n13449, n_12021, n_12908);
  and g24356 (n13450, n_12017, n_12018);
  not g24357 (n_12909, n13449);
  not g24358 (n_12910, n13450);
  and g24359 (n13451, n_12909, n_12910);
  not g24360 (n_12911, n13447);
  and g24361 (n13452, n_12911, n13451);
  not g24362 (n_12912, n13451);
  and g24363 (n13453, n13447, n_12912);
  not g24364 (n_12913, n13452);
  not g24365 (n_12914, n13453);
  and g24366 (n13454, n_12913, n_12914);
  not g24367 (n_12915, n13443);
  not g24368 (n_12916, n13454);
  and g24369 (n13455, n_12915, n_12916);
  not g24373 (n_12917, n13455);
  not g24374 (n_12918, n13458);
  and g24375 (n13459, n_12917, n_12918);
  and g24376 (n13460, n_11980, n_11981);
  not g24377 (n_12919, n13460);
  and g24378 (n13461, n_11984, n_12919);
  not g24382 (n_12920, n13461);
  not g24383 (n_12921, n13464);
  and g24384 (n13465, n_12920, n_12921);
  and g24385 (n13466, n12290, n12295);
  not g24386 (n_12922, n13466);
  and g24387 (n13467, n_11959, n_12922);
  and g24388 (n13468, n_11955, n_11956);
  not g24389 (n_12923, n13467);
  not g24390 (n_12924, n13468);
  and g24391 (n13469, n_12923, n_12924);
  and g24392 (n13470, n12314, n12319);
  not g24393 (n_12925, n13470);
  and g24394 (n13471, n_11976, n_12925);
  and g24395 (n13472, n_11972, n_11973);
  not g24396 (n_12926, n13471);
  not g24397 (n_12927, n13472);
  and g24398 (n13473, n_12926, n_12927);
  not g24399 (n_12928, n13469);
  and g24400 (n13474, n_12928, n13473);
  not g24401 (n_12929, n13473);
  and g24402 (n13475, n13469, n_12929);
  not g24403 (n_12930, n13474);
  not g24404 (n_12931, n13475);
  and g24405 (n13476, n_12930, n_12931);
  not g24406 (n_12932, n13465);
  not g24407 (n_12933, n13476);
  and g24408 (n13477, n_12932, n_12933);
  not g24412 (n_12934, n13477);
  not g24413 (n_12935, n13480);
  and g24414 (n13481, n_12934, n_12935);
  not g24415 (n_12936, n13459);
  and g24416 (n13482, n_12936, n13481);
  not g24417 (n_12937, n13481);
  and g24418 (n13483, n13459, n_12937);
  not g24419 (n_12938, n13482);
  not g24420 (n_12939, n13483);
  and g24421 (n13484, n_12938, n_12939);
  not g24422 (n_12940, n13437);
  not g24423 (n_12941, n13484);
  and g24424 (n13485, n_12940, n_12941);
  and g24425 (n13486, n13437, n13484);
  not g24426 (n_12942, n13485);
  not g24427 (n_12943, n13486);
  and g24428 (n13487, n_12942, n_12943);
  and g24429 (n13488, n_11932, n_11933);
  not g24430 (n_12944, n13488);
  and g24431 (n13489, n_11936, n_12944);
  and g24432 (n13490, n12207, n12265);
  not g24433 (n_12945, n13489);
  not g24434 (n_12946, n13490);
  and g24435 (n13491, n_12945, n_12946);
  and g24436 (n13492, n_11924, n_11925);
  not g24437 (n_12947, n13492);
  and g24438 (n13493, n_11928, n_12947);
  not g24442 (n_12948, n13493);
  not g24443 (n_12949, n13496);
  and g24444 (n13497, n_12948, n_12949);
  and g24445 (n13498, n12222, n12227);
  not g24446 (n_12950, n13498);
  and g24447 (n13499, n_11903, n_12950);
  and g24448 (n13500, n_11899, n_11900);
  not g24449 (n_12951, n13499);
  not g24450 (n_12952, n13500);
  and g24451 (n13501, n_12951, n_12952);
  and g24452 (n13502, n12246, n12251);
  not g24453 (n_12953, n13502);
  and g24454 (n13503, n_11920, n_12953);
  and g24455 (n13504, n_11916, n_11917);
  not g24456 (n_12954, n13503);
  not g24457 (n_12955, n13504);
  and g24458 (n13505, n_12954, n_12955);
  not g24459 (n_12956, n13501);
  and g24460 (n13506, n_12956, n13505);
  not g24461 (n_12957, n13505);
  and g24462 (n13507, n13501, n_12957);
  not g24463 (n_12958, n13506);
  not g24464 (n_12959, n13507);
  and g24465 (n13508, n_12958, n_12959);
  not g24466 (n_12960, n13497);
  not g24467 (n_12961, n13508);
  and g24468 (n13509, n_12960, n_12961);
  not g24472 (n_12962, n13509);
  not g24473 (n_12963, n13512);
  and g24474 (n13513, n_12962, n_12963);
  and g24475 (n13514, n_11879, n_11880);
  not g24476 (n_12964, n13514);
  and g24477 (n13515, n_11883, n_12964);
  not g24481 (n_12965, n13515);
  not g24482 (n_12966, n13518);
  and g24483 (n13519, n_12965, n_12966);
  and g24484 (n13520, n12164, n12169);
  not g24485 (n_12967, n13520);
  and g24486 (n13521, n_11858, n_12967);
  and g24487 (n13522, n_11854, n_11855);
  not g24488 (n_12968, n13521);
  not g24489 (n_12969, n13522);
  and g24490 (n13523, n_12968, n_12969);
  and g24491 (n13524, n12188, n12193);
  not g24492 (n_12970, n13524);
  and g24493 (n13525, n_11875, n_12970);
  and g24494 (n13526, n_11871, n_11872);
  not g24495 (n_12971, n13525);
  not g24496 (n_12972, n13526);
  and g24497 (n13527, n_12971, n_12972);
  not g24498 (n_12973, n13523);
  and g24499 (n13528, n_12973, n13527);
  not g24500 (n_12974, n13527);
  and g24501 (n13529, n13523, n_12974);
  not g24502 (n_12975, n13528);
  not g24503 (n_12976, n13529);
  and g24504 (n13530, n_12975, n_12976);
  not g24505 (n_12977, n13519);
  not g24506 (n_12978, n13530);
  and g24507 (n13531, n_12977, n_12978);
  not g24511 (n_12979, n13531);
  not g24512 (n_12980, n13534);
  and g24513 (n13535, n_12979, n_12980);
  not g24514 (n_12981, n13513);
  and g24515 (n13536, n_12981, n13535);
  not g24516 (n_12982, n13535);
  and g24517 (n13537, n13513, n_12982);
  not g24518 (n_12983, n13536);
  not g24519 (n_12984, n13537);
  and g24520 (n13538, n_12983, n_12984);
  not g24521 (n_12985, n13491);
  not g24522 (n_12986, n13538);
  and g24523 (n13539, n_12985, n_12986);
  and g24524 (n13540, n13491, n13538);
  not g24525 (n_12987, n13539);
  not g24526 (n_12988, n13540);
  and g24527 (n13541, n_12987, n_12988);
  not g24528 (n_12989, n13487);
  and g24529 (n13542, n_12989, n13541);
  not g24530 (n_12990, n13541);
  and g24531 (n13543, n13487, n_12990);
  not g24532 (n_12991, n13542);
  not g24533 (n_12992, n13543);
  and g24534 (n13544, n_12991, n_12992);
  not g24535 (n_12993, n13433);
  not g24536 (n_12994, n13544);
  and g24537 (n13545, n_12993, n_12994);
  and g24538 (n13546, n13433, n13544);
  not g24539 (n_12995, n13545);
  not g24540 (n_12996, n13546);
  and g24541 (n13547, n_12995, n_12996);
  and g24542 (n13548, n_11828, n_11829);
  not g24543 (n_12997, n13548);
  and g24544 (n13549, n_11832, n_12997);
  and g24545 (n13550, n12009, n12135);
  not g24546 (n_12998, n13549);
  not g24547 (n_12999, n13550);
  and g24548 (n13551, n_12998, n_12999);
  and g24549 (n13552, n_11820, n_11821);
  not g24550 (n_13000, n13552);
  and g24551 (n13553, n_11824, n_13000);
  and g24552 (n13554, n12071, n12129);
  not g24553 (n_13001, n13553);
  not g24554 (n_13002, n13554);
  and g24555 (n13555, n_13001, n_13002);
  and g24556 (n13556, n_11812, n_11813);
  not g24557 (n_13003, n13556);
  and g24558 (n13557, n_11816, n_13003);
  not g24562 (n_13004, n13557);
  not g24563 (n_13005, n13560);
  and g24564 (n13561, n_13004, n_13005);
  and g24565 (n13562, n12086, n12091);
  not g24566 (n_13006, n13562);
  and g24567 (n13563, n_11791, n_13006);
  and g24568 (n13564, n_11787, n_11788);
  not g24569 (n_13007, n13563);
  not g24570 (n_13008, n13564);
  and g24571 (n13565, n_13007, n_13008);
  and g24572 (n13566, n12110, n12115);
  not g24573 (n_13009, n13566);
  and g24574 (n13567, n_11808, n_13009);
  and g24575 (n13568, n_11804, n_11805);
  not g24576 (n_13010, n13567);
  not g24577 (n_13011, n13568);
  and g24578 (n13569, n_13010, n_13011);
  not g24579 (n_13012, n13565);
  and g24580 (n13570, n_13012, n13569);
  not g24581 (n_13013, n13569);
  and g24582 (n13571, n13565, n_13013);
  not g24583 (n_13014, n13570);
  not g24584 (n_13015, n13571);
  and g24585 (n13572, n_13014, n_13015);
  not g24586 (n_13016, n13561);
  not g24587 (n_13017, n13572);
  and g24588 (n13573, n_13016, n_13017);
  not g24592 (n_13018, n13573);
  not g24593 (n_13019, n13576);
  and g24594 (n13577, n_13018, n_13019);
  and g24595 (n13578, n_11767, n_11768);
  not g24596 (n_13020, n13578);
  and g24597 (n13579, n_11771, n_13020);
  not g24601 (n_13021, n13579);
  not g24602 (n_13022, n13582);
  and g24603 (n13583, n_13021, n_13022);
  and g24604 (n13584, n12028, n12033);
  not g24605 (n_13023, n13584);
  and g24606 (n13585, n_11746, n_13023);
  and g24607 (n13586, n_11742, n_11743);
  not g24608 (n_13024, n13585);
  not g24609 (n_13025, n13586);
  and g24610 (n13587, n_13024, n_13025);
  and g24611 (n13588, n12052, n12057);
  not g24612 (n_13026, n13588);
  and g24613 (n13589, n_11763, n_13026);
  and g24614 (n13590, n_11759, n_11760);
  not g24615 (n_13027, n13589);
  not g24616 (n_13028, n13590);
  and g24617 (n13591, n_13027, n_13028);
  not g24618 (n_13029, n13587);
  and g24619 (n13592, n_13029, n13591);
  not g24620 (n_13030, n13591);
  and g24621 (n13593, n13587, n_13030);
  not g24622 (n_13031, n13592);
  not g24623 (n_13032, n13593);
  and g24624 (n13594, n_13031, n_13032);
  not g24625 (n_13033, n13583);
  not g24626 (n_13034, n13594);
  and g24627 (n13595, n_13033, n_13034);
  not g24631 (n_13035, n13595);
  not g24632 (n_13036, n13598);
  and g24633 (n13599, n_13035, n_13036);
  not g24634 (n_13037, n13577);
  and g24635 (n13600, n_13037, n13599);
  not g24636 (n_13038, n13599);
  and g24637 (n13601, n13577, n_13038);
  not g24638 (n_13039, n13600);
  not g24639 (n_13040, n13601);
  and g24640 (n13602, n_13039, n_13040);
  not g24641 (n_13041, n13555);
  not g24642 (n_13042, n13602);
  and g24643 (n13603, n_13041, n_13042);
  and g24644 (n13604, n13555, n13602);
  not g24645 (n_13043, n13603);
  not g24646 (n_13044, n13604);
  and g24647 (n13605, n_13043, n_13044);
  and g24648 (n13606, n_11719, n_11720);
  not g24649 (n_13045, n13606);
  and g24650 (n13607, n_11723, n_13045);
  and g24651 (n13608, n11945, n12003);
  not g24652 (n_13046, n13607);
  not g24653 (n_13047, n13608);
  and g24654 (n13609, n_13046, n_13047);
  and g24655 (n13610, n_11711, n_11712);
  not g24656 (n_13048, n13610);
  and g24657 (n13611, n_11715, n_13048);
  not g24661 (n_13049, n13611);
  not g24662 (n_13050, n13614);
  and g24663 (n13615, n_13049, n_13050);
  and g24664 (n13616, n11960, n11965);
  not g24665 (n_13051, n13616);
  and g24666 (n13617, n_11690, n_13051);
  and g24667 (n13618, n_11686, n_11687);
  not g24668 (n_13052, n13617);
  not g24669 (n_13053, n13618);
  and g24670 (n13619, n_13052, n_13053);
  and g24671 (n13620, n11984, n11989);
  not g24672 (n_13054, n13620);
  and g24673 (n13621, n_11707, n_13054);
  and g24674 (n13622, n_11703, n_11704);
  not g24675 (n_13055, n13621);
  not g24676 (n_13056, n13622);
  and g24677 (n13623, n_13055, n_13056);
  not g24678 (n_13057, n13619);
  and g24679 (n13624, n_13057, n13623);
  not g24680 (n_13058, n13623);
  and g24681 (n13625, n13619, n_13058);
  not g24682 (n_13059, n13624);
  not g24683 (n_13060, n13625);
  and g24684 (n13626, n_13059, n_13060);
  not g24685 (n_13061, n13615);
  not g24686 (n_13062, n13626);
  and g24687 (n13627, n_13061, n_13062);
  not g24691 (n_13063, n13627);
  not g24692 (n_13064, n13630);
  and g24693 (n13631, n_13063, n_13064);
  and g24694 (n13632, n_11666, n_11667);
  not g24695 (n_13065, n13632);
  and g24696 (n13633, n_11670, n_13065);
  not g24700 (n_13066, n13633);
  not g24701 (n_13067, n13636);
  and g24702 (n13637, n_13066, n_13067);
  and g24703 (n13638, n11902, n11907);
  not g24704 (n_13068, n13638);
  and g24705 (n13639, n_11645, n_13068);
  and g24706 (n13640, n_11641, n_11642);
  not g24707 (n_13069, n13639);
  not g24708 (n_13070, n13640);
  and g24709 (n13641, n_13069, n_13070);
  and g24710 (n13642, n11926, n11931);
  not g24711 (n_13071, n13642);
  and g24712 (n13643, n_11662, n_13071);
  and g24713 (n13644, n_11658, n_11659);
  not g24714 (n_13072, n13643);
  not g24715 (n_13073, n13644);
  and g24716 (n13645, n_13072, n_13073);
  not g24717 (n_13074, n13641);
  and g24718 (n13646, n_13074, n13645);
  not g24719 (n_13075, n13645);
  and g24720 (n13647, n13641, n_13075);
  not g24721 (n_13076, n13646);
  not g24722 (n_13077, n13647);
  and g24723 (n13648, n_13076, n_13077);
  not g24724 (n_13078, n13637);
  not g24725 (n_13079, n13648);
  and g24726 (n13649, n_13078, n_13079);
  not g24730 (n_13080, n13649);
  not g24731 (n_13081, n13652);
  and g24732 (n13653, n_13080, n_13081);
  not g24733 (n_13082, n13631);
  and g24734 (n13654, n_13082, n13653);
  not g24735 (n_13083, n13653);
  and g24736 (n13655, n13631, n_13083);
  not g24737 (n_13084, n13654);
  not g24738 (n_13085, n13655);
  and g24739 (n13656, n_13084, n_13085);
  not g24740 (n_13086, n13609);
  not g24741 (n_13087, n13656);
  and g24742 (n13657, n_13086, n_13087);
  and g24743 (n13658, n13609, n13656);
  not g24744 (n_13088, n13657);
  not g24745 (n_13089, n13658);
  and g24746 (n13659, n_13088, n_13089);
  not g24747 (n_13090, n13605);
  and g24748 (n13660, n_13090, n13659);
  not g24749 (n_13091, n13659);
  and g24750 (n13661, n13605, n_13091);
  not g24751 (n_13092, n13660);
  not g24752 (n_13093, n13661);
  and g24753 (n13662, n_13092, n_13093);
  not g24754 (n_13094, n13551);
  not g24755 (n_13095, n13662);
  and g24756 (n13663, n_13094, n_13095);
  and g24757 (n13664, n13551, n13662);
  not g24758 (n_13096, n13663);
  not g24759 (n_13097, n13664);
  and g24760 (n13665, n_13096, n_13097);
  not g24761 (n_13098, n13547);
  and g24762 (n13666, n_13098, n13665);
  not g24763 (n_13099, n13665);
  and g24764 (n13667, n13547, n_13099);
  not g24765 (n_13100, n13666);
  not g24766 (n_13101, n13667);
  and g24767 (n13668, n_13100, n_13101);
  not g24768 (n_13102, n13429);
  not g24769 (n_13103, n13668);
  and g24770 (n13669, n_13102, n_13103);
  and g24771 (n13670, n13429, n13668);
  not g24772 (n_13104, n13669);
  not g24773 (n_13105, n13670);
  and g24774 (n13671, n_13104, n_13105);
  not g24775 (n_13106, n13425);
  and g24776 (n13672, n_13106, n13671);
  not g24777 (n_13107, n13671);
  and g24778 (n13673, n13425, n_13107);
  not g24779 (n_13108, n13672);
  not g24780 (n_13109, n13673);
  and g24781 (n13674, n_13108, n_13109);
  not g24782 (n_13110, n13279);
  not g24783 (n_13111, n13674);
  and g24784 (n13675, n_13110, n_13111);
  and g24785 (n13676, n13279, n13674);
  not g24786 (n_13112, n13675);
  not g24787 (n_13113, n13676);
  and g24788 (n13677, n_13112, n_13113);
  and g24789 (n13678, n_12753, n_12754);
  not g24790 (n_13114, n13678);
  and g24791 (n13679, n_12757, n_13114);
  and g24792 (n13680, n13002, n13264);
  not g24793 (n_13115, n13679);
  not g24794 (n_13116, n13680);
  and g24795 (n13681, n_13115, n_13116);
  and g24796 (n13682, n_12745, n_12746);
  not g24797 (n_13117, n13682);
  and g24798 (n13683, n_12749, n_13117);
  and g24799 (n13684, n13132, n13258);
  not g24800 (n_13118, n13683);
  not g24801 (n_13119, n13684);
  and g24802 (n13685, n_13118, n_13119);
  and g24803 (n13686, n_12737, n_12738);
  not g24804 (n_13120, n13686);
  and g24805 (n13687, n_12741, n_13120);
  and g24806 (n13688, n13194, n13252);
  not g24807 (n_13121, n13687);
  not g24808 (n_13122, n13688);
  and g24809 (n13689, n_13121, n_13122);
  and g24810 (n13690, n_12729, n_12730);
  not g24811 (n_13123, n13690);
  and g24812 (n13691, n_12733, n_13123);
  not g24816 (n_13124, n13691);
  not g24817 (n_13125, n13694);
  and g24818 (n13695, n_13124, n_13125);
  and g24819 (n13696, n13209, n13214);
  not g24820 (n_13126, n13696);
  and g24821 (n13697, n_12708, n_13126);
  and g24822 (n13698, n_12704, n_12705);
  not g24823 (n_13127, n13697);
  not g24824 (n_13128, n13698);
  and g24825 (n13699, n_13127, n_13128);
  and g24826 (n13700, n13233, n13238);
  not g24827 (n_13129, n13700);
  and g24828 (n13701, n_12725, n_13129);
  and g24829 (n13702, n_12721, n_12722);
  not g24830 (n_13130, n13701);
  not g24831 (n_13131, n13702);
  and g24832 (n13703, n_13130, n_13131);
  not g24833 (n_13132, n13699);
  and g24834 (n13704, n_13132, n13703);
  not g24835 (n_13133, n13703);
  and g24836 (n13705, n13699, n_13133);
  not g24837 (n_13134, n13704);
  not g24838 (n_13135, n13705);
  and g24839 (n13706, n_13134, n_13135);
  not g24840 (n_13136, n13695);
  not g24841 (n_13137, n13706);
  and g24842 (n13707, n_13136, n_13137);
  not g24846 (n_13138, n13707);
  not g24847 (n_13139, n13710);
  and g24848 (n13711, n_13138, n_13139);
  and g24849 (n13712, n_12684, n_12685);
  not g24850 (n_13140, n13712);
  and g24851 (n13713, n_12688, n_13140);
  not g24855 (n_13141, n13713);
  not g24856 (n_13142, n13716);
  and g24857 (n13717, n_13141, n_13142);
  and g24858 (n13718, n13151, n13156);
  not g24859 (n_13143, n13718);
  and g24860 (n13719, n_12663, n_13143);
  and g24861 (n13720, n_12659, n_12660);
  not g24862 (n_13144, n13719);
  not g24863 (n_13145, n13720);
  and g24864 (n13721, n_13144, n_13145);
  and g24865 (n13722, n13175, n13180);
  not g24866 (n_13146, n13722);
  and g24867 (n13723, n_12680, n_13146);
  and g24868 (n13724, n_12676, n_12677);
  not g24869 (n_13147, n13723);
  not g24870 (n_13148, n13724);
  and g24871 (n13725, n_13147, n_13148);
  not g24872 (n_13149, n13721);
  and g24873 (n13726, n_13149, n13725);
  not g24874 (n_13150, n13725);
  and g24875 (n13727, n13721, n_13150);
  not g24876 (n_13151, n13726);
  not g24877 (n_13152, n13727);
  and g24878 (n13728, n_13151, n_13152);
  not g24879 (n_13153, n13717);
  not g24880 (n_13154, n13728);
  and g24881 (n13729, n_13153, n_13154);
  not g24885 (n_13155, n13729);
  not g24886 (n_13156, n13732);
  and g24887 (n13733, n_13155, n_13156);
  not g24888 (n_13157, n13711);
  and g24889 (n13734, n_13157, n13733);
  not g24890 (n_13158, n13733);
  and g24891 (n13735, n13711, n_13158);
  not g24892 (n_13159, n13734);
  not g24893 (n_13160, n13735);
  and g24894 (n13736, n_13159, n_13160);
  not g24895 (n_13161, n13689);
  not g24896 (n_13162, n13736);
  and g24897 (n13737, n_13161, n_13162);
  and g24898 (n13738, n13689, n13736);
  not g24899 (n_13163, n13737);
  not g24900 (n_13164, n13738);
  and g24901 (n13739, n_13163, n_13164);
  and g24902 (n13740, n_12636, n_12637);
  not g24903 (n_13165, n13740);
  and g24904 (n13741, n_12640, n_13165);
  and g24905 (n13742, n13068, n13126);
  not g24906 (n_13166, n13741);
  not g24907 (n_13167, n13742);
  and g24908 (n13743, n_13166, n_13167);
  and g24909 (n13744, n_12628, n_12629);
  not g24910 (n_13168, n13744);
  and g24911 (n13745, n_12632, n_13168);
  not g24915 (n_13169, n13745);
  not g24916 (n_13170, n13748);
  and g24917 (n13749, n_13169, n_13170);
  and g24918 (n13750, n13083, n13088);
  not g24919 (n_13171, n13750);
  and g24920 (n13751, n_12607, n_13171);
  and g24921 (n13752, n_12603, n_12604);
  not g24922 (n_13172, n13751);
  not g24923 (n_13173, n13752);
  and g24924 (n13753, n_13172, n_13173);
  and g24925 (n13754, n13107, n13112);
  not g24926 (n_13174, n13754);
  and g24927 (n13755, n_12624, n_13174);
  and g24928 (n13756, n_12620, n_12621);
  not g24929 (n_13175, n13755);
  not g24930 (n_13176, n13756);
  and g24931 (n13757, n_13175, n_13176);
  not g24932 (n_13177, n13753);
  and g24933 (n13758, n_13177, n13757);
  not g24934 (n_13178, n13757);
  and g24935 (n13759, n13753, n_13178);
  not g24936 (n_13179, n13758);
  not g24937 (n_13180, n13759);
  and g24938 (n13760, n_13179, n_13180);
  not g24939 (n_13181, n13749);
  not g24940 (n_13182, n13760);
  and g24941 (n13761, n_13181, n_13182);
  not g24945 (n_13183, n13761);
  not g24946 (n_13184, n13764);
  and g24947 (n13765, n_13183, n_13184);
  and g24948 (n13766, n_12583, n_12584);
  not g24949 (n_13185, n13766);
  and g24950 (n13767, n_12587, n_13185);
  not g24954 (n_13186, n13767);
  not g24955 (n_13187, n13770);
  and g24956 (n13771, n_13186, n_13187);
  and g24957 (n13772, n13025, n13030);
  not g24958 (n_13188, n13772);
  and g24959 (n13773, n_12562, n_13188);
  and g24960 (n13774, n_12558, n_12559);
  not g24961 (n_13189, n13773);
  not g24962 (n_13190, n13774);
  and g24963 (n13775, n_13189, n_13190);
  and g24964 (n13776, n13049, n13054);
  not g24965 (n_13191, n13776);
  and g24966 (n13777, n_12579, n_13191);
  and g24967 (n13778, n_12575, n_12576);
  not g24968 (n_13192, n13777);
  not g24969 (n_13193, n13778);
  and g24970 (n13779, n_13192, n_13193);
  not g24971 (n_13194, n13775);
  and g24972 (n13780, n_13194, n13779);
  not g24973 (n_13195, n13779);
  and g24974 (n13781, n13775, n_13195);
  not g24975 (n_13196, n13780);
  not g24976 (n_13197, n13781);
  and g24977 (n13782, n_13196, n_13197);
  not g24978 (n_13198, n13771);
  not g24979 (n_13199, n13782);
  and g24980 (n13783, n_13198, n_13199);
  not g24984 (n_13200, n13783);
  not g24985 (n_13201, n13786);
  and g24986 (n13787, n_13200, n_13201);
  not g24987 (n_13202, n13765);
  and g24988 (n13788, n_13202, n13787);
  not g24989 (n_13203, n13787);
  and g24990 (n13789, n13765, n_13203);
  not g24991 (n_13204, n13788);
  not g24992 (n_13205, n13789);
  and g24993 (n13790, n_13204, n_13205);
  not g24994 (n_13206, n13743);
  not g24995 (n_13207, n13790);
  and g24996 (n13791, n_13206, n_13207);
  and g24997 (n13792, n13743, n13790);
  not g24998 (n_13208, n13791);
  not g24999 (n_13209, n13792);
  and g25000 (n13793, n_13208, n_13209);
  not g25001 (n_13210, n13739);
  and g25002 (n13794, n_13210, n13793);
  not g25003 (n_13211, n13793);
  and g25004 (n13795, n13739, n_13211);
  not g25005 (n_13212, n13794);
  not g25006 (n_13213, n13795);
  and g25007 (n13796, n_13212, n_13213);
  not g25008 (n_13214, n13685);
  not g25009 (n_13215, n13796);
  and g25010 (n13797, n_13214, n_13215);
  and g25011 (n13798, n13685, n13796);
  not g25012 (n_13216, n13797);
  not g25013 (n_13217, n13798);
  and g25014 (n13799, n_13216, n_13217);
  and g25015 (n13800, n_12532, n_12533);
  not g25016 (n_13218, n13800);
  and g25017 (n13801, n_12536, n_13218);
  and g25018 (n13802, n12870, n12996);
  not g25019 (n_13219, n13801);
  not g25020 (n_13220, n13802);
  and g25021 (n13803, n_13219, n_13220);
  and g25022 (n13804, n_12524, n_12525);
  not g25023 (n_13221, n13804);
  and g25024 (n13805, n_12528, n_13221);
  and g25025 (n13806, n12932, n12990);
  not g25026 (n_13222, n13805);
  not g25027 (n_13223, n13806);
  and g25028 (n13807, n_13222, n_13223);
  and g25029 (n13808, n_12516, n_12517);
  not g25030 (n_13224, n13808);
  and g25031 (n13809, n_12520, n_13224);
  not g25035 (n_13225, n13809);
  not g25036 (n_13226, n13812);
  and g25037 (n13813, n_13225, n_13226);
  and g25038 (n13814, n12947, n12952);
  not g25039 (n_13227, n13814);
  and g25040 (n13815, n_12495, n_13227);
  and g25041 (n13816, n_12491, n_12492);
  not g25042 (n_13228, n13815);
  not g25043 (n_13229, n13816);
  and g25044 (n13817, n_13228, n_13229);
  and g25045 (n13818, n12971, n12976);
  not g25046 (n_13230, n13818);
  and g25047 (n13819, n_12512, n_13230);
  and g25048 (n13820, n_12508, n_12509);
  not g25049 (n_13231, n13819);
  not g25050 (n_13232, n13820);
  and g25051 (n13821, n_13231, n_13232);
  not g25052 (n_13233, n13817);
  and g25053 (n13822, n_13233, n13821);
  not g25054 (n_13234, n13821);
  and g25055 (n13823, n13817, n_13234);
  not g25056 (n_13235, n13822);
  not g25057 (n_13236, n13823);
  and g25058 (n13824, n_13235, n_13236);
  not g25059 (n_13237, n13813);
  not g25060 (n_13238, n13824);
  and g25061 (n13825, n_13237, n_13238);
  not g25065 (n_13239, n13825);
  not g25066 (n_13240, n13828);
  and g25067 (n13829, n_13239, n_13240);
  and g25068 (n13830, n_12471, n_12472);
  not g25069 (n_13241, n13830);
  and g25070 (n13831, n_12475, n_13241);
  not g25074 (n_13242, n13831);
  not g25075 (n_13243, n13834);
  and g25076 (n13835, n_13242, n_13243);
  and g25077 (n13836, n12889, n12894);
  not g25078 (n_13244, n13836);
  and g25079 (n13837, n_12450, n_13244);
  and g25080 (n13838, n_12446, n_12447);
  not g25081 (n_13245, n13837);
  not g25082 (n_13246, n13838);
  and g25083 (n13839, n_13245, n_13246);
  and g25084 (n13840, n12913, n12918);
  not g25085 (n_13247, n13840);
  and g25086 (n13841, n_12467, n_13247);
  and g25087 (n13842, n_12463, n_12464);
  not g25088 (n_13248, n13841);
  not g25089 (n_13249, n13842);
  and g25090 (n13843, n_13248, n_13249);
  not g25091 (n_13250, n13839);
  and g25092 (n13844, n_13250, n13843);
  not g25093 (n_13251, n13843);
  and g25094 (n13845, n13839, n_13251);
  not g25095 (n_13252, n13844);
  not g25096 (n_13253, n13845);
  and g25097 (n13846, n_13252, n_13253);
  not g25098 (n_13254, n13835);
  not g25099 (n_13255, n13846);
  and g25100 (n13847, n_13254, n_13255);
  not g25104 (n_13256, n13847);
  not g25105 (n_13257, n13850);
  and g25106 (n13851, n_13256, n_13257);
  not g25107 (n_13258, n13829);
  and g25108 (n13852, n_13258, n13851);
  not g25109 (n_13259, n13851);
  and g25110 (n13853, n13829, n_13259);
  not g25111 (n_13260, n13852);
  not g25112 (n_13261, n13853);
  and g25113 (n13854, n_13260, n_13261);
  not g25114 (n_13262, n13807);
  not g25115 (n_13263, n13854);
  and g25116 (n13855, n_13262, n_13263);
  and g25117 (n13856, n13807, n13854);
  not g25118 (n_13264, n13855);
  not g25119 (n_13265, n13856);
  and g25120 (n13857, n_13264, n_13265);
  and g25121 (n13858, n_12423, n_12424);
  not g25122 (n_13266, n13858);
  and g25123 (n13859, n_12427, n_13266);
  and g25124 (n13860, n12806, n12864);
  not g25125 (n_13267, n13859);
  not g25126 (n_13268, n13860);
  and g25127 (n13861, n_13267, n_13268);
  and g25128 (n13862, n_12415, n_12416);
  not g25129 (n_13269, n13862);
  and g25130 (n13863, n_12419, n_13269);
  not g25134 (n_13270, n13863);
  not g25135 (n_13271, n13866);
  and g25136 (n13867, n_13270, n_13271);
  and g25137 (n13868, n12821, n12826);
  not g25138 (n_13272, n13868);
  and g25139 (n13869, n_12394, n_13272);
  and g25140 (n13870, n_12390, n_12391);
  not g25141 (n_13273, n13869);
  not g25142 (n_13274, n13870);
  and g25143 (n13871, n_13273, n_13274);
  and g25144 (n13872, n12845, n12850);
  not g25145 (n_13275, n13872);
  and g25146 (n13873, n_12411, n_13275);
  and g25147 (n13874, n_12407, n_12408);
  not g25148 (n_13276, n13873);
  not g25149 (n_13277, n13874);
  and g25150 (n13875, n_13276, n_13277);
  not g25151 (n_13278, n13871);
  and g25152 (n13876, n_13278, n13875);
  not g25153 (n_13279, n13875);
  and g25154 (n13877, n13871, n_13279);
  not g25155 (n_13280, n13876);
  not g25156 (n_13281, n13877);
  and g25157 (n13878, n_13280, n_13281);
  not g25158 (n_13282, n13867);
  not g25159 (n_13283, n13878);
  and g25160 (n13879, n_13282, n_13283);
  not g25164 (n_13284, n13879);
  not g25165 (n_13285, n13882);
  and g25166 (n13883, n_13284, n_13285);
  and g25167 (n13884, n_12370, n_12371);
  not g25168 (n_13286, n13884);
  and g25169 (n13885, n_12374, n_13286);
  not g25173 (n_13287, n13885);
  not g25174 (n_13288, n13888);
  and g25175 (n13889, n_13287, n_13288);
  and g25176 (n13890, n12763, n12768);
  not g25177 (n_13289, n13890);
  and g25178 (n13891, n_12349, n_13289);
  and g25179 (n13892, n_12345, n_12346);
  not g25180 (n_13290, n13891);
  not g25181 (n_13291, n13892);
  and g25182 (n13893, n_13290, n_13291);
  and g25183 (n13894, n12787, n12792);
  not g25184 (n_13292, n13894);
  and g25185 (n13895, n_12366, n_13292);
  and g25186 (n13896, n_12362, n_12363);
  not g25187 (n_13293, n13895);
  not g25188 (n_13294, n13896);
  and g25189 (n13897, n_13293, n_13294);
  not g25190 (n_13295, n13893);
  and g25191 (n13898, n_13295, n13897);
  not g25192 (n_13296, n13897);
  and g25193 (n13899, n13893, n_13296);
  not g25194 (n_13297, n13898);
  not g25195 (n_13298, n13899);
  and g25196 (n13900, n_13297, n_13298);
  not g25197 (n_13299, n13889);
  not g25198 (n_13300, n13900);
  and g25199 (n13901, n_13299, n_13300);
  not g25203 (n_13301, n13901);
  not g25204 (n_13302, n13904);
  and g25205 (n13905, n_13301, n_13302);
  not g25206 (n_13303, n13883);
  and g25207 (n13906, n_13303, n13905);
  not g25208 (n_13304, n13905);
  and g25209 (n13907, n13883, n_13304);
  not g25210 (n_13305, n13906);
  not g25211 (n_13306, n13907);
  and g25212 (n13908, n_13305, n_13306);
  not g25213 (n_13307, n13861);
  not g25214 (n_13308, n13908);
  and g25215 (n13909, n_13307, n_13308);
  and g25216 (n13910, n13861, n13908);
  not g25217 (n_13309, n13909);
  not g25218 (n_13310, n13910);
  and g25219 (n13911, n_13309, n_13310);
  not g25220 (n_13311, n13857);
  and g25221 (n13912, n_13311, n13911);
  not g25222 (n_13312, n13911);
  and g25223 (n13913, n13857, n_13312);
  not g25224 (n_13313, n13912);
  not g25225 (n_13314, n13913);
  and g25226 (n13914, n_13313, n_13314);
  not g25227 (n_13315, n13803);
  not g25228 (n_13316, n13914);
  and g25229 (n13915, n_13315, n_13316);
  and g25230 (n13916, n13803, n13914);
  not g25231 (n_13317, n13915);
  not g25232 (n_13318, n13916);
  and g25233 (n13917, n_13317, n_13318);
  not g25234 (n_13319, n13799);
  and g25235 (n13918, n_13319, n13917);
  not g25236 (n_13320, n13917);
  and g25237 (n13919, n13799, n_13320);
  not g25238 (n_13321, n13918);
  not g25239 (n_13322, n13919);
  and g25240 (n13920, n_13321, n_13322);
  not g25241 (n_13323, n13681);
  not g25242 (n_13324, n13920);
  and g25243 (n13921, n_13323, n_13324);
  and g25244 (n13922, n13681, n13920);
  not g25245 (n_13325, n13921);
  not g25246 (n_13326, n13922);
  and g25247 (n13923, n_13325, n_13326);
  not g25248 (n_13327, n13677);
  not g25249 (n_13328, n13923);
  and g25250 (n13924, n_13327, n_13328);
  not g25251 (n_13329, n13275);
  not g25252 (n_13330, n13924);
  and g25253 (n13925, n_13329, n_13330);
  and g25254 (n13926, n_13112, n13923);
  and g25255 (n13927, n_13113, n13926);
  not g25256 (n_13331, n13925);
  not g25257 (n_13332, n13927);
  and g25258 (n13928, n_13331, n_13332);
  and g25259 (n13929, n_13106, n_13107);
  not g25260 (n_13333, n13929);
  and g25261 (n13930, n_13110, n_13333);
  and g25262 (n13931, n13425, n13671);
  not g25263 (n_13334, n13930);
  not g25264 (n_13335, n13931);
  and g25265 (n13932, n_13334, n_13335);
  and g25266 (n13933, n_13098, n_13099);
  not g25267 (n_13336, n13933);
  and g25268 (n13934, n_13102, n_13336);
  and g25269 (n13935, n13547, n13665);
  not g25270 (n_13337, n13934);
  not g25271 (n_13338, n13935);
  and g25272 (n13936, n_13337, n_13338);
  and g25273 (n13937, n_13090, n_13091);
  not g25274 (n_13339, n13937);
  and g25275 (n13938, n_13094, n_13339);
  and g25276 (n13939, n13605, n13659);
  not g25277 (n_13340, n13938);
  not g25278 (n_13341, n13939);
  and g25279 (n13940, n_13340, n_13341);
  and g25280 (n13941, n_13082, n_13083);
  not g25281 (n_13342, n13941);
  and g25282 (n13942, n_13086, n_13342);
  not g25286 (n_13343, n13942);
  not g25287 (n_13344, n13945);
  and g25288 (n13946, n_13343, n_13344);
  not g25292 (n_13345, n13949);
  and g25293 (n13950, n_13078, n_13345);
  and g25294 (n13951, n_13074, n_13075);
  not g25295 (n_13346, n13950);
  not g25296 (n_13347, n13951);
  and g25297 (n13952, n_13346, n_13347);
  not g25301 (n_13348, n13955);
  and g25302 (n13956, n_13061, n_13348);
  and g25303 (n13957, n_13057, n_13058);
  not g25304 (n_13349, n13956);
  not g25305 (n_13350, n13957);
  and g25306 (n13958, n_13349, n_13350);
  not g25307 (n_13351, n13952);
  and g25308 (n13959, n_13351, n13958);
  not g25309 (n_13352, n13958);
  and g25310 (n13960, n13952, n_13352);
  not g25311 (n_13353, n13959);
  not g25312 (n_13354, n13960);
  and g25313 (n13961, n_13353, n_13354);
  not g25314 (n_13355, n13946);
  not g25315 (n_13356, n13961);
  and g25316 (n13962, n_13355, n_13356);
  not g25320 (n_13357, n13962);
  not g25321 (n_13358, n13965);
  and g25322 (n13966, n_13357, n_13358);
  and g25323 (n13967, n_13037, n_13038);
  not g25324 (n_13359, n13967);
  and g25325 (n13968, n_13041, n_13359);
  not g25329 (n_13360, n13968);
  not g25330 (n_13361, n13971);
  and g25331 (n13972, n_13360, n_13361);
  not g25335 (n_13362, n13975);
  and g25336 (n13976, n_13033, n_13362);
  and g25337 (n13977, n_13029, n_13030);
  not g25338 (n_13363, n13976);
  not g25339 (n_13364, n13977);
  and g25340 (n13978, n_13363, n_13364);
  not g25344 (n_13365, n13981);
  and g25345 (n13982, n_13016, n_13365);
  and g25346 (n13983, n_13012, n_13013);
  not g25347 (n_13366, n13982);
  not g25348 (n_13367, n13983);
  and g25349 (n13984, n_13366, n_13367);
  not g25350 (n_13368, n13978);
  and g25351 (n13985, n_13368, n13984);
  not g25352 (n_13369, n13984);
  and g25353 (n13986, n13978, n_13369);
  not g25354 (n_13370, n13985);
  not g25355 (n_13371, n13986);
  and g25356 (n13987, n_13370, n_13371);
  not g25357 (n_13372, n13972);
  not g25358 (n_13373, n13987);
  and g25359 (n13988, n_13372, n_13373);
  not g25363 (n_13374, n13988);
  not g25364 (n_13375, n13991);
  and g25365 (n13992, n_13374, n_13375);
  not g25366 (n_13376, n13966);
  and g25367 (n13993, n_13376, n13992);
  not g25368 (n_13377, n13992);
  and g25369 (n13994, n13966, n_13377);
  not g25370 (n_13378, n13993);
  not g25371 (n_13379, n13994);
  and g25372 (n13995, n_13378, n_13379);
  not g25373 (n_13380, n13940);
  not g25374 (n_13381, n13995);
  and g25375 (n13996, n_13380, n_13381);
  and g25376 (n13997, n13940, n13995);
  not g25377 (n_13382, n13996);
  not g25378 (n_13383, n13997);
  and g25379 (n13998, n_13382, n_13383);
  and g25380 (n13999, n_12989, n_12990);
  not g25381 (n_13384, n13999);
  and g25382 (n14000, n_12993, n_13384);
  and g25383 (n14001, n13487, n13541);
  not g25384 (n_13385, n14000);
  not g25385 (n_13386, n14001);
  and g25386 (n14002, n_13385, n_13386);
  and g25387 (n14003, n_12981, n_12982);
  not g25388 (n_13387, n14003);
  and g25389 (n14004, n_12985, n_13387);
  not g25393 (n_13388, n14004);
  not g25394 (n_13389, n14007);
  and g25395 (n14008, n_13388, n_13389);
  not g25399 (n_13390, n14011);
  and g25400 (n14012, n_12977, n_13390);
  and g25401 (n14013, n_12973, n_12974);
  not g25402 (n_13391, n14012);
  not g25403 (n_13392, n14013);
  and g25404 (n14014, n_13391, n_13392);
  not g25408 (n_13393, n14017);
  and g25409 (n14018, n_12960, n_13393);
  and g25410 (n14019, n_12956, n_12957);
  not g25411 (n_13394, n14018);
  not g25412 (n_13395, n14019);
  and g25413 (n14020, n_13394, n_13395);
  not g25414 (n_13396, n14014);
  and g25415 (n14021, n_13396, n14020);
  not g25416 (n_13397, n14020);
  and g25417 (n14022, n14014, n_13397);
  not g25418 (n_13398, n14021);
  not g25419 (n_13399, n14022);
  and g25420 (n14023, n_13398, n_13399);
  not g25421 (n_13400, n14008);
  not g25422 (n_13401, n14023);
  and g25423 (n14024, n_13400, n_13401);
  not g25427 (n_13402, n14024);
  not g25428 (n_13403, n14027);
  and g25429 (n14028, n_13402, n_13403);
  and g25430 (n14029, n_12936, n_12937);
  not g25431 (n_13404, n14029);
  and g25432 (n14030, n_12940, n_13404);
  not g25436 (n_13405, n14030);
  not g25437 (n_13406, n14033);
  and g25438 (n14034, n_13405, n_13406);
  not g25442 (n_13407, n14037);
  and g25443 (n14038, n_12932, n_13407);
  and g25444 (n14039, n_12928, n_12929);
  not g25445 (n_13408, n14038);
  not g25446 (n_13409, n14039);
  and g25447 (n14040, n_13408, n_13409);
  not g25451 (n_13410, n14043);
  and g25452 (n14044, n_12915, n_13410);
  and g25453 (n14045, n_12911, n_12912);
  not g25454 (n_13411, n14044);
  not g25455 (n_13412, n14045);
  and g25456 (n14046, n_13411, n_13412);
  not g25457 (n_13413, n14040);
  and g25458 (n14047, n_13413, n14046);
  not g25459 (n_13414, n14046);
  and g25460 (n14048, n14040, n_13414);
  not g25461 (n_13415, n14047);
  not g25462 (n_13416, n14048);
  and g25463 (n14049, n_13415, n_13416);
  not g25464 (n_13417, n14034);
  not g25465 (n_13418, n14049);
  and g25466 (n14050, n_13417, n_13418);
  not g25470 (n_13419, n14050);
  not g25471 (n_13420, n14053);
  and g25472 (n14054, n_13419, n_13420);
  not g25473 (n_13421, n14028);
  and g25474 (n14055, n_13421, n14054);
  not g25475 (n_13422, n14054);
  and g25476 (n14056, n14028, n_13422);
  not g25477 (n_13423, n14055);
  not g25478 (n_13424, n14056);
  and g25479 (n14057, n_13423, n_13424);
  not g25480 (n_13425, n14002);
  not g25481 (n_13426, n14057);
  and g25482 (n14058, n_13425, n_13426);
  and g25483 (n14059, n14002, n14057);
  not g25484 (n_13427, n14058);
  not g25485 (n_13428, n14059);
  and g25486 (n14060, n_13427, n_13428);
  not g25487 (n_13429, n13998);
  and g25488 (n14061, n_13429, n14060);
  not g25489 (n_13430, n14060);
  and g25490 (n14062, n13998, n_13430);
  not g25491 (n_13431, n14061);
  not g25492 (n_13432, n14062);
  and g25493 (n14063, n_13431, n_13432);
  not g25494 (n_13433, n13936);
  not g25495 (n_13434, n14063);
  and g25496 (n14064, n_13433, n_13434);
  and g25497 (n14065, n13936, n14063);
  not g25498 (n_13435, n14064);
  not g25499 (n_13436, n14065);
  and g25500 (n14066, n_13435, n_13436);
  and g25501 (n14067, n_12884, n_12886);
  not g25502 (n_13437, n14067);
  and g25503 (n14068, n_12889, n_13437);
  and g25504 (n14069, n_12883, n13417);
  and g25505 (n14070, n_12885, n14069);
  not g25506 (n_13438, n14068);
  not g25507 (n_13439, n14070);
  and g25508 (n14071, n_13438, n_13439);
  and g25509 (n14072, n_12831, n_12833);
  not g25510 (n_13440, n14072);
  and g25511 (n14073, n_12836, n_13440);
  and g25512 (n14074, n_12830, n13356);
  and g25513 (n14075, n_12832, n14074);
  not g25514 (n_13441, n14073);
  not g25515 (n_13442, n14075);
  and g25516 (n14076, n_13441, n_13442);
  and g25517 (n14077, n_12807, n_12808);
  not g25518 (n_13443, n14077);
  and g25519 (n14078, n_12811, n_13443);
  not g25523 (n_13444, n14078);
  not g25524 (n_13445, n14081);
  and g25525 (n14082, n_13444, n_13445);
  not g25529 (n_13446, n14085);
  and g25530 (n14086, n_12803, n_13446);
  and g25531 (n14087, n_12799, n_12800);
  not g25532 (n_13447, n14086);
  not g25533 (n_13448, n14087);
  and g25534 (n14088, n_13447, n_13448);
  and g25535 (n14089, n_12786, n_12784);
  not g25536 (n_13449, n14089);
  and g25537 (n14090, n_12785, n_13449);
  not g25538 (n_13450, n14088);
  and g25539 (n14091, n_13450, n14090);
  not g25540 (n_13451, n14090);
  and g25541 (n14092, n14088, n_13451);
  not g25542 (n_13452, n14091);
  not g25543 (n_13453, n14092);
  and g25544 (n14093, n_13452, n_13453);
  not g25545 (n_13454, n14082);
  not g25546 (n_13455, n14093);
  and g25547 (n14094, n_13454, n_13455);
  not g25554 (n_13456, n14100);
  and g25555 (n14101, n_12826, n_13456);
  and g25556 (n14102, n_12822, n_12823);
  not g25557 (n_13457, n14101);
  not g25558 (n_13458, n14102);
  and g25559 (n14103, n_13457, n_13458);
  not g25560 (n_13459, n14097);
  and g25561 (n14104, n_13459, n14103);
  not g25562 (n_13460, n14094);
  and g25563 (n14105, n_13460, n14104);
  and g25564 (n14106, n_13460, n_13459);
  not g25565 (n_13461, n14103);
  not g25566 (n_13462, n14106);
  and g25567 (n14107, n_13461, n_13462);
  not g25568 (n_13463, n14105);
  not g25569 (n_13464, n14107);
  and g25570 (n14108, n_13463, n_13464);
  not g25571 (n_13465, n14076);
  not g25572 (n_13466, n14108);
  and g25573 (n14109, n_13465, n_13466);
  not g25577 (n_13467, n14109);
  not g25578 (n_13468, n14112);
  and g25579 (n14113, n_13467, n_13468);
  and g25580 (n14114, n_12875, n_12876);
  not g25581 (n_13469, n14114);
  and g25582 (n14115, n_12879, n_13469);
  not g25586 (n_13470, n14115);
  not g25587 (n_13471, n14118);
  and g25588 (n14119, n_13470, n_13471);
  not g25592 (n_13472, n14122);
  and g25593 (n14123, n_12871, n_13472);
  and g25594 (n14124, n_12867, n_12868);
  not g25595 (n_13473, n14123);
  not g25596 (n_13474, n14124);
  and g25597 (n14125, n_13473, n_13474);
  not g25601 (n_13475, n14128);
  and g25602 (n14129, n_12854, n_13475);
  and g25603 (n14130, n_12850, n_12851);
  not g25604 (n_13476, n14129);
  not g25605 (n_13477, n14130);
  and g25606 (n14131, n_13476, n_13477);
  not g25607 (n_13478, n14125);
  and g25608 (n14132, n_13478, n14131);
  not g25609 (n_13479, n14131);
  and g25610 (n14133, n14125, n_13479);
  not g25611 (n_13480, n14132);
  not g25612 (n_13481, n14133);
  and g25613 (n14134, n_13480, n_13481);
  not g25614 (n_13482, n14119);
  not g25615 (n_13483, n14134);
  and g25616 (n14135, n_13482, n_13483);
  not g25620 (n_13484, n14135);
  not g25621 (n_13485, n14138);
  and g25622 (n14139, n_13484, n_13485);
  not g25623 (n_13486, n14113);
  and g25624 (n14140, n_13486, n14139);
  not g25625 (n_13487, n14139);
  and g25626 (n14141, n_13467, n_13487);
  and g25627 (n14142, n_13468, n14141);
  not g25628 (n_13488, n14140);
  not g25629 (n_13489, n14142);
  and g25630 (n14143, n_13488, n_13489);
  not g25631 (n_13490, n14071);
  not g25632 (n_13491, n14143);
  and g25633 (n14144, n_13490, n_13491);
  and g25634 (n14145, n14071, n14143);
  not g25635 (n_13492, n14144);
  not g25636 (n_13493, n14145);
  and g25637 (n14146, n_13492, n_13493);
  not g25638 (n_13494, n14066);
  and g25639 (n14147, n_13494, n14146);
  not g25640 (n_13495, n14146);
  and g25641 (n14148, n14066, n_13495);
  not g25642 (n_13496, n14147);
  not g25643 (n_13497, n14148);
  and g25644 (n14149, n_13496, n_13497);
  not g25645 (n_13498, n13932);
  not g25646 (n_13499, n14149);
  and g25647 (n14150, n_13498, n_13499);
  and g25648 (n14151, n13932, n14149);
  not g25649 (n_13500, n14150);
  not g25650 (n_13501, n14151);
  and g25651 (n14152, n_13500, n_13501);
  and g25652 (n14153, n_13319, n_13320);
  not g25653 (n_13502, n14153);
  and g25654 (n14154, n_13323, n_13502);
  and g25655 (n14155, n13799, n13917);
  not g25656 (n_13503, n14154);
  not g25657 (n_13504, n14155);
  and g25658 (n14156, n_13503, n_13504);
  and g25659 (n14157, n_13311, n_13312);
  not g25660 (n_13505, n14157);
  and g25661 (n14158, n_13315, n_13505);
  and g25662 (n14159, n13857, n13911);
  not g25663 (n_13506, n14158);
  not g25664 (n_13507, n14159);
  and g25665 (n14160, n_13506, n_13507);
  and g25666 (n14161, n_13303, n_13304);
  not g25667 (n_13508, n14161);
  and g25668 (n14162, n_13307, n_13508);
  not g25672 (n_13509, n14162);
  not g25673 (n_13510, n14165);
  and g25674 (n14166, n_13509, n_13510);
  not g25678 (n_13511, n14169);
  and g25679 (n14170, n_13299, n_13511);
  and g25680 (n14171, n_13295, n_13296);
  not g25681 (n_13512, n14170);
  not g25682 (n_13513, n14171);
  and g25683 (n14172, n_13512, n_13513);
  not g25687 (n_13514, n14175);
  and g25688 (n14176, n_13282, n_13514);
  and g25689 (n14177, n_13278, n_13279);
  not g25690 (n_13515, n14176);
  not g25691 (n_13516, n14177);
  and g25692 (n14178, n_13515, n_13516);
  not g25693 (n_13517, n14172);
  and g25694 (n14179, n_13517, n14178);
  not g25695 (n_13518, n14178);
  and g25696 (n14180, n14172, n_13518);
  not g25697 (n_13519, n14179);
  not g25698 (n_13520, n14180);
  and g25699 (n14181, n_13519, n_13520);
  not g25700 (n_13521, n14166);
  not g25701 (n_13522, n14181);
  and g25702 (n14182, n_13521, n_13522);
  not g25706 (n_13523, n14182);
  not g25707 (n_13524, n14185);
  and g25708 (n14186, n_13523, n_13524);
  and g25709 (n14187, n_13258, n_13259);
  not g25710 (n_13525, n14187);
  and g25711 (n14188, n_13262, n_13525);
  not g25715 (n_13526, n14188);
  not g25716 (n_13527, n14191);
  and g25717 (n14192, n_13526, n_13527);
  not g25721 (n_13528, n14195);
  and g25722 (n14196, n_13254, n_13528);
  and g25723 (n14197, n_13250, n_13251);
  not g25724 (n_13529, n14196);
  not g25725 (n_13530, n14197);
  and g25726 (n14198, n_13529, n_13530);
  not g25730 (n_13531, n14201);
  and g25731 (n14202, n_13237, n_13531);
  and g25732 (n14203, n_13233, n_13234);
  not g25733 (n_13532, n14202);
  not g25734 (n_13533, n14203);
  and g25735 (n14204, n_13532, n_13533);
  not g25736 (n_13534, n14198);
  and g25737 (n14205, n_13534, n14204);
  not g25738 (n_13535, n14204);
  and g25739 (n14206, n14198, n_13535);
  not g25740 (n_13536, n14205);
  not g25741 (n_13537, n14206);
  and g25742 (n14207, n_13536, n_13537);
  not g25743 (n_13538, n14192);
  not g25744 (n_13539, n14207);
  and g25745 (n14208, n_13538, n_13539);
  not g25749 (n_13540, n14208);
  not g25750 (n_13541, n14211);
  and g25751 (n14212, n_13540, n_13541);
  not g25752 (n_13542, n14186);
  and g25753 (n14213, n_13542, n14212);
  not g25754 (n_13543, n14212);
  and g25755 (n14214, n14186, n_13543);
  not g25756 (n_13544, n14213);
  not g25757 (n_13545, n14214);
  and g25758 (n14215, n_13544, n_13545);
  not g25759 (n_13546, n14160);
  not g25760 (n_13547, n14215);
  and g25761 (n14216, n_13546, n_13547);
  and g25762 (n14217, n14160, n14215);
  not g25763 (n_13548, n14216);
  not g25764 (n_13549, n14217);
  and g25765 (n14218, n_13548, n_13549);
  and g25766 (n14219, n_13210, n_13211);
  not g25767 (n_13550, n14219);
  and g25768 (n14220, n_13214, n_13550);
  and g25769 (n14221, n13739, n13793);
  not g25770 (n_13551, n14220);
  not g25771 (n_13552, n14221);
  and g25772 (n14222, n_13551, n_13552);
  and g25773 (n14223, n_13202, n_13203);
  not g25774 (n_13553, n14223);
  and g25775 (n14224, n_13206, n_13553);
  not g25779 (n_13554, n14224);
  not g25780 (n_13555, n14227);
  and g25781 (n14228, n_13554, n_13555);
  not g25785 (n_13556, n14231);
  and g25786 (n14232, n_13198, n_13556);
  and g25787 (n14233, n_13194, n_13195);
  not g25788 (n_13557, n14232);
  not g25789 (n_13558, n14233);
  and g25790 (n14234, n_13557, n_13558);
  not g25794 (n_13559, n14237);
  and g25795 (n14238, n_13181, n_13559);
  and g25796 (n14239, n_13177, n_13178);
  not g25797 (n_13560, n14238);
  not g25798 (n_13561, n14239);
  and g25799 (n14240, n_13560, n_13561);
  not g25800 (n_13562, n14234);
  and g25801 (n14241, n_13562, n14240);
  not g25802 (n_13563, n14240);
  and g25803 (n14242, n14234, n_13563);
  not g25804 (n_13564, n14241);
  not g25805 (n_13565, n14242);
  and g25806 (n14243, n_13564, n_13565);
  not g25807 (n_13566, n14228);
  not g25808 (n_13567, n14243);
  and g25809 (n14244, n_13566, n_13567);
  not g25813 (n_13568, n14244);
  not g25814 (n_13569, n14247);
  and g25815 (n14248, n_13568, n_13569);
  and g25816 (n14249, n_13157, n_13158);
  not g25817 (n_13570, n14249);
  and g25818 (n14250, n_13161, n_13570);
  not g25822 (n_13571, n14250);
  not g25823 (n_13572, n14253);
  and g25824 (n14254, n_13571, n_13572);
  not g25828 (n_13573, n14257);
  and g25829 (n14258, n_13153, n_13573);
  and g25830 (n14259, n_13149, n_13150);
  not g25831 (n_13574, n14258);
  not g25832 (n_13575, n14259);
  and g25833 (n14260, n_13574, n_13575);
  not g25837 (n_13576, n14263);
  and g25838 (n14264, n_13136, n_13576);
  and g25839 (n14265, n_13132, n_13133);
  not g25840 (n_13577, n14264);
  not g25841 (n_13578, n14265);
  and g25842 (n14266, n_13577, n_13578);
  not g25843 (n_13579, n14260);
  and g25844 (n14267, n_13579, n14266);
  not g25845 (n_13580, n14266);
  and g25846 (n14268, n14260, n_13580);
  not g25847 (n_13581, n14267);
  not g25848 (n_13582, n14268);
  and g25849 (n14269, n_13581, n_13582);
  not g25850 (n_13583, n14254);
  not g25851 (n_13584, n14269);
  and g25852 (n14270, n_13583, n_13584);
  not g25856 (n_13585, n14270);
  not g25857 (n_13586, n14273);
  and g25858 (n14274, n_13585, n_13586);
  not g25859 (n_13587, n14248);
  and g25860 (n14275, n_13587, n14274);
  not g25861 (n_13588, n14274);
  and g25862 (n14276, n14248, n_13588);
  not g25863 (n_13589, n14275);
  not g25864 (n_13590, n14276);
  and g25865 (n14277, n_13589, n_13590);
  not g25866 (n_13591, n14222);
  not g25867 (n_13592, n14277);
  and g25868 (n14278, n_13591, n_13592);
  and g25869 (n14279, n14222, n14277);
  not g25870 (n_13593, n14278);
  not g25871 (n_13594, n14279);
  and g25872 (n14280, n_13593, n_13594);
  not g25873 (n_13595, n14218);
  and g25874 (n14281, n_13595, n14280);
  not g25875 (n_13596, n14280);
  and g25876 (n14282, n14218, n_13596);
  not g25877 (n_13597, n14281);
  not g25878 (n_13598, n14282);
  and g25879 (n14283, n_13597, n_13598);
  not g25880 (n_13599, n14156);
  not g25881 (n_13600, n14283);
  and g25882 (n14284, n_13599, n_13600);
  and g25883 (n14285, n14156, n14283);
  not g25884 (n_13601, n14284);
  not g25885 (n_13602, n14285);
  and g25886 (n14286, n_13601, n_13602);
  not g25887 (n_13603, n14152);
  not g25888 (n_13604, n14286);
  and g25889 (n14287, n_13603, n_13604);
  not g25890 (n_13605, n13928);
  not g25891 (n_13606, n14287);
  and g25892 (n14288, n_13605, n_13606);
  and g25893 (n14289, n_13500, n14286);
  and g25894 (n14290, n_13501, n14289);
  not g25895 (n_13607, n14288);
  not g25896 (n_13608, n14290);
  and g25897 (n14291, n_13607, n_13608);
  and g25898 (n14292, n_13494, n_13495);
  not g25899 (n_13609, n14292);
  and g25900 (n14293, n_13498, n_13609);
  and g25901 (n14294, n14066, n14146);
  not g25902 (n_13610, n14293);
  not g25903 (n_13611, n14294);
  and g25904 (n14295, n_13610, n_13611);
  and g25905 (n14296, n_13486, n_13487);
  not g25906 (n_13612, n14296);
  and g25907 (n14297, n_13490, n_13612);
  and g25908 (n14298, n_13467, n14139);
  and g25909 (n14299, n_13468, n14298);
  not g25910 (n_13613, n14297);
  not g25911 (n_13614, n14299);
  and g25912 (n14300, n_13613, n_13614);
  not g25916 (n_13615, n14303);
  and g25917 (n14304, n_13482, n_13615);
  and g25918 (n14305, n_13478, n_13479);
  not g25919 (n_13616, n14304);
  not g25920 (n_13617, n14305);
  and g25921 (n14306, n_13616, n_13617);
  and g25922 (n14307, n14103, n_13462);
  not g25923 (n_13618, n14307);
  and g25924 (n14308, n_13465, n_13618);
  and g25925 (n14309, n_13459, n_13461);
  and g25926 (n14310, n_13460, n14309);
  not g25927 (n_13619, n14308);
  not g25928 (n_13620, n14310);
  and g25929 (n14311, n_13619, n_13620);
  not g25933 (n_13621, n14314);
  and g25934 (n14315, n_13454, n_13621);
  and g25935 (n14316, n_13450, n_13451);
  not g25936 (n_13622, n14315);
  not g25937 (n_13623, n14316);
  and g25938 (n14317, n_13622, n_13623);
  not g25939 (n_13624, n14311);
  and g25940 (n14318, n_13624, n14317);
  not g25941 (n_13625, n14317);
  and g25942 (n14319, n_13620, n_13625);
  and g25943 (n14320, n_13619, n14319);
  not g25944 (n_13626, n14318);
  not g25945 (n_13627, n14320);
  and g25946 (n14321, n_13626, n_13627);
  not g25947 (n_13628, n14306);
  not g25948 (n_13629, n14321);
  and g25949 (n14322, n_13628, n_13629);
  and g25950 (n14323, n14306, n_13627);
  and g25951 (n14324, n_13626, n14323);
  not g25952 (n_13630, n14322);
  not g25953 (n_13631, n14324);
  and g25954 (n14325, n_13630, n_13631);
  not g25955 (n_13632, n14300);
  and g25956 (n14326, n_13632, n14325);
  not g25957 (n_13633, n14325);
  and g25958 (n14327, n14300, n_13633);
  not g25959 (n_13634, n14326);
  not g25960 (n_13635, n14327);
  and g25961 (n14328, n_13634, n_13635);
  and g25962 (n14329, n_13429, n_13430);
  not g25963 (n_13636, n14329);
  and g25964 (n14330, n_13433, n_13636);
  and g25965 (n14331, n13998, n14060);
  not g25966 (n_13637, n14330);
  not g25967 (n_13638, n14331);
  and g25968 (n14332, n_13637, n_13638);
  and g25969 (n14333, n_13421, n_13422);
  not g25970 (n_13639, n14333);
  and g25971 (n14334, n_13425, n_13639);
  not g25975 (n_13640, n14334);
  not g25976 (n_13641, n14337);
  and g25977 (n14338, n_13640, n_13641);
  not g25981 (n_13642, n14341);
  and g25982 (n14342, n_13400, n_13642);
  and g25983 (n14343, n_13396, n_13397);
  not g25984 (n_13643, n14342);
  not g25985 (n_13644, n14343);
  and g25986 (n14344, n_13643, n_13644);
  not g25990 (n_13645, n14347);
  and g25991 (n14348, n_13417, n_13645);
  and g25992 (n14349, n_13413, n_13414);
  not g25993 (n_13646, n14348);
  not g25994 (n_13647, n14349);
  and g25995 (n14350, n_13646, n_13647);
  not g25996 (n_13648, n14344);
  and g25997 (n14351, n_13648, n14350);
  not g25998 (n_13649, n14350);
  and g25999 (n14352, n14344, n_13649);
  not g26000 (n_13650, n14351);
  not g26001 (n_13651, n14352);
  and g26002 (n14353, n_13650, n_13651);
  not g26003 (n_13652, n14338);
  not g26004 (n_13653, n14353);
  and g26005 (n14354, n_13652, n_13653);
  not g26009 (n_13654, n14354);
  not g26010 (n_13655, n14357);
  and g26011 (n14358, n_13654, n_13655);
  and g26012 (n14359, n_13376, n_13377);
  not g26013 (n_13656, n14359);
  and g26014 (n14360, n_13380, n_13656);
  not g26018 (n_13657, n14360);
  not g26019 (n_13658, n14363);
  and g26020 (n14364, n_13657, n_13658);
  not g26024 (n_13659, n14367);
  and g26025 (n14368, n_13355, n_13659);
  and g26026 (n14369, n_13351, n_13352);
  not g26027 (n_13660, n14368);
  not g26028 (n_13661, n14369);
  and g26029 (n14370, n_13660, n_13661);
  not g26033 (n_13662, n14373);
  and g26034 (n14374, n_13372, n_13662);
  and g26035 (n14375, n_13368, n_13369);
  not g26036 (n_13663, n14374);
  not g26037 (n_13664, n14375);
  and g26038 (n14376, n_13663, n_13664);
  not g26039 (n_13665, n14370);
  and g26040 (n14377, n_13665, n14376);
  not g26041 (n_13666, n14376);
  and g26042 (n14378, n14370, n_13666);
  not g26043 (n_13667, n14377);
  not g26044 (n_13668, n14378);
  and g26045 (n14379, n_13667, n_13668);
  not g26046 (n_13669, n14364);
  not g26047 (n_13670, n14379);
  and g26048 (n14380, n_13669, n_13670);
  not g26052 (n_13671, n14380);
  not g26053 (n_13672, n14383);
  and g26054 (n14384, n_13671, n_13672);
  not g26055 (n_13673, n14358);
  and g26056 (n14385, n_13673, n14384);
  not g26057 (n_13674, n14384);
  and g26058 (n14386, n14358, n_13674);
  not g26059 (n_13675, n14385);
  not g26060 (n_13676, n14386);
  and g26061 (n14387, n_13675, n_13676);
  not g26062 (n_13677, n14332);
  not g26063 (n_13678, n14387);
  and g26064 (n14388, n_13677, n_13678);
  and g26065 (n14389, n14332, n14387);
  not g26066 (n_13679, n14388);
  not g26067 (n_13680, n14389);
  and g26068 (n14390, n_13679, n_13680);
  not g26069 (n_13681, n14328);
  and g26070 (n14391, n_13681, n14390);
  not g26071 (n_13682, n14390);
  and g26072 (n14392, n14328, n_13682);
  not g26073 (n_13683, n14391);
  not g26074 (n_13684, n14392);
  and g26075 (n14393, n_13683, n_13684);
  not g26076 (n_13685, n14295);
  not g26077 (n_13686, n14393);
  and g26078 (n14394, n_13685, n_13686);
  and g26079 (n14395, n14295, n14393);
  not g26080 (n_13687, n14394);
  not g26081 (n_13688, n14395);
  and g26082 (n14396, n_13687, n_13688);
  and g26083 (n14397, n_13595, n_13596);
  not g26084 (n_13689, n14397);
  and g26085 (n14398, n_13599, n_13689);
  and g26086 (n14399, n14218, n14280);
  not g26087 (n_13690, n14398);
  not g26088 (n_13691, n14399);
  and g26089 (n14400, n_13690, n_13691);
  and g26090 (n14401, n_13587, n_13588);
  not g26091 (n_13692, n14401);
  and g26092 (n14402, n_13591, n_13692);
  not g26096 (n_13693, n14402);
  not g26097 (n_13694, n14405);
  and g26098 (n14406, n_13693, n_13694);
  not g26102 (n_13695, n14409);
  and g26103 (n14410, n_13566, n_13695);
  and g26104 (n14411, n_13562, n_13563);
  not g26105 (n_13696, n14410);
  not g26106 (n_13697, n14411);
  and g26107 (n14412, n_13696, n_13697);
  not g26111 (n_13698, n14415);
  and g26112 (n14416, n_13583, n_13698);
  and g26113 (n14417, n_13579, n_13580);
  not g26114 (n_13699, n14416);
  not g26115 (n_13700, n14417);
  and g26116 (n14418, n_13699, n_13700);
  not g26117 (n_13701, n14412);
  and g26118 (n14419, n_13701, n14418);
  not g26119 (n_13702, n14418);
  and g26120 (n14420, n14412, n_13702);
  not g26121 (n_13703, n14419);
  not g26122 (n_13704, n14420);
  and g26123 (n14421, n_13703, n_13704);
  not g26124 (n_13705, n14406);
  not g26125 (n_13706, n14421);
  and g26126 (n14422, n_13705, n_13706);
  not g26130 (n_13707, n14422);
  not g26131 (n_13708, n14425);
  and g26132 (n14426, n_13707, n_13708);
  and g26133 (n14427, n_13542, n_13543);
  not g26134 (n_13709, n14427);
  and g26135 (n14428, n_13546, n_13709);
  not g26139 (n_13710, n14428);
  not g26140 (n_13711, n14431);
  and g26141 (n14432, n_13710, n_13711);
  not g26145 (n_13712, n14435);
  and g26146 (n14436, n_13521, n_13712);
  and g26147 (n14437, n_13517, n_13518);
  not g26148 (n_13713, n14436);
  not g26149 (n_13714, n14437);
  and g26150 (n14438, n_13713, n_13714);
  not g26154 (n_13715, n14441);
  and g26155 (n14442, n_13538, n_13715);
  and g26156 (n14443, n_13534, n_13535);
  not g26157 (n_13716, n14442);
  not g26158 (n_13717, n14443);
  and g26159 (n14444, n_13716, n_13717);
  not g26160 (n_13718, n14438);
  and g26161 (n14445, n_13718, n14444);
  not g26162 (n_13719, n14444);
  and g26163 (n14446, n14438, n_13719);
  not g26164 (n_13720, n14445);
  not g26165 (n_13721, n14446);
  and g26166 (n14447, n_13720, n_13721);
  not g26167 (n_13722, n14432);
  not g26168 (n_13723, n14447);
  and g26169 (n14448, n_13722, n_13723);
  not g26173 (n_13724, n14448);
  not g26174 (n_13725, n14451);
  and g26175 (n14452, n_13724, n_13725);
  not g26176 (n_13726, n14426);
  and g26177 (n14453, n_13726, n14452);
  not g26178 (n_13727, n14452);
  and g26179 (n14454, n14426, n_13727);
  not g26180 (n_13728, n14453);
  not g26181 (n_13729, n14454);
  and g26182 (n14455, n_13728, n_13729);
  not g26183 (n_13730, n14400);
  not g26184 (n_13731, n14455);
  and g26185 (n14456, n_13730, n_13731);
  and g26186 (n14457, n14400, n14455);
  not g26187 (n_13732, n14456);
  not g26188 (n_13733, n14457);
  and g26189 (n14458, n_13732, n_13733);
  not g26190 (n_13734, n14396);
  not g26191 (n_13735, n14458);
  and g26192 (n14459, n_13734, n_13735);
  not g26193 (n_13736, n14291);
  not g26194 (n_13737, n14459);
  and g26195 (n14460, n_13736, n_13737);
  and g26196 (n14461, n_13687, n14458);
  and g26197 (n14462, n_13688, n14461);
  not g26198 (n_13738, n14460);
  not g26199 (n_13739, n14462);
  and g26200 (n14463, n_13738, n_13739);
  and g26201 (n14464, n_13681, n_13682);
  not g26202 (n_13740, n14464);
  and g26203 (n14465, n_13685, n_13740);
  and g26204 (n14466, n14328, n14390);
  not g26205 (n_13741, n14465);
  not g26206 (n_13742, n14466);
  and g26207 (n14467, n_13741, n_13742);
  and g26208 (n14468, n_13632, n_13631);
  not g26209 (n_13743, n14468);
  and g26210 (n14469, n_13630, n_13743);
  and g26211 (n14470, n_13624, n_13625);
  not g26212 (n_13744, n14469);
  and g26213 (n14471, n_13744, n14470);
  not g26214 (n_13745, n14470);
  and g26215 (n14472, n_13630, n_13745);
  and g26216 (n14473, n_13743, n14472);
  not g26217 (n_13746, n14471);
  not g26218 (n_13747, n14473);
  and g26219 (n14474, n_13746, n_13747);
  and g26220 (n14475, n_13673, n_13674);
  not g26221 (n_13748, n14475);
  and g26222 (n14476, n_13677, n_13748);
  not g26226 (n_13749, n14476);
  not g26227 (n_13750, n14479);
  and g26228 (n14480, n_13749, n_13750);
  not g26232 (n_13751, n14483);
  and g26233 (n14484, n_13669, n_13751);
  and g26234 (n14485, n_13665, n_13666);
  not g26235 (n_13752, n14484);
  not g26236 (n_13753, n14485);
  and g26237 (n14486, n_13752, n_13753);
  not g26241 (n_13754, n14489);
  and g26242 (n14490, n_13652, n_13754);
  and g26243 (n14491, n_13648, n_13649);
  not g26244 (n_13755, n14490);
  not g26245 (n_13756, n14491);
  and g26246 (n14492, n_13755, n_13756);
  not g26247 (n_13757, n14486);
  and g26248 (n14493, n_13757, n14492);
  not g26249 (n_13758, n14492);
  and g26250 (n14494, n14486, n_13758);
  not g26251 (n_13759, n14493);
  not g26252 (n_13760, n14494);
  and g26253 (n14495, n_13759, n_13760);
  not g26254 (n_13761, n14480);
  not g26255 (n_13762, n14495);
  and g26256 (n14496, n_13761, n_13762);
  not g26260 (n_13763, n14496);
  not g26261 (n_13764, n14499);
  and g26262 (n14500, n_13763, n_13764);
  not g26263 (n_13765, n14474);
  not g26264 (n_13766, n14500);
  and g26265 (n14501, n_13765, n_13766);
  not g26269 (n_13767, n14501);
  not g26270 (n_13768, n14504);
  and g26271 (n14505, n_13767, n_13768);
  not g26272 (n_13769, n14467);
  and g26273 (n14506, n_13769, n14505);
  not g26274 (n_13770, n14505);
  and g26275 (n14507, n14467, n_13770);
  not g26276 (n_13771, n14506);
  not g26277 (n_13772, n14507);
  and g26278 (n14508, n_13771, n_13772);
  and g26279 (n14509, n_13726, n_13727);
  not g26280 (n_13773, n14509);
  and g26281 (n14510, n_13730, n_13773);
  not g26285 (n_13774, n14510);
  not g26286 (n_13775, n14513);
  and g26287 (n14514, n_13774, n_13775);
  not g26291 (n_13776, n14517);
  and g26292 (n14518, n_13722, n_13776);
  and g26293 (n14519, n_13718, n_13719);
  not g26294 (n_13777, n14518);
  not g26295 (n_13778, n14519);
  and g26296 (n14520, n_13777, n_13778);
  not g26300 (n_13779, n14523);
  and g26301 (n14524, n_13705, n_13779);
  and g26302 (n14525, n_13701, n_13702);
  not g26303 (n_13780, n14524);
  not g26304 (n_13781, n14525);
  and g26305 (n14526, n_13780, n_13781);
  not g26306 (n_13782, n14520);
  and g26307 (n14527, n_13782, n14526);
  not g26308 (n_13783, n14526);
  and g26309 (n14528, n14520, n_13783);
  not g26310 (n_13784, n14527);
  not g26311 (n_13785, n14528);
  and g26312 (n14529, n_13784, n_13785);
  not g26313 (n_13786, n14514);
  not g26314 (n_13787, n14529);
  and g26315 (n14530, n_13786, n_13787);
  not g26319 (n_13788, n14530);
  not g26320 (n_13789, n14533);
  and g26321 (n14534, n_13788, n_13789);
  not g26322 (n_13790, n14508);
  not g26323 (n_13791, n14534);
  and g26324 (n14535, n_13790, n_13791);
  not g26325 (n_13792, n14463);
  not g26326 (n_13793, n14535);
  and g26327 (n14536, n_13792, n_13793);
  and g26328 (n14537, n_13771, n14534);
  and g26329 (n14538, n_13772, n14537);
  not g26330 (n_13794, n14536);
  not g26331 (n_13795, n14538);
  and g26332 (n14539, n_13794, n_13795);
  and g26333 (n14540, n_13769, n_13767);
  not g26334 (n_13796, n14540);
  and g26335 (n14541, n_13768, n_13796);
  not g26339 (n_13797, n14544);
  and g26340 (n14545, n_13761, n_13797);
  and g26341 (n14546, n_13757, n_13758);
  not g26342 (n_13798, n14546);
  and g26343 (n14547, n_13746, n_13798);
  not g26344 (n_13799, n14545);
  and g26345 (n14548, n_13799, n14547);
  and g26346 (n14549, n_13799, n_13798);
  not g26347 (n_13800, n14549);
  and g26348 (n14550, n14471, n_13800);
  not g26349 (n_13801, n14548);
  not g26350 (n_13802, n14550);
  and g26351 (n14551, n_13801, n_13802);
  not g26352 (n_13803, n14541);
  and g26353 (n14552, n_13803, n14551);
  not g26354 (n_13804, n14551);
  and g26355 (n14553, n_13768, n_13804);
  and g26356 (n14554, n_13796, n14553);
  not g26357 (n_13805, n14552);
  not g26358 (n_13806, n14554);
  and g26359 (n14555, n_13805, n_13806);
  not g26363 (n_13807, n14558);
  and g26364 (n14559, n_13786, n_13807);
  and g26365 (n14560, n_13782, n_13783);
  not g26366 (n_13808, n14559);
  not g26367 (n_13809, n14560);
  and g26368 (n14561, n_13808, n_13809);
  not g26369 (n_13810, n14555);
  and g26370 (n14562, n_13810, n14561);
  not g26371 (n_13811, n14539);
  not g26372 (n_13812, n14562);
  and g26373 (n14563, n_13811, n_13812);
  not g26374 (n_13813, n14561);
  and g26375 (n14564, n_13806, n_13813);
  and g26376 (n14565, n_13805, n14564);
  not g26377 (n_13814, n14563);
  not g26378 (n_13815, n14565);
  and g26379 (n14566, n_13814, n_13815);
  and g26380 (n14567, n_13803, n_13801);
  not g26381 (n_13816, n14567);
  and g26382 (n14568, n_13802, n_13816);
  not g26383 (n_13817, n14566);
  and g26384 (n14569, n_13817, n14568);
  not g26385 (n_13818, n14568);
  and g26386 (n14570, n_13815, n_13818);
  and g26387 (n14571, n_13814, n14570);
  not g26388 (n_13819, n14569);
  not g26389 (n_13820, n14571);
  and g26390 (n14572, n_13819, n_13820);
  and g26391 (n14573, n_13810, n_13813);
  and g26392 (n14574, n_13806, n14561);
  and g26393 (n14575, n_13805, n14574);
  not g26394 (n_13821, n14575);
  not g26397 (n_13822, n14573);
  and g26399 (n14579, n_13822, n_13821);
  not g26400 (n_13823, n14579);
  and g26401 (n14580, n_13811, n_13823);
  and g26402 (n14581, n_13790, n14534);
  and g26403 (n14582, n_13771, n_13791);
  and g26404 (n14583, n_13772, n14582);
  not g26405 (n_13824, n14581);
  not g26406 (n_13825, n14583);
  and g26407 (n14584, n_13824, n_13825);
  and g26408 (n14585, n14463, n14584);
  not g26409 (n_13826, n14584);
  and g26410 (n14586, n_13792, n_13826);
  and g26411 (n14587, n_13687, n_13735);
  and g26412 (n14588, n_13688, n14587);
  and g26413 (n14589, n_13734, n14458);
  not g26414 (n_13827, n14588);
  not g26415 (n_13828, n14589);
  and g26416 (n14590, n_13827, n_13828);
  and g26417 (n14591, n14291, n14590);
  not g26418 (n_13829, n14590);
  and g26419 (n14592, n_13736, n_13829);
  and g26420 (n14593, n_13603, n14286);
  and g26421 (n14594, n_13500, n_13604);
  and g26422 (n14595, n_13501, n14594);
  not g26423 (n_13830, n14593);
  not g26424 (n_13831, n14595);
  and g26425 (n14596, n_13830, n_13831);
  and g26426 (n14597, n13928, n14596);
  not g26427 (n_13832, n14596);
  and g26428 (n14598, n_13605, n_13832);
  and g26429 (n14599, n_13112, n_13328);
  and g26430 (n14600, n_13113, n14599);
  and g26431 (n14601, n_13327, n13923);
  not g26432 (n_13833, n14600);
  not g26433 (n_13834, n14601);
  and g26434 (n14602, n_13833, n_13834);
  and g26435 (n14603, n13275, n14602);
  not g26436 (n_13835, n14602);
  and g26437 (n14604, n_13329, n_13835);
  and g26438 (n14605, n_12761, n13270);
  and g26439 (n14606, n_12322, n_12762);
  and g26440 (n14607, n_12323, n14606);
  not g26441 (n_13836, n14605);
  not g26442 (n_13837, n14607);
  and g26443 (n14608, n_13836, n_13837);
  and g26444 (n14609, n11871, n14608);
  not g26445 (n_13838, n14608);
  and g26446 (n14610, n_12763, n_13838);
  and g26447 (n14611, n_10978, n_11612);
  and g26448 (n14612, n_10979, n14611);
  and g26449 (n14613, n_11611, n11866);
  not g26450 (n_13839, n14612);
  not g26451 (n_13840, n14613);
  and g26452 (n14614, n_13839, n_13840);
  not g26453 (n_13841, n14614);
  and g26454 (n14615, n_11613, n_13841);
  and g26455 (n14616, n_9951, n_9949);
  and g26456 (n14617, n_9950, n14616);
  and g26457 (n14618, n10032, n_9952);
  not g26458 (n_13842, n14617);
  not g26459 (n_13843, n14618);
  and g26460 (n14619, n_13842, n_13843);
  not g26461 (n_13845, n14619);
  and g26462 (n14620, \A[1000] , n_13845);
  not g26463 (n_13846, n14615);
  and g26465 (n14622, n10047, n14614);
  and g26466 (n14623, n10036, n_9957);
  and g26467 (n14624, n_9958, n14623);
  and g26468 (n14625, n_9956, n_9961);
  not g26469 (n_13847, n14624);
  not g26470 (n_13848, n14625);
  and g26471 (n14626, n_13847, n_13848);
  not g26472 (n_13849, n14626);
  and g26473 (n14627, n4472, n_13849);
  and g26474 (n14628, n_9960, n_9963);
  not g26475 (n_13850, n14628);
  and g26476 (n14629, n_9959, n_13850);
  not g26477 (n_13851, n14627);
  not g26478 (n_13852, n14629);
  and g26479 (n14630, n_13851, n_13852);
  not g26480 (n_13853, n14622);
  not g26481 (n_13854, n14630);
  not g26484 (n_13855, n14610);
  and g26485 (n14633, n_13855, n14632);
  not g26486 (n_13856, n14609);
  and g26487 (n14634, n_13856, n14633);
  not g26488 (n_13857, n14604);
  and g26489 (n14635, n_13857, n14634);
  not g26490 (n_13858, n14603);
  and g26491 (n14636, n_13858, n14635);
  not g26492 (n_13859, n14598);
  and g26493 (n14637, n_13859, n14636);
  not g26494 (n_13860, n14597);
  and g26495 (n14638, n_13860, n14637);
  not g26496 (n_13861, n14592);
  and g26497 (n14639, n_13861, n14638);
  not g26498 (n_13862, n14591);
  and g26499 (n14640, n_13862, n14639);
  not g26500 (n_13863, n14586);
  and g26501 (n14641, n_13863, n14640);
  not g26502 (n_13864, n14585);
  and g26503 (n14642, n_13864, n14641);
  not g26504 (n_13865, n14580);
  and g26505 (n14643, n_13865, n14642);
  not g26506 (n_13866, n14578);
  and g26507 (n14644, n_13866, n14643);
  and g26508 (n14645, n14572, n14644);
  not g26509 (n_13867, n14572);
  not g26510 (n_13868, n14644);
  and g26511 (n14646, n_13867, n_13868);
  not g26512 (n_13869, n14645);
  not g26513 (n_13870, n14646);
  and g26514 (n14647, n_13869, n_13870);
  and g26515 (n14648, n_13866, n_13865);
  not g26516 (n_13871, n14642);
  not g26517 (n_13872, n14648);
  and g26518 (n14649, n_13871, n_13872);
  and g26519 (n14650, n_13864, n_13863);
  not g26520 (n_13873, n14640);
  not g26521 (n_13874, n14650);
  and g26522 (n14651, n_13873, n_13874);
  and g26523 (n14652, n_13862, n_13861);
  not g26524 (n_13875, n14638);
  not g26525 (n_13876, n14652);
  and g26526 (n14653, n_13875, n_13876);
  and g26527 (n14654, n_13856, n_13855);
  not g26528 (n_13877, n14632);
  not g26529 (n_13878, n14654);
  and g26530 (n14655, n_13877, n_13878);
  and g26531 (n14656, n_13846, n_13853);
  and g26532 (n14657, n14620, n_13854);
  not g26533 (n_13879, n14656);
  not g26534 (n_13880, n14657);
  and g26535 (n14658, n_13879, n_13880);
  not g26536 (n_13881, n14658);
  and g26537 (n14659, n_13877, n_13881);
  and g26538 (n14660, n14620, n_13851);
  and g26539 (n14661, n_13852, n14660);
  not g26540 (n_13882, n14620);
  and g26541 (n14662, n_13882, n_13854);
  not g26542 (n_13883, n14661);
  not g26543 (n_13884, n14662);
  and g26544 (n14663, n_13883, n_13884);
  not g26545 (n_13885, n14659);
  and g26546 (n14664, n_13885, n14663);
  not g26547 (n_13886, n14634);
  not g26548 (n_13887, n14664);
  and g26549 (n14665, n_13886, n_13887);
  not g26550 (n_13888, n14655);
  and g26551 (n14666, n_13888, n14665);
  and g26552 (n14667, n_13858, n_13857);
  not g26553 (n_13889, n14667);
  and g26554 (n14668, n_13886, n_13889);
  not g26555 (n_13890, n14636);
  not g26556 (n_13891, n14668);
  and g26557 (n14669, n_13890, n_13891);
  not g26558 (n_13892, n14666);
  not g26559 (n_13893, n14669);
  and g26560 (n14670, n_13892, n_13893);
  and g26561 (n14671, n_13860, n_13859);
  not g26562 (n_13894, n14671);
  and g26563 (n14672, n_13890, n_13894);
  not g26564 (n_13895, n14672);
  and g26565 (n14673, n_13875, n_13895);
  not g26566 (n_13896, n14670);
  and g26567 (n14674, n_13896, n14673);
  and g26568 (n14675, n_13873, n14674);
  not g26569 (n_13897, n14653);
  and g26570 (n14676, n_13897, n14675);
  and g26571 (n14677, n_13871, n14676);
  not g26572 (n_13898, n14651);
  and g26573 (n14678, n_13898, n14677);
  and g26574 (n14679, n_13868, n14678);
  not g26575 (n_13899, n14649);
  and g26576 (n14680, n_13899, n14679);
  not g26577 (n_13900, n14647);
  and g26578 (n14681, n_13900, n14680);
  and g26579 (n14682, n_13867, n14644);
  and g26580 (n14683, n_13817, n_13818);
  not g26581 (n_13901, n14682);
  and g26582 (n14684, n_13901, n14683);
  not g26583 (n_13902, n14683);
  and g26584 (n14685, n14644, n_13902);
  and g26585 (n14686, n_13867, n14685);
  not g26592 (n_13903, n14686);
  not g26595 (n_13905, n14684);
  not g26597 (n_13906, n14681);
  and g26599 (n14696, n_13871, n_13898);
  and g26600 (n14697, n_13886, n_13888);
  not g26601 (n_13907, n14697);
  and g26602 (n14698, n14664, n_13907);
  not g26603 (n_13908, n14698);
  and g26604 (n14699, n_13892, n_13908);
  not g26605 (n_13909, n14663);
  and g26606 (n14700, n14659, n_13909);
  and g26607 (n14701, \A[1000] , n_13842);
  and g26608 (n14702, n_13843, n14701);
  not g26609 (n_13910, \A[1000] );
  and g26610 (n14703, n_13910, n_13845);
  not g26611 (n_13911, n14702);
  not g26612 (n_13912, n14703);
  and g26613 (n14704, n_13911, n_13912);
  and g26614 (n14705, n_13887, n14704);
  not g26615 (n_13913, n14700);
  and g26616 (n14706, n_13913, n14705);
  not g26617 (n_13914, n14706);
  and g26618 (n14707, n14659, n_13914);
  and g26619 (n14708, n_13887, n_13913);
  not g26620 (n_13915, n14704);
  not g26621 (n_13916, n14708);
  and g26622 (n14709, n_13915, n_13916);
  not g26623 (n_13917, n14707);
  not g26624 (n_13918, n14709);
  and g26625 (n14710, n_13917, n_13918);
  not g26626 (n_13919, n14699);
  and g26627 (n14711, n_13919, n14710);
  not g26628 (n_13920, n14711);
  and g26629 (n14712, n14697, n_13920);
  not g26630 (n_13921, n14710);
  and g26631 (n14713, n14699, n_13921);
  not g26632 (n_13922, n14712);
  not g26633 (n_13923, n14713);
  and g26634 (n14714, n_13922, n_13923);
  not g26635 (n_13924, n14714);
  and g26636 (n14715, n_13892, n_13924);
  and g26637 (n14716, n_13890, n14666);
  and g26638 (n14717, n_13891, n14716);
  not g26639 (n_13925, n14673);
  and g26640 (n14718, n14670, n_13925);
  not g26641 (n_13926, n14674);
  not g26642 (n_13927, n14718);
  and g26643 (n14719, n_13926, n_13927);
  not g26644 (n_13928, n14717);
  not g26645 (n_13929, n14719);
  and g26646 (n14720, n_13928, n_13929);
  not g26647 (n_13930, n14715);
  and g26648 (n14721, n_13930, n14720);
  not g26649 (n_13931, n14721);
  and g26650 (n14722, n14673, n_13931);
  and g26651 (n14723, n_13930, n_13928);
  not g26652 (n_13932, n14723);
  and g26653 (n14724, n14719, n_13932);
  not g26654 (n_13933, n14722);
  not g26655 (n_13934, n14724);
  and g26656 (n14725, n_13933, n_13934);
  not g26657 (n_13935, n14725);
  and g26658 (n14726, n14674, n_13935);
  and g26659 (n14727, n_13873, n_13897);
  and g26660 (n14728, n_13926, n14727);
  not g26661 (n_13936, n14676);
  not g26662 (n_13937, n14696);
  and g26663 (n14729, n_13936, n_13937);
  not g26664 (n_13938, n14678);
  not g26665 (n_13939, n14729);
  and g26666 (n14730, n_13938, n_13939);
  not g26667 (n_13940, n14728);
  not g26668 (n_13941, n14730);
  and g26669 (n14731, n_13940, n_13941);
  not g26670 (n_13942, n14726);
  and g26671 (n14732, n_13942, n14731);
  not g26672 (n_13943, n14732);
  and g26673 (n14733, n14696, n_13943);
  and g26674 (n14734, n_13942, n_13940);
  not g26675 (n_13944, n14734);
  and g26676 (n14735, n14730, n_13944);
  not g26677 (n_13945, n14733);
  not g26678 (n_13946, n14735);
  and g26679 (n14736, n_13945, n_13946);
  not g26680 (n_13947, n14680);
  and g26681 (n14737, n14678, n_13947);
  not g26682 (n_13948, n14736);
  and g26683 (n14738, n_13948, n14737);
  and g26684 (n14739, n14680, n_13945);
  and g26685 (n14740, n_13946, n14739);
  and g26686 (n14741, n_13868, n_13899);
  not g26687 (n_13949, n14740);
  and g26688 (n14742, n_13949, n14741);
  not g26689 (n_13950, n14738);
  not g26690 (n_13951, n14742);
  and g26691 (n14743, n_13950, n_13951);
  and g26692 (n14744, n14680, n_13906);
  not g26693 (n_13952, n14743);
  and g26694 (n14745, n_13952, n14744);
  and g26695 (n14746, n14681, n_13950);
  and g26696 (n14747, n_13951, n14746);
  not g26697 (n_13953, n14747);
  and g26698 (n14748, n_13900, n_13953);
  not g26699 (n_13954, n14748);
  and g26700 (n14749, n_13906, n_13954);
  not g26701 (n_13955, n14745);
  and g26702 (n14750, n_13955, n14749);
  and g26706 (n14754, n_13905, n_13903);
  and g26707 (n14755, n_13906, n14754);
  not g26708 (n_13956, n14755);
  and g26709 (n14756, n14692, n_13956);
  not g26710 (n_13957, n14695);
  not g26711 (n_13958, n14756);
  and g26712 (n14757, n_13957, n_13958);
  not g26713 (n_13959, n14753);
  not g26714 (n_13960, n14757);
  and g26715 (n14758, n_13959, n_13960);
  not g26716 (n_13961, n14750);
  and g26717 (n14759, n_13961, n14758);
  or g26718 (maj, n_13957, n14759);
  and g26719 (n14695, n_13963, n_13906, n_13905, n_13903);
  not g26720 (n_13963, n14692);
  and g26721 (n14753, n_13900, n_13905, n14680, n_13903);
  and g26722 (n_13964, n_13867, n_13817);
  and g26724 (n_13966, n14650, n_13818);
  and g26725 (n14692, n14640, n_13964, n14648, n_13966);
  and g26726 (n14578, n_13822, n_13794, n_13795, n_13821);
  and g26727 (n14632, n_13846, n14620, n_13853, n_13854);
  and g26728 (n14533, n_13774, n_13785, n_13775, n_13784);
  and g26729 (n14558, n_13777, n_13780, n_13778, n_13781);
  and g26730 (n14504, n_13763, n_13746, n_13747, n_13764);
  and g26731 (n14513, n_13707, n_13724, n_13708, n_13725);
  and g26732 (n14544, n_13752, n_13755, n_13753, n_13756);
  and g26733 (n14499, n_13749, n_13760, n_13750, n_13759);
  and g26734 (n14425, n_13693, n_13704, n_13694, n_13703);
  and g26735 (n14451, n_13710, n_13721, n_13711, n_13720);
  and g26736 (n14517, n_13713, n_13716, n_13714, n_13717);
  and g26737 (n14523, n_13696, n_13699, n_13697, n_13700);
  and g26738 (n14314, n_13447, n_13449, n_12785, n_13448);
  and g26739 (n14303, n_13473, n_13476, n_13474, n_13477);
  and g26740 (n14479, n_13654, n_13671, n_13655, n_13672);
  and g26741 (n14483, n_13660, n_13663, n_13661, n_13664);
  and g26742 (n14489, n_13643, n_13646, n_13644, n_13647);
  and g26743 (n14405, n_13568, n_13585, n_13569, n_13586);
  and g26744 (n14431, n_13523, n_13540, n_13524, n_13541);
  and g26745 (n14097, n_13444, n_13453, n_13445, n_13452);
  and g26746 (n14435, n_13512, n_13515, n_13513, n_13516);
  and g26747 (n14441, n_13529, n_13532, n_13530, n_13533);
  and g26748 (n14409, n_13557, n_13560, n_13558, n_13561);
  and g26749 (n14415, n_13574, n_13577, n_13575, n_13578);
  and g26750 (n14112, n_13464, n_13441, n_13442, n_13463);
  and g26751 (n14138, n_13470, n_13481, n_13471, n_13480);
  and g26752 (n14081, n_12788, n_12805, n_12789, n_12806);
  and g26753 (n14085, n_12794, n_12797, n_12795, n_12798);
  and g26754 (n14357, n_13640, n_13651, n_13641, n_13650);
  and g26755 (n14383, n_13657, n_13668, n_13658, n_13667);
  and g26756 (n14247, n_13554, n_13565, n_13555, n_13564);
  and g26757 (n14273, n_13571, n_13582, n_13572, n_13581);
  and g26758 (n14185, n_13509, n_13520, n_13510, n_13519);
  and g26759 (n14211, n_13526, n_13537, n_13527, n_13536);
  and g26760 (n14118, n_12856, n_12873, n_12857, n_12874);
  and g26761 (n14122, n_12862, n_12865, n_12863, n_12866);
  and g26762 (n14128, n_12845, n_12848, n_12846, n_12849);
  and g26763 (n14100, n_12817, n_12820, n_12818, n_12821);
  and g26764 (n14363, n_13357, n_13374, n_13358, n_13375);
  and g26765 (n14367, n_13346, n_13349, n_13347, n_13350);
  and g26766 (n14373, n_13363, n_13366, n_13364, n_13367);
  and g26767 (n14337, n_13402, n_13419, n_13403, n_13420);
  and g26768 (n14341, n_13391, n_13394, n_13392, n_13395);
  and g26769 (n14347, n_13408, n_13411, n_13409, n_13412);
  and g26770 (n13328, n_12791, n_12802, n_12792, n_12801);
  and g26771 (n14227, n_13183, n_13200, n_13184, n_13201);
  and g26772 (n14253, n_13138, n_13155, n_13139, n_13156);
  and g26773 (n14165, n_13284, n_13301, n_13285, n_13302);
  and g26774 (n14191, n_13239, n_13256, n_13240, n_13257);
  and g26775 (n14169, n_13290, n_13293, n_13291, n_13294);
  and g26776 (n14175, n_13273, n_13276, n_13274, n_13277);
  and g26777 (n14195, n_13245, n_13248, n_13246, n_13249);
  and g26778 (n14201, n_13228, n_13231, n_13229, n_13232);
  and g26779 (n14231, n_13189, n_13192, n_13190, n_13193);
  and g26780 (n14237, n_13172, n_13175, n_13173, n_13176);
  and g26781 (n14257, n_13144, n_13147, n_13145, n_13148);
  and g26782 (n14263, n_13127, n_13130, n_13128, n_13131);
  and g26783 (n13388, n_12842, n_12853, n_12843, n_12852);
  and g26784 (n13410, n_12859, n_12870, n_12860, n_12869);
  and g26785 (n13355, n_12814, n_12825, n_12815, n_12824);
  and g26786 (n13312, n_12084, n_12101, n_12085, n_12102);
  and g26787 (n13965, n_13343, n_13354, n_13344, n_13353);
  and g26788 (n13991, n_13360, n_13371, n_13361, n_13370);
  and g26789 (n14027, n_13388, n_13399, n_13389, n_13398);
  and g26790 (n14053, n_13405, n_13416, n_13406, n_13415);
  and g26791 (n13394, n_12228, n_12245, n_12229, n_12246);
  and g26792 (n13372, n_12273, n_12290, n_12274, n_12291);
  and g26793 (n13339, n_12172, n_12189, n_12173, n_12190);
  and g26794 (n13945, n_13063, n_13080, n_13064, n_13081);
  and g26795 (n13949, n_13069, n_13072, n_13070, n_13073);
  and g26796 (n13955, n_13052, n_13055, n_13053, n_13056);
  and g26797 (n13971, n_13018, n_13035, n_13019, n_13036);
  and g26798 (n13975, n_13024, n_13027, n_13025, n_13028);
  and g26799 (n13981, n_13007, n_13010, n_13008, n_13011);
  and g26800 (n14007, n_12962, n_12979, n_12963, n_12980);
  and g26801 (n14011, n_12968, n_12971, n_12969, n_12972);
  and g26802 (n14017, n_12951, n_12954, n_12952, n_12955);
  and g26803 (n14033, n_12917, n_12934, n_12918, n_12935);
  and g26804 (n14037, n_12923, n_12926, n_12924, n_12927);
  and g26805 (n14043, n_12906, n_12909, n_12907, n_12910);
  and g26806 (n13764, n_13169, n_13180, n_13170, n_13179);
  and g26807 (n13786, n_13186, n_13197, n_13187, n_13196);
  and g26808 (n13710, n_13124, n_13135, n_13125, n_13134);
  and g26809 (n13732, n_13141, n_13152, n_13142, n_13151);
  and g26810 (n13882, n_13270, n_13281, n_13271, n_13280);
  and g26811 (n13904, n_13287, n_13298, n_13288, n_13297);
  and g26812 (n13828, n_13225, n_13236, n_13226, n_13235);
  and g26813 (n13850, n_13242, n_13253, n_13243, n_13252);
  and g26814 (n12450, n_12070, n_12081, n_12071, n_12080);
  and g26815 (n12474, n_12087, n_12098, n_12088, n_12097);
  and g26816 (n12519, n_12122, n_12133, n_12123, n_12132);
  and g26817 (n13888, n_12351, n_12368, n_12352, n_12369);
  and g26818 (n13866, n_12396, n_12413, n_12397, n_12414);
  and g26819 (n13834, n_12452, n_12469, n_12453, n_12470);
  and g26820 (n13812, n_12497, n_12514, n_12498, n_12515);
  and g26821 (n13770, n_12564, n_12581, n_12565, n_12582);
  and g26822 (n13748, n_12609, n_12626, n_12610, n_12627);
  and g26823 (n13716, n_12665, n_12682, n_12666, n_12683);
  and g26824 (n13694, n_12710, n_12727, n_12711, n_12728);
  and g26825 (n12628, n_12214, n_12225, n_12215, n_12224);
  and g26826 (n12652, n_12231, n_12242, n_12232, n_12241);
  and g26827 (n12686, n_12259, n_12270, n_12260, n_12269);
  and g26828 (n12710, n_12276, n_12287, n_12277, n_12286);
  and g26829 (n12559, n_12158, n_12169, n_12159, n_12168);
  and g26830 (n12583, n_12175, n_12186, n_12176, n_12185);
  and g26831 (n12432, n_10066, n_10077, n_10067, n_10078);
  and g26832 (n12456, n_10035, n_10046, n_10036, n_10047);
  and g26833 (n12501, n_9995, n_10006, n_9996, n_10007);
  and g26834 (n13630, n_13049, n_13060, n_13050, n_13059);
  and g26835 (n13652, n_13066, n_13077, n_13067, n_13076);
  and g26836 (n13576, n_13004, n_13015, n_13005, n_13014);
  and g26837 (n13598, n_13021, n_13032, n_13022, n_13031);
  and g26838 (n13512, n_12948, n_12959, n_12949, n_12958);
  and g26839 (n13534, n_12965, n_12976, n_12966, n_12975);
  and g26840 (n13458, n_12903, n_12914, n_12904, n_12913);
  and g26841 (n13480, n_12920, n_12931, n_12921, n_12930);
  and g26842 (n12610, n_10294, n_10305, n_10295, n_10306);
  and g26843 (n12634, n_10263, n_10274, n_10264, n_10275);
  and g26844 (n12668, n_10223, n_10234, n_10224, n_10235);
  and g26845 (n12692, n_10192, n_10203, n_10193, n_10204);
  and g26846 (n12541, n_10143, n_10154, n_10144, n_10155);
  and g26847 (n12565, n_10112, n_10123, n_10113, n_10124);
  and g26848 (n13636, n_11647, n_11664, n_11648, n_11665);
  and g26849 (n13614, n_11692, n_11709, n_11693, n_11710);
  and g26850 (n13582, n_11748, n_11765, n_11749, n_11766);
  and g26851 (n13560, n_11793, n_11810, n_11794, n_11811);
  and g26852 (n13518, n_11860, n_11877, n_11861, n_11878);
  and g26853 (n13496, n_11905, n_11922, n_11906, n_11923);
  and g26854 (n13464, n_11961, n_11978, n_11962, n_11979);
  and g26855 (n13442, n_12006, n_12023, n_12007, n_12024);
  and g26856 (n12775, n_12337, n_12348, n_12338, n_12347);
  and g26857 (n12799, n_12354, n_12365, n_12355, n_12364);
  and g26858 (n12833, n_12382, n_12393, n_12383, n_12392);
  and g26859 (n12857, n_12399, n_12410, n_12400, n_12409);
  and g26860 (n12901, n_12438, n_12449, n_12439, n_12448);
  and g26861 (n12925, n_12455, n_12466, n_12456, n_12465);
  and g26862 (n12959, n_12483, n_12494, n_12484, n_12493);
  and g26863 (n12983, n_12500, n_12511, n_12501, n_12510);
  and g26864 (n13037, n_12550, n_12561, n_12551, n_12560);
  and g26865 (n13061, n_12567, n_12578, n_12568, n_12577);
  and g26866 (n13095, n_12595, n_12606, n_12596, n_12605);
  and g26867 (n13119, n_12612, n_12623, n_12613, n_12622);
  and g26868 (n13163, n_12651, n_12662, n_12652, n_12661);
  and g26869 (n13187, n_12668, n_12679, n_12669, n_12678);
  and g26870 (n13221, n_12696, n_12707, n_12697, n_12706);
  and g26871 (n13245, n_12713, n_12724, n_12714, n_12723);
  and g26872 (n10173, n_10057, n_10063, n_4975, n_10062);
  and g26873 (n10187, n_10068, n_10074, n_5072, n_10073);
  and g26874 (n_13967, n_5066, n_5062);
  and g26875 (n5589, n5580, n_5067, n_5068, n_13967);
  and g26876 (n_13968, n_4965, n_4961);
  and g26877 (n5504, n5491, n_4966, n_4967, n_13968);
  and g26878 (n10137, n_10026, n_10032, n_4867, n_10031);
  and g26879 (n10151, n_10037, n_10043, n_4748, n_10042);
  and g26880 (n_13969, n_4742, n_4738);
  and g26881 (n5300, n5291, n_4743, n_4744, n_13969);
  and g26882 (n_13970, n_4801, n_4799);
  and g26883 (n5408, n5395, n_4845, n_4859, n_13970);
  and g26884 (n10077, n_9980, n_9969, n_4644, n_9979);
  and g26885 (n10093, n_9986, n_9992, n_4384, n_9991);
  and g26886 (n10107, n_9997, n_10003, n_4481, n_10002);
  and g26887 (n_13971, n_4475, n_4471);
  and g26888 (n5061, n5052, n_4476, n_4477, n_13971);
  and g26889 (n_13972, n_4374, n_4370);
  and g26890 (n4976, n4963, n_4375, n_4376, n_13972);
  and g26891 (n12757, n_11558, n_11569, n_11559, n_11570);
  and g26892 (n12781, n_11527, n_11538, n_11528, n_11539);
  and g26893 (n12815, n_11487, n_11498, n_11488, n_11499);
  and g26894 (n12839, n_11456, n_11467, n_11457, n_11468);
  and g26895 (n12883, n_11407, n_11418, n_11408, n_11419);
  and g26896 (n12907, n_11376, n_11387, n_11377, n_11388);
  and g26897 (n12941, n_11336, n_11347, n_11337, n_11348);
  and g26898 (n12965, n_11305, n_11316, n_11306, n_11317);
  and g26899 (n13019, n_11247, n_11258, n_11248, n_11259);
  and g26900 (n13043, n_11216, n_11227, n_11217, n_11228);
  and g26901 (n13077, n_11176, n_11187, n_11177, n_11188);
  and g26902 (n13101, n_11145, n_11156, n_11146, n_11157);
  and g26903 (n13145, n_11096, n_11107, n_11097, n_11108);
  and g26904 (n13169, n_11065, n_11076, n_11066, n_11077);
  and g26905 (n13203, n_11025, n_11036, n_11026, n_11037);
  and g26906 (n13227, n_10994, n_11005, n_10995, n_11006);
  and g26907 (n10427, n_10285, n_10291, n_5970, n_10290);
  and g26908 (n10441, n_10296, n_10302, n_5979, n_10301);
  and g26909 (n_13973, n_5195, n_5193);
  and g26910 (n6384, n6375, n_5239, n_5975, n_13973);
  and g26911 (n_13974, n_5287, n_5285);
  and g26912 (n6369, n6356, n_5331, n_5962, n_13974);
  and g26913 (n10391, n_10254, n_10260, n_5950, n_10259);
  and g26914 (n10405, n_10265, n_10271, n_5929, n_10270);
  and g26915 (n_13975, n_5383, n_5381);
  and g26916 (n6315, n6306, n_5427, n_5925, n_13975);
  and g26917 (n_13976, n_5475, n_5473);
  and g26918 (n6343, n6330, n_5519, n_5942, n_13976);
  and g26919 (n10347, n_10214, n_10220, n_6022, n_10219);
  and g26920 (n10361, n_10225, n_10231, n_6031, n_10230);
  and g26921 (n_13977, n_5575, n_5573);
  and g26922 (n6451, n6442, n_5619, n_6027, n_13977);
  and g26923 (n_13978, n_5667, n_5665);
  and g26924 (n6436, n6423, n_5711, n_6014, n_13978);
  and g26925 (n10311, n_10183, n_10189, n_6080, n_10188);
  and g26926 (n10325, n_10194, n_10200, n_6059, n_10199);
  and g26927 (n_13979, n_5763, n_5761);
  and g26928 (n6487, n6478, n_5807, n_6055, n_13979);
  and g26929 (n_13980, n_5855, n_5853);
  and g26930 (n6515, n6502, n_5899, n_6072, n_13980);
  and g26931 (n10258, n_10134, n_10140, n_3921, n_10139);
  and g26932 (n10272, n_10145, n_10151, n_4018, n_10150);
  and g26933 (n_13981, n_4012, n_4008);
  and g26934 (n4643, n4634, n_4013, n_4014, n_13981);
  and g26935 (n_13982, n_3911, n_3907);
  and g26936 (n4558, n4545, n_3912, n_3913, n_13982);
  and g26937 (n10222, n_10103, n_10109, n_4269, n_10108);
  and g26938 (n10236, n_10114, n_10120, n_4248, n_10119);
  and g26939 (n_13983, n_4090, n_4088);
  and g26940 (n4845, n4836, n_4134, n_4244, n_13983);
  and g26941 (n_13984, n_4182, n_4180);
  and g26942 (n4873, n4860, n_4226, n_4261, n_13984);
  and g26943 (n11914, n_11633, n_11644, n_11634, n_11643);
  and g26944 (n11938, n_11650, n_11661, n_11651, n_11660);
  and g26945 (n11972, n_11678, n_11689, n_11679, n_11688);
  and g26946 (n11996, n_11695, n_11706, n_11696, n_11705);
  and g26947 (n12040, n_11734, n_11745, n_11735, n_11744);
  and g26948 (n12064, n_11751, n_11762, n_11752, n_11761);
  and g26949 (n12098, n_11779, n_11790, n_11780, n_11789);
  and g26950 (n12122, n_11796, n_11807, n_11797, n_11806);
  and g26951 (n12176, n_11846, n_11857, n_11847, n_11856);
  and g26952 (n12200, n_11863, n_11874, n_11864, n_11873);
  and g26953 (n12234, n_11891, n_11902, n_11892, n_11901);
  and g26954 (n12258, n_11908, n_11919, n_11909, n_11918);
  and g26955 (n12302, n_11947, n_11958, n_11948, n_11957);
  and g26956 (n12326, n_11964, n_11975, n_11965, n_11974);
  and g26957 (n12360, n_11992, n_12003, n_11993, n_12002);
  and g26958 (n12384, n_12009, n_12020, n_12010, n_12019);
  and g26959 (n11896, n_10919, n_10930, n_10920, n_10931);
  and g26960 (n11920, n_10888, n_10899, n_10889, n_10900);
  and g26961 (n11954, n_10848, n_10859, n_10849, n_10860);
  and g26962 (n11978, n_10817, n_10828, n_10818, n_10829);
  and g26963 (n12022, n_10768, n_10779, n_10769, n_10780);
  and g26964 (n12046, n_10737, n_10748, n_10738, n_10749);
  and g26965 (n12080, n_10697, n_10708, n_10698, n_10709);
  and g26966 (n12104, n_10666, n_10677, n_10667, n_10678);
  and g26967 (n12158, n_10608, n_10619, n_10609, n_10620);
  and g26968 (n12182, n_10577, n_10588, n_10578, n_10589);
  and g26969 (n12216, n_10537, n_10548, n_10538, n_10549);
  and g26970 (n12240, n_10506, n_10517, n_10507, n_10518);
  and g26971 (n12284, n_10457, n_10468, n_10458, n_10469);
  and g26972 (n12308, n_10426, n_10437, n_10427, n_10438);
  and g26973 (n12342, n_10386, n_10397, n_10387, n_10398);
  and g26974 (n12366, n_10355, n_10366, n_10356, n_10367);
  and g26975 (n11821, n_11549, n_11555, n_1727, n_11554);
  and g26976 (n11835, n_11560, n_11566, n_1824, n_11565);
  and g26977 (n_13985, n_1818, n_1814);
  and g26978 (n2645, n2636, n_1819, n_1820, n_13985);
  and g26979 (n_13986, n_1717, n_1713);
  and g26980 (n2560, n2547, n_1718, n_1719, n_13986);
  and g26981 (n11785, n_11518, n_11524, n_1619, n_11523);
  and g26982 (n11799, n_11529, n_11535, n_1500, n_11534);
  and g26983 (n_13987, n_1494, n_1490);
  and g26984 (n2356, n2347, n_1495, n_1496, n_13987);
  and g26985 (n_13988, n_1553, n_1551);
  and g26986 (n2464, n2451, n_1597, n_1611, n_13988);
  and g26987 (n11741, n_11478, n_11484, n_1041, n_11483);
  and g26988 (n11755, n_11489, n_11495, n_1138, n_11494);
  and g26989 (n_13989, n_1132, n_1128);
  and g26990 (n2027, n2018, n_1133, n_1134, n_13989);
  and g26991 (n_13990, n_1031, n_1027);
  and g26992 (n1942, n1929, n_1032, n_1033, n_13990);
  and g26993 (n11705, n_11447, n_11453, n_1389, n_11452);
  and g26994 (n11719, n_11458, n_11464, n_1368, n_11463);
  and g26995 (n_13991, n_1210, n_1208);
  and g26996 (n2229, n2220, n_1254, n_1364, n_13991);
  and g26997 (n_13992, n_1302, n_1300);
  and g26998 (n2257, n2244, n_1346, n_1381, n_13992);
  and g26999 (n11653, n_11398, n_11404, n_321, n_11403);
  and g27000 (n11667, n_11409, n_11415, n_418, n_11414);
  and g27001 (n_13993, n_412, n_408);
  and g27002 (n1373, n1364, n_413, n_414, n_13993);
  and g27003 (n_13994, n_311, n_307);
  and g27004 (n1288, n1275, n_312, n_313, n_13994);
  and g27005 (n11617, n_11367, n_11373, n_213, n_11372);
  and g27006 (n11631, n_11378, n_11384, n_94, n_11383);
  and g27007 (n_13995, n_88, n_84);
  and g27008 (n1084, n1075, n_89, n_90, n_13995);
  and g27009 (n_13996, n_147, n_145);
  and g27010 (n1192, n1179, n_191, n_205, n_13996);
  and g27011 (n11573, n_11327, n_11333, n_861, n_11332);
  and g27012 (n11587, n_11338, n_11344, n_870, n_11343);
  and g27013 (n_13997, n_507, n_505);
  and g27014 (n1768, n1759, n_551, n_866, n_13997);
  and g27015 (n_13998, n_599, n_597);
  and g27016 (n1753, n1740, n_643, n_853, n_13998);
  and g27017 (n11537, n_11296, n_11302, n_919, n_11301);
  and g27018 (n11551, n_11307, n_11313, n_898, n_11312);
  and g27019 (n_13999, n_695, n_693);
  and g27020 (n1804, n1795, n_739, n_894, n_13999);
  and g27021 (n_14000, n_787, n_785);
  and g27022 (n1832, n1819, n_831, n_911, n_14000);
  and g27023 (n11477, n_11238, n_11244, n_3575, n_11243);
  and g27024 (n11491, n_11249, n_11255, n_3584, n_11254);
  and g27025 (n_14001, n_2709, n_2707);
  and g27026 (n4174, n4165, n_2753, n_3580, n_14001);
  and g27027 (n_14002, n_2801, n_2799);
  and g27028 (n4159, n4146, n_2845, n_3567, n_14002);
  and g27029 (n11441, n_11207, n_11213, n_3555, n_11212);
  and g27030 (n11455, n_11218, n_11224, n_3534, n_11223);
  and g27031 (n_14003, n_2897, n_2895);
  and g27032 (n4105, n4096, n_2941, n_3530, n_14003);
  and g27033 (n_14004, n_2989, n_2987);
  and g27034 (n4133, n4120, n_3033, n_3547, n_14004);
  and g27035 (n11397, n_11167, n_11173, n_3453, n_11172);
  and g27036 (n11411, n_11178, n_11184, n_3462, n_11183);
  and g27037 (n_14005, n_3089, n_3087);
  and g27038 (n4012, n4003, n_3133, n_3458, n_14005);
  and g27039 (n_14006, n_3181, n_3179);
  and g27040 (n3997, n3984, n_3225, n_3445, n_14006);
  and g27041 (n11361, n_11136, n_11142, n_3511, n_11141);
  and g27042 (n11375, n_11147, n_11153, n_3490, n_11152);
  and g27043 (n_14007, n_3277, n_3275);
  and g27044 (n4048, n4039, n_3321, n_3486, n_14007);
  and g27045 (n_14008, n_3369, n_3367);
  and g27046 (n4076, n4063, n_3413, n_3503, n_14008);
  and g27047 (n11309, n_11087, n_11093, n_3675, n_11092);
  and g27048 (n11323, n_11098, n_11104, n_3684, n_11103);
  and g27049 (n_14009, n_2325, n_2323);
  and g27050 (n4303, n4294, n_2369, n_3680, n_14009);
  and g27051 (n_14010, n_2417, n_2415);
  and g27052 (n4288, n4275, n_2461, n_3667, n_14010);
  and g27053 (n11273, n_11056, n_11062, n_3655, n_11061);
  and g27054 (n11287, n_11067, n_11073, n_3634, n_11072);
  and g27055 (n_14011, n_2513, n_2511);
  and g27056 (n4234, n4225, n_2557, n_3630, n_14011);
  and g27057 (n_14012, n_2605, n_2603);
  and g27058 (n4262, n4249, n_2649, n_3647, n_14012);
  and g27059 (n11229, n_11016, n_11022, n_3727, n_11021);
  and g27060 (n11243, n_11027, n_11033, n_3736, n_11032);
  and g27061 (n_14013, n_2133, n_2131);
  and g27062 (n4370, n4361, n_2177, n_3732, n_14013);
  and g27063 (n_14014, n_2225, n_2223);
  and g27064 (n4355, n4342, n_2269, n_3719, n_14014);
  and g27065 (n11193, n_10985, n_10991, n_3785, n_10990);
  and g27066 (n11207, n_10996, n_11002, n_3764, n_11001);
  and g27067 (n_14015, n_2037, n_2035);
  and g27068 (n4406, n4397, n_2081, n_3760, n_14015);
  and g27069 (n_14016, n_1945, n_1943);
  and g27070 (n4434, n4421, n_1989, n_3777, n_14016);
  and g27071 (n11119, n_10910, n_10916, n_9741, n_10915);
  and g27072 (n11133, n_10921, n_10927, n_9838, n_10926);
  and g27073 (n_14017, n_9832, n_9828);
  and g27074 (n9915, n9906, n_9833, n_9834, n_14017);
  and g27075 (n_14018, n_9731, n_9727);
  and g27076 (n9830, n9817, n_9732, n_9733, n_14018);
  and g27077 (n11083, n_10879, n_10885, n_9633, n_10884);
  and g27078 (n11097, n_10890, n_10896, n_9514, n_10895);
  and g27079 (n_14019, n_9508, n_9504);
  and g27080 (n9626, n9617, n_9509, n_9510, n_14019);
  and g27081 (n_14020, n_9567, n_9565);
  and g27082 (n9734, n9721, n_9611, n_9625, n_14020);
  and g27083 (n11039, n_10839, n_10845, n_9055, n_10844);
  and g27084 (n11053, n_10850, n_10856, n_9152, n_10855);
  and g27085 (n_14021, n_9146, n_9142);
  and g27086 (n9297, n9288, n_9147, n_9148, n_14021);
  and g27087 (n_14022, n_9045, n_9041);
  and g27088 (n9212, n9199, n_9046, n_9047, n_14022);
  and g27089 (n11003, n_10808, n_10814, n_9403, n_10813);
  and g27090 (n11017, n_10819, n_10825, n_9382, n_10824);
  and g27091 (n_14023, n_9224, n_9222);
  and g27092 (n9499, n9490, n_9268, n_9378, n_14023);
  and g27093 (n_14024, n_9316, n_9314);
  and g27094 (n9527, n9514, n_9360, n_9395, n_14024);
  and g27095 (n10951, n_10759, n_10765, n_8335, n_10764);
  and g27096 (n10965, n_10770, n_10776, n_8432, n_10775);
  and g27097 (n_14025, n_8426, n_8422);
  and g27098 (n8643, n8634, n_8427, n_8428, n_14025);
  and g27099 (n_14026, n_8325, n_8321);
  and g27100 (n8558, n8545, n_8326, n_8327, n_14026);
  and g27101 (n10915, n_10728, n_10734, n_8227, n_10733);
  and g27102 (n10929, n_10739, n_10745, n_8108, n_10744);
  and g27103 (n_14027, n_8102, n_8098);
  and g27104 (n8354, n8345, n_8103, n_8104, n_14027);
  and g27105 (n_14028, n_8161, n_8159);
  and g27106 (n8462, n8449, n_8205, n_8219, n_14028);
  and g27107 (n10871, n_10688, n_10694, n_8875, n_10693);
  and g27108 (n10885, n_10699, n_10705, n_8884, n_10704);
  and g27109 (n_14029, n_8521, n_8519);
  and g27110 (n9038, n9029, n_8565, n_8880, n_14029);
  and g27111 (n_14030, n_8613, n_8611);
  and g27112 (n9023, n9010, n_8657, n_8867, n_14030);
  and g27113 (n10835, n_10657, n_10663, n_8933, n_10662);
  and g27114 (n10849, n_10668, n_10674, n_8912, n_10673);
  and g27115 (n_14031, n_8709, n_8707);
  and g27116 (n9074, n9065, n_8753, n_8908, n_14031);
  and g27117 (n_14032, n_8801, n_8799);
  and g27118 (n9102, n9089, n_8845, n_8925, n_14032);
  and g27119 (n10775, n_10599, n_10605, n_6895, n_10604);
  and g27120 (n10789, n_10610, n_10616, n_6992, n_10615);
  and g27121 (n_14033, n_6986, n_6982);
  and g27122 (n7335, n7326, n_6987, n_6988, n_14033);
  and g27123 (n_14034, n_6885, n_6881);
  and g27124 (n7250, n7237, n_6886, n_6887, n_14034);
  and g27125 (n10739, n_10568, n_10574, n_6787, n_10573);
  and g27126 (n10753, n_10579, n_10585, n_6668, n_10584);
  and g27127 (n_14035, n_6662, n_6658);
  and g27128 (n7046, n7037, n_6663, n_6664, n_14035);
  and g27129 (n_14036, n_6721, n_6719);
  and g27130 (n7154, n7141, n_6765, n_6779, n_14036);
  and g27131 (n10695, n_10528, n_10534, n_6209, n_10533);
  and g27132 (n10709, n_10539, n_10545, n_6306, n_10544);
  and g27133 (n_14037, n_6300, n_6296);
  and g27134 (n6717, n6708, n_6301, n_6302, n_14037);
  and g27135 (n_14038, n_6199, n_6195);
  and g27136 (n6632, n6619, n_6200, n_6201, n_14038);
  and g27137 (n10659, n_10497, n_10503, n_6557, n_10502);
  and g27138 (n10673, n_10508, n_10514, n_6536, n_10513);
  and g27139 (n_14039, n_6378, n_6376);
  and g27140 (n6919, n6910, n_6422, n_6532, n_14039);
  and g27141 (n_14040, n_6470, n_6468);
  and g27142 (n6947, n6934, n_6514, n_6549, n_14040);
  and g27143 (n10607, n_10448, n_10454, n_7873, n_10453);
  and g27144 (n10621, n_10459, n_10465, n_7882, n_10464);
  and g27145 (n_14041, n_7098, n_7096);
  and g27146 (n8110, n8101, n_7142, n_7878, n_14041);
  and g27147 (n_14042, n_7190, n_7188);
  and g27148 (n8095, n8082, n_7234, n_7865, n_14042);
  and g27149 (n10571, n_10417, n_10423, n_7853, n_10422);
  and g27150 (n10585, n_10428, n_10434, n_7832, n_10433);
  and g27151 (n_14043, n_7286, n_7284);
  and g27152 (n8041, n8032, n_7330, n_7828, n_14043);
  and g27153 (n_14044, n_7378, n_7376);
  and g27154 (n8069, n8056, n_7422, n_7845, n_14044);
  and g27155 (n10527, n_10377, n_10383, n_7925, n_10382);
  and g27156 (n10541, n_10388, n_10394, n_7934, n_10393);
  and g27157 (n_14045, n_7478, n_7476);
  and g27158 (n8177, n8168, n_7522, n_7930, n_14045);
  and g27159 (n_14046, n_7570, n_7568);
  and g27160 (n8162, n8149, n_7614, n_7917, n_14046);
  and g27161 (n10491, n_10346, n_10352, n_7983, n_10351);
  and g27162 (n10505, n_10357, n_10363, n_7962, n_10362);
  and g27163 (n_14047, n_7666, n_7664);
  and g27164 (n8213, n8204, n_7710, n_7958, n_14047);
  and g27165 (n_14048, n_7758, n_7756);
  and g27166 (n8241, n8228, n_7802, n_7975, n_14048);
endmodule
