//# 62 inputs
//# 152 outputs
//# 638 D-type flipflops
//# 5378 inverters
//# 2573 gates (1114 ANDs + 849 NANDs + 512 ORs + 98 NORs)



module s13207 (clock, g43, g49, g633, g634, g635, g645, g647,
     g648, g690, g694, g698, g702, g722, g723, g751, g752, g753, g754,
     g755, g756, g757, g781, g941, g962, g1000, g1008, g1016, g1080,
     g1234, g1554, g206, g291, g372, g453, g534, g594, g785, g1006,
     g1015, g1017, g1246, g1724, g1783, g1798, g1804, g1810, g1817,
     g1824, g1829, g1870, g1871, g1894, g1911, g1944, g2662, g2844,
     g2888, g3077, g3096, g3130, g3159, g3191, g3829, g3859, g3860,
     g4267, g4316, g4370, g4371, g4372, g4373, g4655, g4657, g4660,
     g4661, g4663, g4664, g5143, g5164, g5571, g5669, g5678, g5682,
     g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269, g6425,
     g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063,
     g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290,
     g7291, g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425,
     g7474, g7504, g7505, g7506, g7507, g7508, g7514, g7729, g7730,
     g7731, g7732, g8216, g8217, g8218, g8219, g8234, g8661, g8663,
     g8872, g8958, g9128, g9132, g9204, g9280, g9297, g9299, g9305,
     g9308, g9310, g9312, g9314, g9378);
  input clock, g43, g49, g633, g634, g635, g645, g647, g648, g690,
       g694, g698, g702, g722, g723, g751, g752, g753, g754, g755,
       g756, g757, g781, g941, g962, g1000, g1008, g1016, g1080, g1234,
       g1554;
  output g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017,
       g1246, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829,
       g1870, g1871, g1894, g1911, g1944, g2662, g2844, g2888, g3077,
       g3096, g3130, g3159, g3191, g3829, g3859, g3860, g4267, g4316,
       g4370, g4371, g4372, g4373, g4655, g4657, g4660, g4661, g4663,
       g4664, g5143, g5164, g5571, g5669, g5678, g5682, g5684, g5687,
       g5729, g6207, g6212, g6223, g6236, g6269, g6425, g6648, g6653,
       g6675, g6849, g6850, g6895, g6909, g7048, g7063, g7103, g7283,
       g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291, g7292,
       g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504,
       g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732,
       g8216, g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958,
       g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310,
       g9312, g9314, g9378;
  wire clock, g43, g49, g633, g634, g635, g645, g647, g648, g690, g694,
       g698, g702, g722, g723, g751, g752, g753, g754, g755, g756,
       g757, g781, g941, g962, g1000, g1008, g1016, g1080, g1234, g1554;
  wire g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017,
       g1246, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829,
       g1870, g1871, g1894, g1911, g1944, g2662, g2844, g2888, g3077,
       g3096, g3130, g3159, g3191, g3829, g3859, g3860, g4267, g4316,
       g4370, g4371, g4372, g4373, g4655, g4657, g4660, g4661, g4663,
       g4664, g5143, g5164, g5571, g5669, g5678, g5682, g5684, g5687,
       g5729, g6207, g6212, g6223, g6236, g6269, g6425, g6648, g6653,
       g6675, g6849, g6850, g6895, g6909, g7048, g7063, g7103, g7283,
       g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291, g7292,
       g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504,
       g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732,
       g8216, g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958,
       g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310,
       g9312, g9314, g9378;
  wire g652, g866, g871, g929, g933, g936, g940, g942;
  wire g944, g969, g971, g972, g973, g979, g984, g985;
  wire g990, g995, g998, g999, g1033, g1037, g1041, g1045;
  wire g1049, g1053, g1057, g1061, g1065, g1069, g1077, g1087;
  wire g1092, g1097, g1098, g1102, g1106, g1110, g1114, g1118;
  wire g1122, g1126, g1130, g1134, g1138, g1142, g1149, g1166;
  wire g1176, g1179, g1189, g1253, g1257, g1263, g1266, g1267;
  wire g1268, g1269, g1304, g1313, g1354, g1360, g1363, g1364;
  wire g1365, g1366, g1367, g1368, g1369, g1370, g1371, g1372;
  wire g1373, g1374, g1375, g1408, g1415, g1416, g1421, g1428;
  wire g1430, g1435, g1439, g1444, g1450, g1454, g1462, g1467;
  wire g1472, g1481, g1489, g1494, g1499, g1504, g1509, g1514;
  wire g1519, g_1796, g_1800, g_1801, g_1820, g_1821, g_1822, g_1823;
  wire g_1824, g_1827, g_1828, g_1829, g_1830, g_1831, g_1832, g_1833;
  wire g_1834, g_1835, g_1844, n_0, n_1, n_2, n_3, n_4;
  wire n_5, n_6, n_7, n_8, n_9, n_12, n_15, n_17;
  wire n_19, n_22, n_24, n_25, n_26, n_27, n_28, n_29;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45;
  wire n_46, n_47, n_48, n_49, n_50, n_52, n_53, n_55;
  wire n_56, n_57, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_100, n_101, n_103, n_104, n_105, n_106, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_115, n_116, n_117;
  wire n_118, n_119, n_120, n_121, n_122, n_124, n_125, n_126;
  wire n_127, n_128, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_165, n_166, n_167, n_168, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_219, n_221, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_253;
  wire n_254, n_255, n_256, n_257, n_258, n_260, n_261, n_262;
  wire n_263, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_276, n_277, n_278, n_280, n_281;
  wire n_282, n_283, n_285, n_286, n_287, n_288, n_290, n_291;
  wire n_292, n_293, n_295, n_296, n_297, n_298, n_299, n_300;
  wire n_301, n_302, n_304, n_305, n_306, n_307, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_326, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395;
  wire n_396, n_397, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444;
  wire n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476;
  wire n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484;
  wire n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492;
  wire n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500;
  wire n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508;
  wire n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516;
  wire n_517, n_519, n_520, n_521, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533;
  wire n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541;
  wire n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581;
  wire n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589;
  wire n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597;
  wire n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605;
  wire n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613;
  wire n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621;
  wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
  wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669;
  wire n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677;
  wire n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_706;
  wire n_708, n_709, n_710, n_712, n_713, n_714, n_715, n_716;
  wire n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724;
  wire n_725, n_726, n_727, n_728, n_729, n_730, n_731, new_I6791_;
  wire new_I6864_, new_I8094_, new_I8446_, new_I11008_, new_g1616_,
       new_g2216_, new_g2298_, new_g2407_;
  wire new_g2562_, new_g2573_, new_g2584_, new_g2605_, new_g2665_,
       new_g2668_, new_g2712_, new_g2727_;
  wire new_g2728_, new_g2734_, new_g2746_, new_g2752_, new_g2770_,
       new_g2784_, new_g2959_, new_g3019_;
  wire new_g3029_, new_g3038_, new_g3052_, new_g3062_, new_g3124_,
       new_g3533_, new_g3549_, new_g3568_;
  wire new_g3583_, new_g3605_, new_g3617_, new_g3635_, new_g3644_,
       new_g3666_, new_g3684_, new_g3694_;
  wire new_g3700_, new_g3707_, new_g3712_, new_g3716_, new_g3728_,
       new_g3732_, new_g3735_, new_g3750_;
  wire new_g3753_, new_g3754_, new_g3757_, new_g3768_, new_g3769_,
       new_g3778_, new_g3779_;
  assign g9378 = 1'b1;
  assign g9314 = 1'b1;
  assign g9312 = 1'b1;
  assign g9310 = 1'b1;
  assign g9308 = 1'b1;
  assign g9305 = 1'b1;
  assign g9299 = 1'b1;
  assign g9297 = 1'b1;
  assign g9280 = 1'b1;
  assign g9204 = 1'b0;
  assign g9132 = g8234;
  assign g9128 = 1'b0;
  assign g8958 = 1'b1;
  assign g8872 = 1'b1;
  assign g8663 = g7063;
  assign g8661 = 1'b0;
  assign g8219 = g6675;
  assign g8218 = g6425;
  assign g8217 = g6653;
  assign g8216 = g6648;
  assign g7732 = g6223;
  assign g7731 = g6236;
  assign g7730 = g6212;
  assign g7729 = 1'b0;
  assign g7508 = g5687;
  assign g7507 = g5684;
  assign g7506 = g5682;
  assign g7505 = g5678;
  assign g7504 = g5669;
  assign g7474 = 1'b1;
  assign g7298 = 1'b0;
  assign g7295 = 1'b1;
  assign g7294 = 1'b1;
  assign g7293 = 1'b1;
  assign g7292 = 1'b1;
  assign g7291 = 1'b1;
  assign g7290 = 1'b1;
  assign g7289 = 1'b1;
  assign g7288 = 1'b1;
  assign g7287 = 1'b1;
  assign g7286 = 1'b1;
  assign g7285 = 1'b1;
  assign g7284 = 1'b1;
  assign g7283 = 1'b1;
  assign g6909 = g1008;
  assign g6895 = 1'b1;
  assign g6849 = 1'b0;
  assign g6269 = g1000;
  assign g6207 = 1'b0;
  assign g5729 = g49;
  assign g5164 = 1'b0;
  assign g5143 = g1554;
  assign g4664 = 1'b0;
  assign g4663 = 1'b0;
  assign g4661 = 1'b0;
  assign g4660 = 1'b0;
  assign g4316 = 1'b0;
  assign g3860 = g3829;
  assign g3859 = g3829;
  assign g3191 = 1'b0;
  assign g3159 = 1'b0;
  assign g3130 = 1'b0;
  assign g3096 = 1'b0;
  assign g3077 = 1'b0;
  assign g2844 = 1'b0;
  assign g1911 = 1'b0;
  assign g1870 = 1'b0;
  assign g1829 = 1'b0;
  assign g1824 = 1'b0;
  assign g1817 = 1'b0;
  assign g1810 = 1'b0;
  assign g1804 = 1'b0;
  assign g1798 = 1'b0;
  assign g1783 = 1'b0;
  assign g1017 = 1'b0;
  assign g1015 = 1'b0;
  assign g1006 = 1'b0;
  assign g594 = g206;
  assign g534 = g206;
  assign g453 = g206;
  assign g372 = g206;
  assign g291 = g206;
  fflopd g1102_reg(.CK (clock), .D (n_684), .Q (g1102));
  fflopd g1087_reg(.CK (clock), .D (n_683), .Q (g1087));
  fflopd g1110_reg(.CK (clock), .D (n_674), .Q (g1110));
  fflopd g1126_reg(.CK (clock), .D (n_679), .Q (g1126));
  fflopd g1118_reg(.CK (clock), .D (n_677), .Q (g1118));
  fflopd g1106_reg(.CK (clock), .D (n_681), .Q (g1106));
  fflopd g1122_reg(.CK (clock), .D (n_676), .Q (g1122));
  fflopd g1114_reg(.CK (clock), .D (n_675), .Q (g1114));
  not g24689 (n_684, n_682);
  not g24690 (n_683, n_678);
  fflopd g1142_reg(.CK (clock), .D (n_672), .Q (g1142));
  fflopd g1098_reg(.CK (clock), .D (n_673), .Q (g1098));
  nand g24692__2398 (n_682, n_680, n_307);
  nand g24691__5107 (n_681, n_680, n_263);
  nand g24699__6260 (n_679, n_680, n_363);
  nand g24693__4319 (n_678, n_680, n_225);
  nand g24696__8428 (n_677, n_680, n_345);
  nand g24695__5526 (n_676, n_680, n_323);
  nand g24694__6783 (n_675, n_680, n_272);
  nand g24697__3680 (n_674, n_680, n_305);
  nor g24698__1617 (n_673, g1097, n_260);
  nor g24700__2802 (n_672, g1097, n_341);
  fflopd g1065_reg(.CK (clock), .D (n_671), .Q (g1065));
  fflopd g13_reg(.CK (clock), .D (n_669), .Q (g5669));
  fflopd g1069_reg(.CK (clock), .D (n_670), .Q (g1069));
  not g24701 (n_680, g1097);
  nand g24759__1705 (n_671, n_659, n_663);
  nand g24760__5122 (n_670, n_647, n_658);
  fflopd g1504_reg(.CK (clock), .D (n_660), .Q (g1504));
  fflopd g1296_reg(.CK (clock), .D (n_656), .Q (new_g3778_));
  fflopd g1462_reg(.CK (clock), .D (n_666), .Q (g1462));
  fflopd g1514_reg(.CK (clock), .D (n_664), .Q (g1514));
  not g24820 (n_669, n_668);
  fflopd g1097_reg(.CK (clock), .D (g_1835), .Q (g1097));
  fflopd g1519_reg(.CK (clock), .D (n_667), .Q (g1519));
  fflopd g1467_reg(.CK (clock), .D (n_661), .Q (g1467));
  fflopd g1509_reg(.CK (clock), .D (n_662), .Q (g1509));
  fflopd g1073_reg(.CK (clock), .D (n_665), .Q (g4267));
  nand g24839__8246 (n_668, n_652, n_651);
  fflopd g1057_reg(.CK (clock), .D (n_655), .Q (g1057));
  fflopd g1328_reg(.CK (clock), .D (n_653), .Q (new_g3779_));
  fflopd g1061_reg(.CK (clock), .D (n_654), .Q (g1061));
  nand g24725__7098 (n_667, n_582, n_642);
  fflopd g1185_reg(.CK (clock), .D (g_1834), .Q (g_1835));
  nand g24724__6131 (n_666, n_649, n_594);
  nand g24772__1881 (n_665, n_560, n_644);
  nand g24726__5115 (n_664, n_638, n_596);
  fflopd g1405_reg(.CK (clock), .D (n_636), .Q (new_g2665_));
  nand g24825__7482 (n_663, n_646, n_639);
  nand g24730__4733 (n_662, n_599, n_645);
  nand g24731__6161 (n_661, n_598, n_650);
  nand g24732__9315 (n_660, n_583, n_641);
  nand g24803__9945 (n_659, g1065, n_657);
  nand g24804__2883 (n_658, g1069, n_657);
  nor g24728__2346 (n_656, g1304, n_643);
  nand g24757__1666 (n_655, n_617, n_625);
  nand g24758__7410 (n_654, n_578, n_623);
  nand g24840__6417 (n_653, n_652, n_628);
  fflopd g1284_reg(.CK (clock), .D (n_627), .Q (new_g3583_));
  fflopd g1041_reg(.CK (clock), .D (n_621), .Q (g1041));
  fflopd g1049_reg(.CK (clock), .D (n_620), .Q (g1049));
  fflopd g1412_reg(.CK (clock), .D (n_635), .Q (new_g2668_));
  fflopd g1130_reg(.CK (clock), .D (n_633), .Q (g1130));
  nand g24881__5477 (n_651, n_12, n_624);
  fflopd g1134_reg(.CK (clock), .D (n_632), .Q (g1134));
  fflopd g1149_reg(.CK (clock), .D (n_619), .Q (g1149));
  fflopd g1138_reg(.CK (clock), .D (n_631), .Q (g1138));
  fflopd g1300_reg(.CK (clock), .D (n_626), .Q (new_g3644_));
  fflopd g1045_reg(.CK (clock), .D (n_630), .Q (g1045));
  fflopd g1432_reg(.CK (clock), .D (n_618), .Q (new_I6791_));
  fflopd g1053_reg(.CK (clock), .D (n_634), .Q (g1053));
  fflopd g1037_reg(.CK (clock), .D (n_629), .Q (g1037));
  nand g24765__2398 (n_650, g1467, n_648);
  nand g24762__5107 (n_649, g1462, n_648);
  nand g24866__6260 (n_647, n_646, n_613);
  nand g24766__4319 (n_645, g1509, n_640);
  nand g24854__8428 (n_644, n_646, n_610);
  fflopd g1230_reg(.CK (clock), .D (n_616), .Q (new_g2752_));
  fflopd g1327_reg(.CK (clock), .D (n_615), .Q (new_g2784_));
  fflopd g1092_reg(.CK (clock), .D (n_611), .Q (g1092));
  wire w, w0, w1, w2;
  nand g24771__5526 (n_643, w0, w2);
  nand g4 (w2, w1, new_g3778_);
  not g1 (w1, n_604);
  nand g0 (w0, w, n_604);
  not g (w, new_g3778_);
  nand g24768__6783 (n_642, g1519, n_637);
  nand g24769__3680 (n_641, g1504, n_640);
  nor g24918__1617 (n_639, n_554, n_609);
  nand g24767__2802 (n_638, g1514, n_637);
  fflopd g1155_reg(.CK (clock), .D (g_1833), .Q (g_1834));
  nor g24729__1705 (n_636, new_g3617_, n_607);
  nand g24876__5122 (n_657, n_595, n_614);
  not g24737 (n_635, n_608);
  nand g24756__8246 (n_634, n_541, n_585);
  nand g24761__7098 (n_633, n_557, n_593);
  nand g24763__6131 (n_632, n_592, n_535);
  nand g24764__1881 (n_631, n_539, n_591);
  nand g24755__5115 (n_630, n_540, n_603);
  nand g24770__7482 (n_629, n_538, n_587);
  wire w3, w4, w5, w6;
  nand g24915__4733 (n_628, w4, w6);
  nand g8 (w6, w5, new_g3779_);
  not g7 (w5, n_576);
  nand g6 (w4, w3, n_576);
  not g5 (w3, new_g3779_);
  fflopd g1494_reg(.CK (clock), .D (n_588), .Q (g1494));
  nor g24745__6161 (n_627, g1304, n_581);
  nor g24738__9315 (n_626, g1304, n_580);
  nand g24801__9945 (n_625, g1057, n_622);
  nand g24942__2883 (n_624, new_g3779_, n_577);
  nand g24802__2346 (n_623, g1061, n_622);
  nand g24739__1666 (n_621, n_548, n_602);
  nand g24740__7410 (n_620, n_550, n_605);
  nand g24743__6417 (n_619, n_549, n_589);
  nand g24796__5477 (n_618, n_475, n_600);
  nand g24865__2398 (n_617, n_646, n_572);
  nand g24841__5107 (n_616, n_493, n_575);
  nand g24907__6260 (n_615, n_652, n_570);
  fflopd g1486_reg(.CK (clock), .D (n_564), .Q (new_I11008_));
  nand g24785__4319 (n_637, n_606, n_574);
  fflopd g1288_reg(.CK (clock), .D (n_568), .Q (new_g3605_));
  fflopd g1280_reg(.CK (clock), .D (n_569), .Q (new_g3568_));
  fflopd g1292_reg(.CK (clock), .D (n_567), .Q (new_g3635_));
  fflopd g1439_reg(.CK (clock), .D (n_571), .Q (g1439));
  nand g24959__8428 (n_614, n_553, n_612);
  nor g24946__5526 (n_613, g1069, n_612);
  nand g24805__6783 (n_611, n_544, n_573);
  not g24954 (n_610, n_579);
  nand g24945__3680 (n_609, g1061, n_612);
  nand g24741__1617 (n_608, n_565, n_496);
  fflopd g1154_reg(.CK (clock), .D (g_1832), .Q (g_1833));
  nand g24744__2802 (n_607, n_430, n_566);
  nand g24786__1705 (n_640, n_606, n_563);
  nand g24787__5122 (n_648, n_606, n_561);
  nand g24799__8246 (n_605, g1049, n_584);
  nand g24843__7098 (n_604, new_g3644_, n_537);
  nand g24798__6131 (n_603, g1045, n_601);
  nand g24797__1881 (n_602, g1041, n_601);
  nand g24869__5115 (n_600, g6675, n_534);
  nand g24776__7482 (n_599, n_285, n_597);
  nand g24775__4733 (n_598, n_597, n_372);
  nand g24774__6161 (n_596, n_597, n_362);
  fflopd g1326_reg(.CK (clock), .D (n_533), .Q (new_g2770_));
  nand g24877__9315 (n_622, n_595, n_555);
  fflopd g1472_reg(.CK (clock), .D (n_546), .Q (g1472));
  fflopd g1499_reg(.CK (clock), .D (n_551), .Q (g1499));
  fflopd g1454_reg(.CK (clock), .D (n_556), .Q (g1454));
  fflopd g1034_reg(.CK (clock), .D (n_543), .Q (g6425));
  nand g24814__9945 (n_594, n_597, n_393);
  nand g24808__2883 (n_593, g1130, n_547);
  nand g24809__2346 (n_592, g1134, n_590);
  nand g24810__1666 (n_591, g1138, n_590);
  nand g24811__7410 (n_589, g1149, n_586);
  nand g24812__6417 (n_588, n_542, n_512);
  nand g24813__5477 (n_587, g1037, n_586);
  nand g24800__2398 (n_585, g1053, n_584);
  nand g24815__5107 (n_583, n_297, n_597);
  nand g24816__6260 (n_582, n_337, n_597);
  wire w7, w8, w9, w10;
  nand g24817__4319 (n_581, w8, w10);
  nand g12 (w10, w9, new_g3583_);
  not g11 (w9, n_523);
  nand g10 (w8, w7, n_523);
  not g9 (w7, new_g3583_);
  wire w11, w12, w13, w14;
  nand g24818__8428 (n_580, w12, w14);
  nand g16 (w14, w13, new_g3644_);
  not g15 (w13, n_536);
  nand g14 (w12, w11, n_536);
  not g13 (w11, new_g3644_);
  nand g24974__5526 (n_579, g1069, n_558);
  nand g24826__6783 (n_578, n_646, n_552);
  not g25007 (n_577, n_576);
  nand g24885__3680 (n_575, g2662, n_516);
  nand g24868__1617 (n_574, n_562, n_392);
  nand g24836__2802 (n_573, g1092, n_559);
  nor g25011__1705 (n_572, n_478, n_530);
  nand g24870__5122 (n_571, n_519, n_465);
  fflopd g1435_reg(.CK (clock), .D (n_522), .Q (g1435));
  fflopd g1077_reg(.CK (clock), .D (n_524), .Q (g1077));
  nand g25026__8246 (n_576, new_g2784_, n_532);
  fflopd g1489_reg(.CK (clock), .D (n_528), .Q (g1489));
  fflopd g1450_reg(.CK (clock), .D (n_517), .Q (g1450));
  wire w15, w16, w17, w18;
  nand g24960__6131 (n_570, w16, w18);
  nand g20 (w18, w17, new_g2784_);
  not g19 (w17, n_531);
  nand g18 (w16, w15, n_531);
  not g17 (w15, new_g2784_);
  nor g24779__1881 (n_569, g1304, n_526);
  nand g24780__5115 (n_568, n_471, n_529);
  nor g24781__7482 (n_567, g1304, n_527);
  nand g24806__4733 (n_566, g1408, new_g2665_);
  nand g24807__6161 (n_565, g1415, new_g2668_);
  fflopd g1153_reg(.CK (clock), .D (n_525), .Q (g_1832));
  wire w19, w20, w21, w22;
  nand g24819__9315 (n_564, w20, w22);
  nand g24 (w22, w21, new_I11008_);
  not g23 (w21, n_545);
  nand g22 (w20, w19, n_545);
  not g21 (w19, new_I11008_);
  nand g24830__9945 (n_563, n_361, n_562);
  nand g24832__2883 (n_561, n_562, n_371);
  nand g24835__2346 (n_560, g4267, n_559);
  not g25008 (n_612, n_558);
  nand g24871__1666 (n_557, n_70, n_646);
  nand g24838__7410 (n_556, n_437, n_511);
  nand g25022__6417 (n_555, n_553, n_554);
  nor g25012__5477 (n_552, g1061, n_554);
  wire w23, w24, w25, w26;
  nand g24852__2398 (n_551, w24, w26);
  nand g28 (w26, w25, g1499);
  not g27 (w25, n_482);
  nand g26 (w24, w23, n_482);
  not g25 (w23, g1499);
  nand g24853__5107 (n_550, n_646, n_460);
  nand g24855__6260 (n_549, n_646, n_298);
  nand g24856__4319 (n_548, n_646, n_379);
  nand g24861__8428 (n_547, n_95, n_595);
  nor g24864__5526 (n_546, n_545, n_495);
  nand g24867__6783 (n_544, n_210, n_646);
  nor g25027__3680 (n_558, n_45, n_554);
  fflopd g1276_reg(.CK (clock), .D (n_506), .Q (new_g3549_));
  fflopd g1229_reg(.CK (clock), .D (n_510), .Q (new_g2734_));
  nor g24773__1617 (n_543, n_184, n_515);
  nand g24833__2802 (n_542, n_136, n_509);
  nand g24828__1705 (n_541, n_646, n_438);
  nand g24829__5122 (n_540, n_646, n_375);
  nand g24824__8246 (n_539, n_646, n_183);
  nand g24822__7098 (n_538, n_646, n_283);
  not g24880 (n_537, n_536);
  nand g24872__6131 (n_535, n_646, n_211);
  not g24903 (n_534, n_521);
  nand g24972__1881 (n_533, n_652, n_513);
  nand g24875__5115 (n_590, n_595, n_175);
  nand g24878__7482 (n_584, n_595, n_435);
  nand g24873__4733 (n_601, n_595, n_370);
  nand g24874__6161 (n_586, n_595, n_278);
  nor g24879__9315 (n_597, g6648, n_545);
  not g25029 (n_532, n_531);
  not g25030 (n_530, n_554);
  not g24850 (n_529, n_514);
  wire w27, w28, w29, w30;
  nand g24857__9945 (n_528, w28, w30);
  nand g32 (w30, w29, n_507);
  not g31 (w29, n_508);
  nand g30 (w28, w27, n_508);
  not g29 (w27, n_507);
  wire w31, w32, w33, w34;
  nand g24858__2883 (n_527, w32, w34);
  nand g36 (w34, w33, new_g3635_);
  not g35 (w33, n_483);
  nand g34 (w32, w31, n_483);
  not g33 (w31, new_g3635_);
  wire w35, w36, w37, w38;
  nand g24859__2346 (n_526, w36, w38);
  nand g40 (w38, w37, new_g3568_);
  not g39 (w37, n_488);
  nand g38 (w36, w35, n_488);
  not g37 (w35, new_g3568_);
  nand g24863__1666 (n_525, n_34, n_498);
  fflopd g1033_reg(.CK (clock), .D (n_503), .Q (g1033));
  fflopd g1357_reg(.CK (clock), .D (n_501), .Q (new_g3757_));
  fflopd g1325_reg(.CK (clock), .D (n_499), .Q (new_g2746_));
  fflopd g1481_reg(.CK (clock), .D (n_491), .Q (g1481));
  fflopd g1444_reg(.CK (clock), .D (n_486), .Q (g1444));
  fflopd g1081_reg(.CK (clock), .D (n_492), .Q (g1944));
  nand g24831__7410 (n_524, n_346, n_500);
  nand g24887__6417 (n_523, new_g3568_, n_489);
  nand g24882__5477 (n_522, n_126, n_520);
  fflopd g1408_reg(.CK (clock), .D (n_494), .Q (g1408));
  fflopd g1415_reg(.CK (clock), .D (n_497), .Q (g1415));
  nand g24908__2398 (n_521, g1439, n_520);
  nand g24909__5107 (n_519, n_7, n_520);
  nand g24924__6260 (n_517, n_487, n_433);
  wire w39, w40, w41, w42;
  nand g24961__4319 (n_516, w40, w42);
  nand g45 (w42, w41, n_68);
  not g44 (w41, n_480);
  nand g42 (w40, w39, n_480);
  not g41 (w39, n_68);
  not g24906 (n_559, n_595);
  nand g24896__8428 (n_536, new_g3635_, n_484);
  fflopd g1272_reg(.CK (clock), .D (n_490), .Q (new_g3533_));
  not g24905 (n_562, n_545);
  not g24851 (n_515, n_504);
  nand g24860__5526 (n_514, n_166, n_473);
  wire w43, w44, w45, w46;
  nand g25013__6783 (n_513, w44, w46);
  nand g50 (w46, w45, new_g2770_);
  not g48 (w45, n_476);
  nand g47 (w44, w43, n_476);
  not g46 (w43, new_g2770_);
  nand g25041__3680 (n_531, new_g2770_, n_477);
  fflopd g38_reg(.CK (clock), .D (n_470), .Q (g5687));
  fflopd g16_reg(.CK (clock), .D (g_1822), .Q (g5678));
  fflopd g33_reg(.CK (clock), .D (n_468), .Q (g5684));
  nand g25042__1617 (n_554, g1057, n_479);
  nand g24920__2802 (n_512, g1494, n_481);
  nand g24922__1705 (n_511, g1450, n_467);
  nor g24935__5122 (n_510, n_255, n_464);
  nor g24912__8246 (n_509, n_507, n_508);
  nor g24834__7098 (n_506, g1304, n_474);
  nor g24926__6131 (n_545, n_508, n_221);
  nand g24927__1881 (n_595, n_553, n_505);
  nor g24928__5115 (n_646, n_505, n_71);
  nand g24862__7482 (n_504, n_154, n_502);
  nand g24837__4733 (n_503, g8234, n_502);
  nor g25020__6161 (n_501, n_439, n_461);
  nor g24883__9315 (n_500, g7424, n_458);
  fflopd g1320_reg(.CK (clock), .D (n_450), .Q (new_g3707_));
  fflopd g1317_reg(.CK (clock), .D (n_445), .Q (new_g3666_));
  fflopd g1321_reg(.CK (clock), .D (n_449), .Q (new_g3728_));
  fflopd g1323_reg(.CK (clock), .D (n_447), .Q (new_g3768_));
  fflopd g1319_reg(.CK (clock), .D (n_451), .Q (new_g3694_));
  fflopd g1318_reg(.CK (clock), .D (n_452), .Q (new_g3684_));
  fflopd g1324_reg(.CK (clock), .D (n_446), .Q (new_g2728_));
  fflopd g1322_reg(.CK (clock), .D (n_454), .Q (new_g3750_));
  fflopd g1313_reg(.CK (clock), .D (n_453), .Q (g1313));
  fflopd g1228_reg(.CK (clock), .D (n_459), .Q (new_g2712_));
  nand g24971__9945 (n_499, n_652, n_462);
  nand g24911__2883 (n_498, new_g2216_, n_463);
  nand g24914__2346 (n_497, n_8, n_496);
  nor g24917__1666 (n_495, g1472, n_448);
  nand g24919__7410 (n_494, n_493, n_456);
  nand g24921__6417 (n_492, n_457, n_90);
  wire w47, w48, w49, w50;
  nand g24923__5477 (n_491, w48, w50);
  nand g54 (w50, w49, g1481);
  not g53 (w49, n_606);
  nand g52 (w48, w47, n_606);
  not g51 (w47, g1481);
  not g24904 (n_490, n_472);
  not g24930 (n_489, n_488);
  nand g24938__2398 (n_487, n_78, n_485);
  nand g24944__5107 (n_486, n_30, n_485);
  not g24956 (n_484, n_483);
  not g24957 (n_482, n_481);
  not g24929 (n_520, n_466);
  nand g25040__6260 (n_480, new_g2734_, n_443);
  not g25062 (n_479, n_478);
  not g25076 (n_477, n_476);
  nand g24931__4319 (n_475, n_469, n_50);
  wire w51, w52, w53, w54;
  nand g24916__8428 (n_474, w52, w54);
  nand g58 (w54, w53, new_g3549_);
  not g57 (w53, n_428);
  nand g56 (w52, w51, n_428);
  not g55 (w51, new_g3549_);
  fflopd g1404_reg(.CK (clock), .D (g_1821), .Q (g_1822));
  wire w55, w56, w57, w58;
  nand g24910__5526 (n_473, w56, w58);
  nand g62 (w58, w57, new_g3605_);
  not g61 (w57, n_426);
  nand g60 (w56, w55, n_426);
  not g59 (w55, new_g3605_);
  nand g24913__6783 (n_472, n_471, n_432);
  fflopd g1354_reg(.CK (clock), .D (n_440), .Q (g1354));
  fflopd g1416_reg(.CK (clock), .D (n_441), .Q (g1416));
  nand g24933__3680 (n_470, n_469, n_198);
  nand g24936__1617 (n_468, n_469, n_127);
  nor g24937__2802 (n_467, g1454, n_444);
  nand g24950__1705 (n_466, g1435, n_469);
  nand g24932__5122 (n_465, n_469, n_120);
  wire w59, w60, w61, w62;
  nand g25010__8246 (n_464, w60, w62);
  nand g66 (w62, w61, new_g2734_);
  not g65 (w61, n_442);
  nand g64 (w60, w59, n_442);
  not g63 (w59, new_g2734_);
  nand g24976__7098 (n_505, new_g2216_, n_606);
  nand g24978__6131 (n_483, new_g3605_, n_427);
  nand g24979__1881 (n_481, n_606, n_188);
  nand g24951__5115 (n_488, new_g3549_, n_429);
  nand g24980__7482 (n_508, g1481, n_606);
  not g24955 (n_463, n_431);
  wire w63, w64, w65, w66;
  nand g25059__4733 (n_462, w64, w66);
  nand g70 (w66, w65, new_g2746_);
  not g69 (w65, n_424);
  nand g68 (w64, w63, n_424);
  not g67 (w63, new_g2746_);
  wire w67, w68, w69, w70;
  nand g25060__6161 (n_461, w68, w70);
  nand g74 (w70, w69, new_g3757_);
  not g73 (w69, n_414);
  nand g72 (w68, w67, n_414);
  not g71 (w67, new_g3757_);
  nor g25066__9315 (n_460, n_390, n_455);
  nand g25021__9945 (n_459, n_493, n_421);
  nand g24939__2883 (n_458, n_385, n_423);
  nand g24941__2346 (n_457, g1944, n_420);
  nor g24943__1666 (n_456, g1428, new_g2665_);
  fflopd g1421_reg(.CK (clock), .D (n_422), .Q (g1421));
  nand g25070__7410 (n_478, g1053, n_455);
  nor g24925__6417 (n_502, n_419, n_338);
  nand g25086__5477 (n_476, new_g2746_, n_425);
  nand g24968__2398 (n_454, n_652, n_344);
  nand g24963__5107 (n_453, g1313, n_652);
  nand g24964__6260 (n_452, n_652, n_128);
  nand g24965__4319 (n_451, n_652, n_200);
  nand g24966__8428 (n_450, n_652, n_246);
  nand g24967__5526 (n_449, n_652, n_301);
  nor g24962__6783 (n_448, g6648, n_360);
  nand g24969__3680 (n_447, n_652, n_381);
  nand g24970__1617 (n_446, n_652, n_417);
  nand g24973__2802 (n_445, n_652, n_116);
  not g25004 (n_485, n_444);
  nor g24977__1705 (n_496, new_g3617_, g1430);
  not g25077 (n_443, n_442);
  nand g25016__5122 (n_441, n_436, n_84);
  nor g25053__8246 (n_440, n_439, n_415);
  nor g25068__7098 (n_438, g1053, n_434);
  nand g25019__6131 (n_437, n_436, n_142);
  nand g25081__1881 (n_435, n_553, n_434);
  fflopd g1250_reg(.CK (clock), .D (n_416), .Q (g6653));
  nand g25023__5115 (n_444, g1444, n_436);
  fflopd g1227_reg(.CK (clock), .D (n_418), .Q (new_g3062_));
  nand g25009__7482 (n_433, n_436, n_176);
  wire w71, w72, w73, w74;
  nand g24958__4733 (n_432, w72, w74);
  nand g78 (w74, w73, new_g2407_);
  not g77 (w73, new_g3533_);
  nand g76 (w72, w71, new_g3533_);
  not g75 (w71, new_g2407_);
  nand g24975__6161 (n_431, g1176, g652);
  not g24982 (n_430, g1428);
  fflopd g1403_reg(.CK (clock), .D (g_1820), .Q (g_1821));
  not g25006 (n_429, n_428);
  not g25005 (n_427, n_426);
  not g24983 (n_469, g1430);
  not g24984 (n_606, g6648);
  not g25088 (n_425, n_424);
  nor g25018__9315 (n_423, g1166, n_330);
  nor g25017__9945 (n_422, new_g2407_, n_64);
  wire w75, w76, w77, w78;
  nand g25048__2883 (n_421, w76, w78);
  nand g82 (w78, w77, new_g2712_);
  not g81 (w77, n_409);
  nand g80 (w76, w75, n_409);
  not g79 (w75, new_g2712_);
  not g25090 (n_455, n_434);
  nand g25025__2346 (n_428, new_g2407_, new_g3533_);
  nand g25024__1666 (n_426, new_g2407_, n_731);
  fflopd g1339_reg(.CK (clock), .D (n_400), .Q (new_g3753_));
  fflopd g1342_reg(.CK (clock), .D (n_405), .Q (new_g3716_));
  fflopd g1333_reg(.CK (clock), .D (n_407), .Q (new_g3712_));
  fflopd g1360_reg(.CK (clock), .D (n_399), .Q (g1360));
  not g24981 (n_420, g1176);
  nor g24940__7410 (n_419, g1000, n_412);
  fflopd g1428_reg(.CK (clock), .D (new_g2407_), .Q (g1428));
  nand g25087__6417 (n_442, new_g2712_, n_410);
  fflopd g1430_reg(.CK (clock), .D (n_411), .Q (g1430));
  fflopd g1351_reg(.CK (clock), .D (n_406), .Q (new_g3769_));
  fflopd g1345_reg(.CK (clock), .D (n_404), .Q (new_g3735_));
  fflopd g1336_reg(.CK (clock), .D (n_408), .Q (new_g3732_));
  fflopd g1348_reg(.CK (clock), .D (n_403), .Q (new_g3754_));
  fflopd g1330_reg(.CK (clock), .D (n_413), .Q (new_g3700_));
  fflopd g1251_reg(.CK (clock), .D (n_402), .Q (g6648));
  not g24985 (n_652, new_g2727_);
  nand g25054__5477 (n_418, n_493, n_394);
  wire w79, w80, w81, w82;
  nand g25083__2398 (n_417, w80, w82);
  nand g86 (w82, w81, new_g2728_);
  not g85 (w81, n_386);
  nand g84 (w80, w79, n_386);
  not g83 (w79, new_g2728_);
  nand g25015__5107 (n_416, g1253, n_401);
  nand g25098__6260 (n_424, new_g2728_, n_387);
  not g25031 (n_436, new_g2407_);
  wire w83, w84, w85, w86;
  nand g25084__4319 (n_415, w84, w86);
  nand g90 (w86, w85, g1354);
  not g89 (w85, n_388);
  nand g88 (w84, w83, n_388);
  not g87 (w83, g1354);
  fflopd g1329_reg(.CK (clock), .D (g1267), .Q (new_g2727_));
  nand g25097__8428 (n_414, g1354, n_389);
  fflopd g1402_reg(.CK (clock), .D (n_721), .Q (g_1820));
  fflopd g1176_reg(.CK (clock), .D (n_397), .Q (g1176));
  nand g25101__5526 (n_434, g1049, n_391);
  nor g25035__6783 (n_413, new_g3700_, n_439);
  nand g25014__3680 (n_412, g999, g998);
  not g25028 (n_411, new_I8094_);
  fflopd g1166_reg(.CK (clock), .D (g7423), .Q (g1166));
  not g25089 (n_410, n_409);
  nor g25039__1617 (n_408, n_439, n_125);
  not g25045 (n_407, n_396);
  fflopd g1307_reg(.CK (clock), .D (n_383), .Q (new_g2407_));
  nor g25052__2802 (n_406, n_439, n_380);
  nor g25049__1705 (n_405, n_439, n_245);
  nor g25050__5122 (n_404, n_439, n_302);
  nor g25051__8246 (n_403, n_439, n_343);
  not g25047 (n_402, n_401);
  nor g25055__7098 (n_400, n_439, n_201);
  not g25046 (n_399, n_395);
  fflopd g1226_reg(.CK (clock), .D (n_382), .Q (new_g3052_));
  fflopd g1084_reg(.CK (clock), .D (n_384), .Q (g2888));
  fflopd g1252_reg(.CK (clock), .D (new_I6864_), .Q (new_I8094_));
  nand g25038__1881 (n_397, n_17, n_367);
  nand g25057__5115 (n_396, new_I8446_, n_52);
  nand g25058__7482 (n_395, new_I8446_, n_334);
  fflopd g1267_reg(.CK (clock), .D (n_377), .Q (g1267));
  nand g25061__4733 (n_401, new_I8446_, n_353);
  wire w87, w88, w89, w90;
  nand g25085__6161 (n_394, w88, w90);
  nand g94 (w90, w89, new_g3062_);
  not g93 (w89, n_373);
  nand g92 (w88, w87, n_373);
  not g91 (w87, new_g3062_);
  nor g25107__9315 (n_393, n_392, n_368);
  not g25118 (n_391, n_390);
  not g25119 (n_389, n_388);
  not g25121 (n_387, n_386);
  not g25064 (n_385, g7423);
  nand g25100__9945 (n_409, new_g3062_, n_374);
  fflopd g999_reg(.CK (clock), .D (n_365), .Q (g999));
  nand g25056__2883 (n_384, n_340, n_366);
  not g25063 (n_383, new_I6864_);
  nand g25080__2346 (n_382, n_493, n_364);
  fflopd g1167_reg(.CK (clock), .D (g7424), .Q (g7423));
  not g25065 (n_439, new_I8446_);
  wire w91, w92, w93, w94;
  nand g25114__1666 (n_381, w92, w94);
  nand g98 (w94, w93, new_g3768_);
  not g97 (w93, n_356);
  nand g96 (w92, w91, n_356);
  not g95 (w91, new_g3768_);
  wire w95, w96, w97, w98;
  nand g25115__7410 (n_380, w96, w98);
  nand g102 (w98, w97, new_g3769_);
  not g101 (w97, n_358);
  nand g100 (w96, w95, n_358);
  not g99 (w95, new_g3769_);
  nor g25126__6417 (n_379, n_310, n_378);
  nand g25132__5477 (n_388, new_g3769_, n_359);
  nand g25136__2398 (n_386, new_g3768_, n_357);
  nand g25130__5107 (n_390, g1045, n_378);
  nor g25067__6260 (n_377, g1268, g1269);
  fflopd g1260_reg(.CK (clock), .D (n_347), .Q (new_I6864_));
  fflopd g1254_reg(.CK (clock), .D (n_348), .Q (g2662));
  fflopd g1247_reg(.CK (clock), .D (n_350), .Q (new_I8446_));
  fflopd g1225_reg(.CK (clock), .D (n_351), .Q (new_g3038_));
  nor g25127__8428 (n_375, g1045, n_369);
  not g25139 (n_374, n_373);
  nor g25145__5526 (n_372, g1467, n_371);
  nand g25147__6783 (n_370, n_553, n_369);
  nand g25148__3680 (n_368, g1519, n_371);
  nor g25082__1617 (n_367, g4371, n_723);
  nand g25079__2802 (n_366, g2888, n_332);
  nor g25078__1705 (n_365, g6425, n_339);
  wire w99, w100, w101, w102;
  nand g25117__5122 (n_364, w100, w102);
  nand g106 (w102, w101, new_g3052_);
  not g105 (w101, n_335);
  nand g104 (w100, w99, n_335);
  not g103 (w99, new_g3052_);
  not g25104 (n_363, n_352);
  fflopd g1170_reg(.CK (clock), .D (g7425), .Q (g7424));
  nor g25122__8246 (n_362, n_361, n_333);
  nand g25144__7098 (n_360, g1467, n_342);
  not g25161 (n_359, n_358);
  not g25159 (n_357, n_356);
  not g25162 (n_378, n_369);
  nand g25156__6131 (n_373, new_g3052_, n_336);
  fflopd g984_reg(.CK (clock), .D (n_329), .Q (g984));
  nand g25095__5115 (n_354, new_g3716_, n_326);
  nand g25112__7482 (n_353, n_709, n_349);
  nand g25105__4733 (n_352, n_725, n_322);
  nand g25108__6161 (n_351, n_493, n_324);
  nand g25109__9315 (n_350, g1263, n_349);
  nand g25110__9945 (n_348, g1257, n_349);
  nand g25111__2883 (n_347, g1266, n_349);
  fflopd g20_reg(.CK (clock), .D (n_313), .Q (g5682));
  not g25120 (n_346, g7425);
  nor g25125__2346 (n_345, n_287, n_314);
  fflopd g1268_reg(.CK (clock), .D (n_318), .Q (g1268));
  wire w103, w104, w105, w106;
  nand g25153__1666 (n_344, w104, w106);
  nand g110 (w106, w105, new_g3750_);
  not g109 (w105, n_315);
  nand g108 (w104, w103, n_315);
  not g107 (w103, new_g3750_);
  wire w107, w108, w109, w110;
  nand g25154__7410 (n_343, w108, w110);
  nand g114 (w110, w109, new_g3754_);
  not g113 (w109, n_319);
  nand g112 (w108, w107, n_319);
  not g111 (w107, new_g3754_);
  nand g25178__6417 (n_358, new_g3754_, n_320);
  nand g25175__5477 (n_356, new_g3750_, n_316);
  not g25091 (n_471, g1304);
  not g25185 (n_371, n_342);
  nand g25179__2398 (n_369, g1041, n_311);
  wire w111, w112, w113, w114;
  nand g25116__5107 (n_341, w112, w114);
  nand g118 (w114, w113, g1142);
  not g117 (w113, n_321);
  nand g116 (w112, w111, n_321);
  not g115 (w111, g1142);
  nand g25113__6260 (n_340, n_15, n_331);
  nand g25106__4319 (n_339, n_309, n_328);
  fflopd g888_reg(.CK (clock), .D (n_304), .Q (g785));
  fflopd g966_reg(.CK (clock), .D (n_338), .Q (g1871));
  fflopd g1224_reg(.CK (clock), .D (n_306), .Q (new_g3029_));
  fflopd g1304_reg(.CK (clock), .D (g_1801), .Q (g1304));
  nor g25188__8428 (n_337, g1519, n_392);
  not g25160 (n_336, n_335);
  wire w115, w116, w117, w118;
  nand g25141__5526 (n_334, w116, w118);
  nand g122 (w118, w117, g1360);
  not g121 (w117, n_312);
  nand g120 (w116, w115, n_312);
  not g119 (w115, g1360);
  nand g25191__6783 (n_333, g1509, n_392);
  nor g25093__3680 (n_332, g1077, n_331);
  nor g25204__1617 (n_342, n_75, n_392);
  fflopd g1173_reg(.CK (clock), .D (n_330), .Q (g7425));
  nor g25143__2802 (n_329, g979, n_328);
  nor g25129__5122 (n_326, n_19, n_290);
  wire w119, w120, w121, w122;
  nand g25151__7098 (n_324, w120, w122);
  nand g126 (w122, w121, new_g3038_);
  not g125 (w121, n_280);
  nand g124 (w120, w119, n_280);
  not g123 (w119, new_g3038_);
  wire w123, w124, w125, w126;
  nand g25149__6131 (n_323, w124, w126);
  nand g130 (w126, w125, g1122);
  not g129 (w125, n_299);
  nand g128 (w124, w123, n_299);
  not g127 (w123, g1122);
  nand g25150__1881 (n_322, g1126, n_321);
  fflopd g1220_reg(.CK (clock), .D (n_286), .Q (new_g2562_));
  not g25211 (n_320, n_319);
  nand g25152__5115 (n_318, n_53, n_282);
  not g25210 (n_316, n_315);
  not g25182 (n_314, n_300);
  nand g25196__4733 (n_313, g1360, n_312);
  not g25207 (n_311, n_310);
  nand g25176__6161 (n_335, new_g3038_, n_281);
  nor g25157__9315 (n_349, new_g2734_, n_291);
  nor g25123__9945 (n_309, g7103, n_274);
  fflopd g1312_reg(.CK (clock), .D (g_1800), .Q (g_1801));
  nand g25140__2883 (n_307, n_273, n_236);
  nand g25146__2346 (n_306, n_493, n_270);
  not g25158 (n_305, n_292);
  nor g25163__1666 (n_304, g785, n_265);
  not g25183 (n_330, n_293);
  nor g25155__7410 (n_331, n_46, n_269);
  fflopd g1389_reg(.CK (clock), .D (g4657), .Q (g6212));
  wire w127, w128, w129, w130;
  nand g25200__6417 (n_302, w128, w130);
  nand g134 (w130, w129, new_g3735_);
  not g133 (w129, n_276);
  nand g132 (w128, w127, n_276);
  not g131 (w127, new_g3735_);
  wire w131, w132, w133, w134;
  nand g25199__5477 (n_301, w132, w134);
  nand g138 (w134, w133, new_g3728_);
  not g137 (w133, n_266);
  nand g136 (w132, w131, n_266);
  not g135 (w131, new_g3728_);
  nand g25193__2398 (n_300, g1118, n_299);
  nor g25219__5107 (n_298, n_208, n_296);
  nor g25239__6260 (n_297, n_206, n_295);
  nand g25222__4319 (n_310, g1037, n_296);
  nand g25228__8428 (n_315, new_g3728_, n_267);
  nand g25229__5526 (n_319, new_g3735_, n_268);
  not g25184 (n_338, n_328);
  nand g25258__6783 (n_392, n_56, n_295);
  nand g25201__1617 (n_293, g1142, n_288);
  nand g25166__2802 (n_292, n_727, n_250);
  nand g25167__1705 (n_291, new_g2712_, n_253);
  nand g25192__5122 (n_290, new_g3732_, n_258);
  nor g25172__7098 (n_287, n_271, n_249);
  nand g25189__6131 (n_286, n_493, n_254);
  fflopd g995_reg(.CK (clock), .D (n_251), .Q (g995));
  fflopd g1214_reg(.CK (clock), .D (n_256), .Q (new_g2584_));
  nor g25248__1881 (n_285, g1509, n_361);
  nor g25216__5115 (n_283, g1037, n_277);
  nor g25197__7482 (n_282, new_g3019_, n_247);
  not g25235 (n_281, n_280);
  nand g25252__4733 (n_278, n_553, n_277);
  nand g25202__6161 (n_321, new_g1616_, n_288);
  nor g25231__9315 (n_312, n_257, n_276);
  nand g25203__9945 (n_328, g43, n_262);
  fflopd g1223_reg(.CK (clock), .D (n_261), .Q (new_g3019_));
  fflopd g973_reg(.CK (clock), .D (n_240), .Q (g973));
  fflopd g1311_reg(.CK (clock), .D (g1246), .Q (g_1800));
  nand g25169__2883 (n_274, n_6, n_243);
  nand g25173__2346 (n_273, n_242, n_160);
  wire w135, w136, w137, w138;
  nand g25186__1666 (n_272, w136, w138);
  nand g142 (w138, w137, g1114);
  not g141 (w137, n_271);
  nand g140 (w136, w135, n_271);
  not g139 (w135, g1114);
  wire w139, w140, w141, w142;
  nand g25194__7410 (n_270, w140, w142);
  nand g146 (w142, w141, new_g3029_);
  not g145 (w141, n_227);
  nand g144 (w140, w139, n_227);
  not g143 (w139, new_g3029_);
  nand g25195__6417 (n_269, g1179, g652);
  fflopd g1217_reg(.CK (clock), .D (n_237), .Q (new_g2573_));
  fflopd g1253_reg(.CK (clock), .D (n_234), .Q (g1253));
  not g25290 (n_268, n_276);
  not g25260 (n_267, n_266);
  nand g25250__5477 (n_265, g866, new_g3124_);
  not g25289 (n_296, n_277);
  not g25264 (n_295, n_361);
  nand g25256__2398 (n_280, new_g3029_, n_228);
  nor g25227__5107 (g4657, n_713, n_231);
  fflopd g1263_reg(.CK (clock), .D (n_229), .Q (g1263));
  nand g25257__6260 (n_299, new_g1616_, n_232);
  wire w143, w144, w145, w146;
  nand g25187__4319 (n_263, w144, w146);
  nand g150 (w146, w145, g1106);
  not g149 (w145, n_235);
  nand g148 (w144, w143, n_235);
  not g147 (w143, g1106);
  not g25234 (n_262, n_244);
  nand g25190__8428 (n_261, n_493, n_224);
  wire w147, w148, w149, w150;
  nand g25198__5526 (n_260, w148, w150);
  nand g154 (w150, w149, g1098);
  not g153 (w149, n_241);
  nand g152 (w148, w147, n_241);
  not g151 (w147, g1098);
  fflopd g1189_reg(.CK (clock), .D (n_233), .Q (g1189));
  nor g25212__6783 (n_258, new_g3712_, n_257);
  nor g25215__3680 (n_256, n_255, n_124);
  fflopd g889_reg(.CK (clock), .D (n_219), .Q (new_g3124_));
  nor g25230__1617 (n_288, n_43, n_248);
  fflopd g1207_reg(.CK (clock), .D (n_215), .Q (new_g2605_));
  fflopd g1211_reg(.CK (clock), .D (n_213), .Q (new_g2298_));
  wire w151, w152, w153, w154;
  nand g25240__2802 (n_254, w152, w154);
  nand g158 (w154, w153, new_g2562_);
  not g157 (w153, n_193);
  nand g156 (w152, w151, n_193);
  not g155 (w151, new_g2562_);
  nor g25241__1705 (n_253, n_48, n_226);
  nand g25246__8246 (n_251, n_159, n_216);
  nand g25249__7098 (n_250, g1110, n_271);
  nand g25251__6131 (n_249, g1114, n_248);
  nand g25253__1881 (n_247, n_88, n_212);
  wire w155, w156, w157, w158;
  nand g25254__5115 (n_246, w156, w158);
  nand g162 (w158, w157, new_g3707_);
  not g161 (w157, n_202);
  nand g160 (w156, w155, n_202);
  not g159 (w155, new_g3707_);
  wire w159, w160, w161, w162;
  nand g25255__7482 (n_245, w160, w162);
  nand g166 (w162, w161, new_g3716_);
  not g165 (w161, n_204);
  nand g164 (w160, w159, n_204);
  not g163 (w159, new_g3716_);
  nand g25278__4733 (n_266, new_g3707_, n_203);
  nand g25310__6161 (n_277, g1149, n_209);
  nand g25311__9315 (n_276, new_g3716_, n_205);
  nand g25284__9945 (n_361, g1504, n_207);
  nand g25237__2883 (n_244, g973, n_239);
  nor g25218__2346 (n_243, g1000, n_199);
  fflopd g1266_reg(.CK (clock), .D (n_189), .Q (g1266));
  nor g25217__1666 (n_242, n_22, n_241);
  fflopd g1245_reg(.CK (clock), .D (g_1796), .Q (g1246));
  fflopd g1179_reg(.CK (clock), .D (g4373), .Q (g1179));
  fflopd g1257_reg(.CK (clock), .D (n_196), .Q (g1257));
  fflopd g940_reg(.CK (clock), .D (n_190), .Q (g940));
  fflopd g990_reg(.CK (clock), .D (n_195), .Q (g990));
  nor g25244__7410 (n_240, g6850, n_239);
  nand g25245__6417 (n_237, n_493, n_197);
  nand g25247__5477 (n_236, g1102, n_235);
  not g25259 (n_234, n_233);
  not g25262 (n_232, n_248);
  nand g25267__2398 (n_231, n_110, n_194);
  fflopd g866_reg(.CK (clock), .D (new_g2959_), .Q (g866));
  not g25286 (n_229, n_214);
  not g25287 (n_228, n_227);
  nand g25293__6260 (n_226, new_g3052_, n_162);
  wire w163, w164, w165, w166;
  nand g25238__4319 (n_225, w164, w166);
  nand g170 (w166, w165, new_g1616_);
  not g169 (w165, g1087);
  nand g168 (w164, w163, g1087);
  not g167 (w163, new_g1616_);
  wire w167, w168, w169, w170;
  nand g25243__8428 (n_224, w168, w170);
  nand g174 (w170, w169, new_g3019_);
  not g173 (w169, n_180);
  nand g172 (w168, w167, n_180);
  not g171 (w167, new_g3019_);
  nand g25265__5526 (n_221, n_93, n_182);
  nor g25269__3680 (n_219, g785, n_187);
  fflopd g1269_reg(.CK (clock), .D (n_173), .Q (g1269));
  nand g25273__1617 (n_233, n_167, n_731);
  not g25263 (g7103, n_239);
  nand g25276__2802 (n_257, new_g3735_, n_729);
  fflopd g1461_reg(.CK (clock), .D (n_161), .Q (g3829));
  nand g25280__1705 (n_248, n_60, n_217);
  nand g25297__5122 (n_216, g6850, n_168);
  nand g25299__8246 (n_215, new_g2605_, n_493);
  nand g25300__7098 (n_214, new_g2298_, n_178);
  nand g25301__6131 (n_213, n_493, n_112);
  nor g25302__1881 (n_212, new_g3038_, n_163);
  nor g25294__5115 (n_211, n_210, n_165);
  not g25312 (n_209, n_208);
  not g25313 (n_207, n_206);
  not g25315 (n_205, n_204);
  not g25316 (n_203, n_202);
  nand g25306__7482 (n_227, new_g3019_, n_181);
  fflopd g985_reg(.CK (clock), .D (n_185), .Q (g985));
  nand g25305__4733 (n_255, g2662, n_493);
  nand g25308__6161 (n_271, new_g1616_, n_217);
  fflopd g874_reg(.CK (clock), .D (n_144), .Q (new_g2959_));
  fflopd g1244_reg(.CK (clock), .D (new_g3617_), .Q (g_1796));
  wire w171, w172, w173, w174;
  nand g25298__9315 (n_201, w172, w174);
  nand g178 (w174, w173, new_g3753_);
  not g177 (w173, n_148);
  nand g176 (w172, w171, n_148);
  not g175 (w171, new_g3753_);
  wire w175, w176, w177, w178;
  nand g25296__9945 (n_200, w176, w178);
  nand g182 (w178, w177, new_g3694_);
  not g181 (w177, n_146);
  nand g180 (w176, w175, n_146);
  not g179 (w175, new_g3694_);
  nand g25303__2883 (n_199, g998, n_92);
  wire w179, w180, w181, w182;
  nand g25291__2346 (n_198, w180, w182);
  nand g186 (w182, w181, g5687);
  not g185 (w181, n_717);
  nand g184 (w180, w179, n_717);
  not g183 (w179, g5687);
  wire w183, w184, w185, w186;
  nand g25292__1666 (n_197, w184, w186);
  nand g190 (w186, w185, new_g2573_);
  not g189 (w185, n_138);
  nand g188 (w184, w183, n_138);
  not g187 (w183, new_g2573_);
  nor g25295__7410 (n_196, new_g2298_, n_156);
  fflopd g871_reg(.CK (clock), .D (n_153), .Q (g871));
  fflopd g936_reg(.CK (clock), .D (n_140), .Q (g936));
  nor g25281__6417 (n_239, g1871, n_151);
  fflopd g1186_reg(.CK (clock), .D (g4372), .Q (g4373));
  fflopd g1158_reg(.CK (clock), .D (g_1829), .Q (new_g2216_));
  nand g25350__5477 (n_195, n_158, n_134);
  nor g25320__2398 (n_194, g1365, n_715);
  nand g25326__5107 (n_193, new_g2573_, n_139);
  not g25343 (n_190, n_171);
  nor g25304__6260 (n_189, new_g2298_, n_177);
  nand g25333__4319 (n_204, new_g3753_, n_149);
  nand g25334__8428 (n_202, new_g3694_, n_147);
  nand g25307__5526 (n_241, new_g1616_, g1087);
  fflopd g1409_reg(.CK (clock), .D (n_152), .Q (g1724));
  nand g25329__6783 (n_208, g1138, n_137);
  nand g25330__3680 (n_206, g1499, n_188);
  nand g25309__1617 (n_235, new_g1616_, n_145);
  nor g25322__2802 (n_187, new_g3124_, n_170);
  nand g25352__1705 (n_186, n_118, n_109);
  nor g25351__5122 (n_185, n_98, n_184);
  nor g25348__8246 (n_183, g1138, n_174);
  nor g25321__7098 (n_182, n_42, n_130);
  not g25345 (n_181, n_180);
  not g25344 (n_178, n_177);
  fflopd g1460_reg(.CK (clock), .D (n_176), .Q (g206));
  not g25317 (n_493, new_g3617_);
  nand g25359__5115 (n_175, n_553, n_174);
  nand g25354__7482 (n_173, new_g2298_, n_117);
  nand g25355__4733 (n_172, n_108, n_133);
  nand g25356__6161 (n_171, g4655, n_170);
  nand g25357__9315 (n_168, n_106, n_119);
  not g25314 (n_167, n_166);
  nand g25358__9945 (n_165, g1130, n_174);
  not g25369 (g7048, g944);
  nand g25361__2883 (n_163, n_87, n_132);
  nor g25362__2346 (n_162, n_62, n_113);
  not g25370 (n_161, n_143);
  nor g25335__1666 (n_217, n_27, n_160);
  nand g25422__7410 (n_159, g995, n_157);
  nand g25423__6417 (n_158, g990, n_157);
  nand g25349__5477 (n_156, new_g2605_, n_135);
  nor g25347__2398 (g7514, n_154, n_150);
  wire w187, w188, w189, w190;
  nand g25365__5107 (n_153, w188, w190);
  nand g194 (w190, w189, g871);
  not g193 (w189, n_105);
  nand g192 (w188, w187, n_105);
  not g191 (w187, g871);
  nand g25360__6260 (n_152, n_40, n_94);
  fflopd g1159_reg(.CK (clock), .D (g_1828), .Q (g_1829));
  nand g25353__4319 (n_151, n_103, n_39);
  fflopd g998_reg(.CK (clock), .D (g_1824), .Q (g998));
  fflopd g1182_reg(.CK (clock), .D (g4370), .Q (g4372));
  fflopd g1231_reg(.CK (clock), .D (g5571), .Q (new_g3617_));
  fflopd g979_reg(.CK (clock), .D (n_150), .Q (g979));
  fflopd g1148_reg(.CK (clock), .D (g_1831), .Q (new_g1616_));
  not g25371 (n_149, n_148);
  not g25372 (n_147, n_146);
  not g25373 (n_145, n_160);
  not g25375 (n_144, n_170);
  fflopd g944_reg(.CK (clock), .D (n_101), .Q (g944));
  nand g25378__8428 (n_143, g1444, n_142);
  not g25401 (n_140, n_131);
  not g25404 (n_139, n_138);
  not g25405 (n_137, n_174);
  not g25403 (n_188, n_136);
  nand g25331__6783 (n_166, new_g3605_, n_104);
  nand g25368__3680 (n_180, n_122, n_135);
  nand g25367__1617 (n_177, n_85, n_135);
  nand g25418__2802 (n_134, g6850, n_82);
  nor g25407__1705 (n_133, g1371, g1375);
  nor g25419__5122 (n_132, new_g3062_, n_69);
  nand g25421__8246 (n_131, g942, n_121);
  nand g25385__7098 (n_130, g1472, n_76);
  wire w191, w192, w193, w194;
  nand g25366__1881 (n_128, w192, w194);
  nand g198 (w194, w193, new_g3684_);
  not g197 (w193, n_115);
  nand g196 (w192, w191, n_115);
  not g195 (w191, new_g3684_);
  wire w195, w196, w197, w198;
  nand g25364__5115 (n_127, w196, w198);
  nand g202 (w198, w197, g5684);
  not g201 (w197, n_126);
  nand g200 (w196, w195, n_126);
  not g199 (w195, g5684);
  wire w199, w200, w201, w202;
  nand g25363__7482 (n_125, w200, w202);
  nand g207 (w202, w201, new_g3732_);
  not g205 (w201, n_72);
  nand g204 (w200, w199, n_72);
  not g203 (w199, new_g3732_);
  wire w203, w204, w205, w206;
  nand g25346__4733 (n_124, w204, w206);
  nand g211 (w206, w205, new_g2584_);
  not g210 (w205, n_111);
  nand g209 (w204, w203, n_111);
  not g208 (w203, new_g2584_);
  nand g25428__6161 (n_138, new_g2584_, n_122);
  nand g25424__9315 (g4655, n_100, n_121);
  fflopd g933_reg(.CK (clock), .D (n_55), .Q (g933));
  nand g25426__9945 (n_136, g1489, n_59);
  nand g25397__2883 (n_160, g1087, n_91);
  nand g25429__2346 (n_174, g1092, n_77);
  not g25400 (n_120, n_96);
  nand g25388__1666 (n_119, g990, n_86);
  nor g25389__7410 (n_118, g1369, g1374);
  nor g25416__6417 (n_117, new_g2573_, n_80);
  nand g25415__5477 (n_116, n_115, n_719);
  nand g25413__5107 (n_113, new_g3029_, n_66);
  nand g25412__6260 (n_112, n_111, n_67);
  nor g25410__4319 (n_110, g1364, g1363);
  nor g25387__8428 (n_109, g1373, g1372);
  nor g25408__5526 (n_108, g1366, g1370);
  not g25402 (n_176, n_97);
  fflopd g652_reg(.CK (clock), .D (g_1844), .Q (g652));
  nand g25396__3680 (n_146, new_g3684_, n_47);
  nand g25395__1617 (n_148, new_g3732_, n_73);
  nor g25393__2802 (n_184, g985, n_106);
  nand g25399__1705 (n_170, g871, n_105);
  nor g25409__5122 (n_104, n_2, n_35);
  nor g25384__8246 (n_103, g969, g972);
  not g25432 (n_101, n_100);
  not g25480 (n_157, n_98);
  not g25475 (n_142, n_79);
  fflopd g1236_reg(.CK (clock), .D (g1894), .Q (g5571));
  nor g25427__7098 (n_135, n_89, n_41);
  fflopd g1005_reg(.CK (clock), .D (g_1823), .Q (g_1824));
  fflopd g1147_reg(.CK (clock), .D (g_1830), .Q (g_1831));
  nand g25425__6131 (n_97, g1450, n_31);
  fflopd g1157_reg(.CK (clock), .D (g_1827), .Q (g_1828));
  nand g25420__1881 (n_96, g1439, n_29);
  nand g25417__5115 (n_95, n_210, n_553);
  nand g25381__7482 (n_94, n_83, g7063);
  nor g25386__4733 (n_93, n_9, n_44);
  nor g25390__6161 (n_150, g979, n_92);
  fflopd g1160_reg(.CK (clock), .D (g4371), .Q (g4370));
  not g25471 (n_91, n_36);
  nand g25433__9315 (n_90, g1080, n_5);
  fflopd g1372_reg(.CK (clock), .D (n_89), .Q (g1372));
  fflopd g1367_reg(.CK (clock), .D (n_65), .Q (g1367));
  fflopd g1370_reg(.CK (clock), .D (n_88), .Q (g1370));
  fflopd g1364_reg(.CK (clock), .D (n_87), .Q (g1364));
  nor g25449__9945 (n_86, g995, n_81);
  fflopd g1375_reg(.CK (clock), .D (n_85), .Q (g1375));
  nand g25458__2883 (n_84, n_63, n_83);
  nor g25459__2346 (n_82, g990, n_81);
  nand g25484__1666 (n_80, new_g2584_, n_61);
  nand g25509__7410 (n_79, g1454, n_78);
  not g25469 (n_77, n_26);
  not g25476 (n_76, n_75);
  not g25479 (n_73, n_72);
  not g25483 (n_71, n_553);
  nor g25486__6417 (n_70, g1130, n_210);
  nand g25494__5477 (n_69, n_68, n_49);
  nand g25495__2398 (n_67, n_85, n_57);
  nor g25502__5107 (n_66, n_68, n_65);
  nand g25516__6260 (n_98, g6850, n_81);
  nand g25464__4319 (n_121, g940, n_1);
  nand g25463__8428 (n_106, g995, n_3);
  nand g25461__5526 (n_64, g1416, n_63);
  fflopd g1366_reg(.CK (clock), .D (n_68), .Q (g1366));
  fflopd g1369_reg(.CK (clock), .D (n_62), .Q (g1369));
  fflopd g1374_reg(.CK (clock), .D (n_61), .Q (g1374));
  not g25474 (n_60, n_33);
  not g25472 (n_59, n_37);
  fflopd g1371_reg(.CK (clock), .D (n_57), .Q (g1371));
  not g25470 (n_56, n_28);
  fflopd g971_reg(.CK (clock), .D (n_154), .Q (g971));
  wire w207, w208, w209, w210;
  nand g25414__6783 (n_55, w208, w210);
  nand g215 (w210, w209, g929);
  not g214 (w209, g933);
  nand g213 (w208, w207, g933);
  not g212 (w207, g929);
  fflopd g1368_reg(.CK (clock), .D (n_53), .Q (g1368));
  wire w211, w212, w213, w214;
  nand g25411__3680 (n_52, w212, w214);
  nand g219 (w214, w213, new_g3700_);
  not g218 (w213, new_g3712_);
  nand g217 (w212, w211, new_g3712_);
  not g216 (w211, new_g3700_);
  nor g25485__2802 (n_50, g1439, g6675);
  fflopd g1365_reg(.CK (clock), .D (n_49), .Q (g1365));
  fflopd g1363_reg(.CK (clock), .D (n_48), .Q (g1363));
  fflopd g1373_reg(.CK (clock), .D (n_24), .Q (g1373));
  not g25481 (n_47, n_115);
  fflopd g646_reg(.CK (clock), .D (n_46), .Q (g_1844));
  not g25482 (n_122, n_111);
  nand g25462__1705 (n_100, g936, n_0);
  not g25478 (n_105, n_25);
  fflopd g929_reg(.CK (clock), .D (n_4), .Q (g929));
  nand g25506__5122 (n_45, g1065, g1061);
  nand g25492__8246 (n_44, g1499, g1494);
  fflopd g1156_reg(.CK (clock), .D (g1944), .Q (g_1827));
  nand g25496__7098 (n_43, g1126, g1122);
  nand g25500__6131 (n_42, g1514, g1489);
  nand g25489__1881 (n_41, new_g2562_, new_g2573_);
  nand g25493__5115 (n_40, g1724, g1416);
  nor g25460__7482 (n_39, g962, g971);
  fflopd g972_reg(.CK (clock), .D (g979), .Q (g972));
  fflopd g1004_reg(.CK (clock), .D (g43), .Q (g_1823));
  nand g25488__4733 (n_38, new_g3583_, new_g3568_);
  fflopd g1240_reg(.CK (clock), .D (g1234), .Q (g1894));
  nand g25515__6161 (n_72, new_g3712_, new_g3700_);
  nand g25510__9315 (n_75, g1462, g1519);
  nand g25517__9945 (n_115, new_g3666_, g1313);
  fflopd g1163_reg(.CK (clock), .D (g4267), .Q (g4371));
  nand g25513__2883 (g8234, g43, g1033);
  nand g25518__2346 (n_111, new_g2298_, new_g2605_);
  nand g25519__1666 (n_553, new_g2216_, g4267);
  nand g25501__7410 (n_37, g1494, g1481);
  nand g25499__6417 (n_36, g1102, g1098);
  nand g25503__5477 (n_35, new_g3644_, new_g3778_);
  nand g25504__2398 (n_34, g1077, g2888);
  nand g25507__5107 (n_33, g1118, g1114);
  nand g25505__6260 (n_32, new_g3757_, g1354);
  fflopd g942_reg(.CK (clock), .D (g941), .Q (g942));
  fflopd g969_reg(.CK (clock), .D (g1871), .Q (g969));
  nor g25457__4319 (n_31, g1454, g1444);
  nand g25490__8428 (n_30, g1454, g1450);
  nor g25487__5526 (n_29, g1435, new_I6791_);
  fflopd g1146_reg(.CK (clock), .D (g2888), .Q (g_1830));
  nand g25498__6783 (n_28, g1514, g1509);
  nand g25491__3680 (n_27, g1110, g1106);
  nand g25497__1617 (n_26, g1134, g1130);
  nand g25514__2802 (n_25, g933, g929);
  nand g25508__1705 (n_92, g43, g984);
  nand g25512__5122 (n_126, g1439, new_I6791_);
  nand g25511__8246 (g7063, new_g2668_, new_g2665_);
  not g25564 (n_24, new_g2573_);
  not g25526 (n_22, g1098);
  not g25555 (n_19, new_g3753_);
  not g25533 (n_17, g4267);
  not g25534 (n_15, g2888);
  not g25537 (n_507, g1489);
  not g25540 (n_48, new_g3062_);
  not g25553 (n_83, g1416);
  not g25562 (n_89, new_g2584_);
  not g25549 (g6223, new_I11008_);
  not g25536 (n_46, new_g2216_);
  not g25543 (n_87, new_g2712_);
  not g25563 (n_65, new_g3019_);
  not g25541 (n_62, new_g3038_);
  not g25546 (n_63, g1421);
  not g25525 (n_81, g985);
  not g25542 (n_154, g6425);
  not g25565 (g6675, new_I6791_);
  not g25567 (g6850, g43);
  not g25521 (n_12, g5669);
  not g25550 (n_9, g1467);
  not g25548 (n_8, new_g2668_);
  not g25535 (n_7, g1439);
  not g25554 (n_6, g979);
  not g25532 (n_5, g1944);
  not g25523 (n_4, g929);
  not g25529 (n_3, g990);
  not g25527 (n_2, new_g3635_);
  not g25520 (n_1, g936);
  not g25545 (n_0, g940);
  not g25557 (n_61, new_g2562_);
  not g25538 (n_88, new_g3052_);
  not g25556 (n_78, g1450);
  not g25539 (n_49, new_g2734_);
  not g25566 (n_53, new_g3029_);
  not g25544 (n_57, new_g2298_);
  not g25560 (n_85, new_g2605_);
  not g25558 (n_68, new_g2752_);
  not g25561 (n_210, g1092);
  not g3 (g6236, n_706);
  nor g2 (n_706, g1189, g5678);
  not g25767 (n_709, n_708);
  nor g25768 (n_708, g1263, g1257);
  nor g25770 (n_710, g1179, g4370);
  not g25771 (n_713, n_712);
  nor g25772 (n_712, n_172, n_186);
  not g25773 (n_715, n_714);
  nor g25774 (n_714, g1368, g1367);
  not g25775 (n_717, n_716);
  nor g25776 (n_716, g5684, n_126);
  not g25777 (n_719, n_718);
  nor g25778 (n_718, new_g3666_, g1313);
  nand g25779 (n_721, g1360, n_720);
  nor g25780 (n_720, n_354, new_g3700_);
  nand g25781 (n_723, n_710, n_722);
  nor g25782 (n_722, g4373, g4372);
  nand g25783 (n_725, g1122, n_724);
  nor g25784 (n_724, n_288, n_299);
  nand g25785 (n_727, g1106, n_726);
  nor g25786 (n_726, n_217, n_235);
  nor g25787 (n_729, n_32, n_728);
  nand g25788 (n_728, new_g3754_, new_g3769_);
  nor g25789 (n_731, n_38, n_730);
  nand g25790 (n_730, new_g3533_, new_g3549_);
endmodule





module fflopd(CK, D, Q);
  input CK, D;
  output Q;
  wire CK, D;
  wire Q;
  wire next_state;
  reg  qi;
  assign #1 Q = qi;
  assign next_state = D;
  always 
    @(posedge CK) 
      qi <= next_state;
  initial 
    qi <= 1'b0;
endmodule